`include "macros.h"

module fft1024
#(
		//--- data bit-width
			parameter width = 24,
		//--- fft size
			parameter size=1024
)
(
		//--- control
			input                   clk, rst, stall,              
		//--- inputs
			input    [width-1:0]    x0_in,                        
			input    [width-1:0]    x1_in,                        
			input    [width-1:0]    x2_in,                        
			input    [width-1:0]    x3_in,                        
			input    [width-1:0]    x4_in,                        
			input    [width-1:0]    x5_in,                        
			input    [width-1:0]    x6_in,                        
			input    [width-1:0]    x7_in,                        
			input    [width-1:0]    x8_in,                        
			input    [width-1:0]    x9_in,                        
			input    [width-1:0]    x10_in,                       
			input    [width-1:0]    x11_in,                       
			input    [width-1:0]    x12_in,                       
			input    [width-1:0]    x13_in,                       
			input    [width-1:0]    x14_in,                       
			input    [width-1:0]    x15_in,                       
			input    [width-1:0]    x16_in,                       
			input    [width-1:0]    x17_in,                       
			input    [width-1:0]    x18_in,                       
			input    [width-1:0]    x19_in,                       
			input    [width-1:0]    x20_in,                       
			input    [width-1:0]    x21_in,                       
			input    [width-1:0]    x22_in,                       
			input    [width-1:0]    x23_in,                       
			input    [width-1:0]    x24_in,                       
			input    [width-1:0]    x25_in,                       
			input    [width-1:0]    x26_in,                       
			input    [width-1:0]    x27_in,                       
			input    [width-1:0]    x28_in,                       
			input    [width-1:0]    x29_in,                       
			input    [width-1:0]    x30_in,                       
			input    [width-1:0]    x31_in,                       
			input    [width-1:0]    x32_in,                       
			input    [width-1:0]    x33_in,                       
			input    [width-1:0]    x34_in,                       
			input    [width-1:0]    x35_in,                       
			input    [width-1:0]    x36_in,                       
			input    [width-1:0]    x37_in,                       
			input    [width-1:0]    x38_in,                       
			input    [width-1:0]    x39_in,                       
			input    [width-1:0]    x40_in,                       
			input    [width-1:0]    x41_in,                       
			input    [width-1:0]    x42_in,                       
			input    [width-1:0]    x43_in,                       
			input    [width-1:0]    x44_in,                       
			input    [width-1:0]    x45_in,                       
			input    [width-1:0]    x46_in,                       
			input    [width-1:0]    x47_in,                       
			input    [width-1:0]    x48_in,                       
			input    [width-1:0]    x49_in,                       
			input    [width-1:0]    x50_in,                       
			input    [width-1:0]    x51_in,                       
			input    [width-1:0]    x52_in,                       
			input    [width-1:0]    x53_in,                       
			input    [width-1:0]    x54_in,                       
			input    [width-1:0]    x55_in,                       
			input    [width-1:0]    x56_in,                       
			input    [width-1:0]    x57_in,                       
			input    [width-1:0]    x58_in,                       
			input    [width-1:0]    x59_in,                       
			input    [width-1:0]    x60_in,                       
			input    [width-1:0]    x61_in,                       
			input    [width-1:0]    x62_in,                       
			input    [width-1:0]    x63_in,                       
			input    [width-1:0]    x64_in,                       
			input    [width-1:0]    x65_in,                       
			input    [width-1:0]    x66_in,                       
			input    [width-1:0]    x67_in,                       
			input    [width-1:0]    x68_in,                       
			input    [width-1:0]    x69_in,                       
			input    [width-1:0]    x70_in,                       
			input    [width-1:0]    x71_in,                       
			input    [width-1:0]    x72_in,                       
			input    [width-1:0]    x73_in,                       
			input    [width-1:0]    x74_in,                       
			input    [width-1:0]    x75_in,                       
			input    [width-1:0]    x76_in,                       
			input    [width-1:0]    x77_in,                       
			input    [width-1:0]    x78_in,                       
			input    [width-1:0]    x79_in,                       
			input    [width-1:0]    x80_in,                       
			input    [width-1:0]    x81_in,                       
			input    [width-1:0]    x82_in,                       
			input    [width-1:0]    x83_in,                       
			input    [width-1:0]    x84_in,                       
			input    [width-1:0]    x85_in,                       
			input    [width-1:0]    x86_in,                       
			input    [width-1:0]    x87_in,                       
			input    [width-1:0]    x88_in,                       
			input    [width-1:0]    x89_in,                       
			input    [width-1:0]    x90_in,                       
			input    [width-1:0]    x91_in,                       
			input    [width-1:0]    x92_in,                       
			input    [width-1:0]    x93_in,                       
			input    [width-1:0]    x94_in,                       
			input    [width-1:0]    x95_in,                       
			input    [width-1:0]    x96_in,                       
			input    [width-1:0]    x97_in,                       
			input    [width-1:0]    x98_in,                       
			input    [width-1:0]    x99_in,                       
			input    [width-1:0]    x100_in,                      
			input    [width-1:0]    x101_in,                      
			input    [width-1:0]    x102_in,                      
			input    [width-1:0]    x103_in,                      
			input    [width-1:0]    x104_in,                      
			input    [width-1:0]    x105_in,                      
			input    [width-1:0]    x106_in,                      
			input    [width-1:0]    x107_in,                      
			input    [width-1:0]    x108_in,                      
			input    [width-1:0]    x109_in,                      
			input    [width-1:0]    x110_in,                      
			input    [width-1:0]    x111_in,                      
			input    [width-1:0]    x112_in,                      
			input    [width-1:0]    x113_in,                      
			input    [width-1:0]    x114_in,                      
			input    [width-1:0]    x115_in,                      
			input    [width-1:0]    x116_in,                      
			input    [width-1:0]    x117_in,                      
			input    [width-1:0]    x118_in,                      
			input    [width-1:0]    x119_in,                      
			input    [width-1:0]    x120_in,                      
			input    [width-1:0]    x121_in,                      
			input    [width-1:0]    x122_in,                      
			input    [width-1:0]    x123_in,                      
			input    [width-1:0]    x124_in,                      
			input    [width-1:0]    x125_in,                      
			input    [width-1:0]    x126_in,                      
			input    [width-1:0]    x127_in,                      
			input    [width-1:0]    x128_in,                      
			input    [width-1:0]    x129_in,                      
			input    [width-1:0]    x130_in,                      
			input    [width-1:0]    x131_in,                      
			input    [width-1:0]    x132_in,                      
			input    [width-1:0]    x133_in,                      
			input    [width-1:0]    x134_in,                      
			input    [width-1:0]    x135_in,                      
			input    [width-1:0]    x136_in,                      
			input    [width-1:0]    x137_in,                      
			input    [width-1:0]    x138_in,                      
			input    [width-1:0]    x139_in,                      
			input    [width-1:0]    x140_in,                      
			input    [width-1:0]    x141_in,                      
			input    [width-1:0]    x142_in,                      
			input    [width-1:0]    x143_in,                      
			input    [width-1:0]    x144_in,                      
			input    [width-1:0]    x145_in,                      
			input    [width-1:0]    x146_in,                      
			input    [width-1:0]    x147_in,                      
			input    [width-1:0]    x148_in,                      
			input    [width-1:0]    x149_in,                      
			input    [width-1:0]    x150_in,                      
			input    [width-1:0]    x151_in,                      
			input    [width-1:0]    x152_in,                      
			input    [width-1:0]    x153_in,                      
			input    [width-1:0]    x154_in,                      
			input    [width-1:0]    x155_in,                      
			input    [width-1:0]    x156_in,                      
			input    [width-1:0]    x157_in,                      
			input    [width-1:0]    x158_in,                      
			input    [width-1:0]    x159_in,                      
			input    [width-1:0]    x160_in,                      
			input    [width-1:0]    x161_in,                      
			input    [width-1:0]    x162_in,                      
			input    [width-1:0]    x163_in,                      
			input    [width-1:0]    x164_in,                      
			input    [width-1:0]    x165_in,                      
			input    [width-1:0]    x166_in,                      
			input    [width-1:0]    x167_in,                      
			input    [width-1:0]    x168_in,                      
			input    [width-1:0]    x169_in,                      
			input    [width-1:0]    x170_in,                      
			input    [width-1:0]    x171_in,                      
			input    [width-1:0]    x172_in,                      
			input    [width-1:0]    x173_in,                      
			input    [width-1:0]    x174_in,                      
			input    [width-1:0]    x175_in,                      
			input    [width-1:0]    x176_in,                      
			input    [width-1:0]    x177_in,                      
			input    [width-1:0]    x178_in,                      
			input    [width-1:0]    x179_in,                      
			input    [width-1:0]    x180_in,                      
			input    [width-1:0]    x181_in,                      
			input    [width-1:0]    x182_in,                      
			input    [width-1:0]    x183_in,                      
			input    [width-1:0]    x184_in,                      
			input    [width-1:0]    x185_in,                      
			input    [width-1:0]    x186_in,                      
			input    [width-1:0]    x187_in,                      
			input    [width-1:0]    x188_in,                      
			input    [width-1:0]    x189_in,                      
			input    [width-1:0]    x190_in,                      
			input    [width-1:0]    x191_in,                      
			input    [width-1:0]    x192_in,                      
			input    [width-1:0]    x193_in,                      
			input    [width-1:0]    x194_in,                      
			input    [width-1:0]    x195_in,                      
			input    [width-1:0]    x196_in,                      
			input    [width-1:0]    x197_in,                      
			input    [width-1:0]    x198_in,                      
			input    [width-1:0]    x199_in,                      
			input    [width-1:0]    x200_in,                      
			input    [width-1:0]    x201_in,                      
			input    [width-1:0]    x202_in,                      
			input    [width-1:0]    x203_in,                      
			input    [width-1:0]    x204_in,                      
			input    [width-1:0]    x205_in,                      
			input    [width-1:0]    x206_in,                      
			input    [width-1:0]    x207_in,                      
			input    [width-1:0]    x208_in,                      
			input    [width-1:0]    x209_in,                      
			input    [width-1:0]    x210_in,                      
			input    [width-1:0]    x211_in,                      
			input    [width-1:0]    x212_in,                      
			input    [width-1:0]    x213_in,                      
			input    [width-1:0]    x214_in,                      
			input    [width-1:0]    x215_in,                      
			input    [width-1:0]    x216_in,                      
			input    [width-1:0]    x217_in,                      
			input    [width-1:0]    x218_in,                      
			input    [width-1:0]    x219_in,                      
			input    [width-1:0]    x220_in,                      
			input    [width-1:0]    x221_in,                      
			input    [width-1:0]    x222_in,                      
			input    [width-1:0]    x223_in,                      
			input    [width-1:0]    x224_in,                      
			input    [width-1:0]    x225_in,                      
			input    [width-1:0]    x226_in,                      
			input    [width-1:0]    x227_in,                      
			input    [width-1:0]    x228_in,                      
			input    [width-1:0]    x229_in,                      
			input    [width-1:0]    x230_in,                      
			input    [width-1:0]    x231_in,                      
			input    [width-1:0]    x232_in,                      
			input    [width-1:0]    x233_in,                      
			input    [width-1:0]    x234_in,                      
			input    [width-1:0]    x235_in,                      
			input    [width-1:0]    x236_in,                      
			input    [width-1:0]    x237_in,                      
			input    [width-1:0]    x238_in,                      
			input    [width-1:0]    x239_in,                      
			input    [width-1:0]    x240_in,                      
			input    [width-1:0]    x241_in,                      
			input    [width-1:0]    x242_in,                      
			input    [width-1:0]    x243_in,                      
			input    [width-1:0]    x244_in,                      
			input    [width-1:0]    x245_in,                      
			input    [width-1:0]    x246_in,                      
			input    [width-1:0]    x247_in,                      
			input    [width-1:0]    x248_in,                      
			input    [width-1:0]    x249_in,                      
			input    [width-1:0]    x250_in,                      
			input    [width-1:0]    x251_in,                      
			input    [width-1:0]    x252_in,                      
			input    [width-1:0]    x253_in,                      
			input    [width-1:0]    x254_in,                      
			input    [width-1:0]    x255_in,                      
			input    [width-1:0]    x256_in,                      
			input    [width-1:0]    x257_in,                      
			input    [width-1:0]    x258_in,                      
			input    [width-1:0]    x259_in,                      
			input    [width-1:0]    x260_in,                      
			input    [width-1:0]    x261_in,                      
			input    [width-1:0]    x262_in,                      
			input    [width-1:0]    x263_in,                      
			input    [width-1:0]    x264_in,                      
			input    [width-1:0]    x265_in,                      
			input    [width-1:0]    x266_in,                      
			input    [width-1:0]    x267_in,                      
			input    [width-1:0]    x268_in,                      
			input    [width-1:0]    x269_in,                      
			input    [width-1:0]    x270_in,                      
			input    [width-1:0]    x271_in,                      
			input    [width-1:0]    x272_in,                      
			input    [width-1:0]    x273_in,                      
			input    [width-1:0]    x274_in,                      
			input    [width-1:0]    x275_in,                      
			input    [width-1:0]    x276_in,                      
			input    [width-1:0]    x277_in,                      
			input    [width-1:0]    x278_in,                      
			input    [width-1:0]    x279_in,                      
			input    [width-1:0]    x280_in,                      
			input    [width-1:0]    x281_in,                      
			input    [width-1:0]    x282_in,                      
			input    [width-1:0]    x283_in,                      
			input    [width-1:0]    x284_in,                      
			input    [width-1:0]    x285_in,                      
			input    [width-1:0]    x286_in,                      
			input    [width-1:0]    x287_in,                      
			input    [width-1:0]    x288_in,                      
			input    [width-1:0]    x289_in,                      
			input    [width-1:0]    x290_in,                      
			input    [width-1:0]    x291_in,                      
			input    [width-1:0]    x292_in,                      
			input    [width-1:0]    x293_in,                      
			input    [width-1:0]    x294_in,                      
			input    [width-1:0]    x295_in,                      
			input    [width-1:0]    x296_in,                      
			input    [width-1:0]    x297_in,                      
			input    [width-1:0]    x298_in,                      
			input    [width-1:0]    x299_in,                      
			input    [width-1:0]    x300_in,                      
			input    [width-1:0]    x301_in,                      
			input    [width-1:0]    x302_in,                      
			input    [width-1:0]    x303_in,                      
			input    [width-1:0]    x304_in,                      
			input    [width-1:0]    x305_in,                      
			input    [width-1:0]    x306_in,                      
			input    [width-1:0]    x307_in,                      
			input    [width-1:0]    x308_in,                      
			input    [width-1:0]    x309_in,                      
			input    [width-1:0]    x310_in,                      
			input    [width-1:0]    x311_in,                      
			input    [width-1:0]    x312_in,                      
			input    [width-1:0]    x313_in,                      
			input    [width-1:0]    x314_in,                      
			input    [width-1:0]    x315_in,                      
			input    [width-1:0]    x316_in,                      
			input    [width-1:0]    x317_in,                      
			input    [width-1:0]    x318_in,                      
			input    [width-1:0]    x319_in,                      
			input    [width-1:0]    x320_in,                      
			input    [width-1:0]    x321_in,                      
			input    [width-1:0]    x322_in,                      
			input    [width-1:0]    x323_in,                      
			input    [width-1:0]    x324_in,                      
			input    [width-1:0]    x325_in,                      
			input    [width-1:0]    x326_in,                      
			input    [width-1:0]    x327_in,                      
			input    [width-1:0]    x328_in,                      
			input    [width-1:0]    x329_in,                      
			input    [width-1:0]    x330_in,                      
			input    [width-1:0]    x331_in,                      
			input    [width-1:0]    x332_in,                      
			input    [width-1:0]    x333_in,                      
			input    [width-1:0]    x334_in,                      
			input    [width-1:0]    x335_in,                      
			input    [width-1:0]    x336_in,                      
			input    [width-1:0]    x337_in,                      
			input    [width-1:0]    x338_in,                      
			input    [width-1:0]    x339_in,                      
			input    [width-1:0]    x340_in,                      
			input    [width-1:0]    x341_in,                      
			input    [width-1:0]    x342_in,                      
			input    [width-1:0]    x343_in,                      
			input    [width-1:0]    x344_in,                      
			input    [width-1:0]    x345_in,                      
			input    [width-1:0]    x346_in,                      
			input    [width-1:0]    x347_in,                      
			input    [width-1:0]    x348_in,                      
			input    [width-1:0]    x349_in,                      
			input    [width-1:0]    x350_in,                      
			input    [width-1:0]    x351_in,                      
			input    [width-1:0]    x352_in,                      
			input    [width-1:0]    x353_in,                      
			input    [width-1:0]    x354_in,                      
			input    [width-1:0]    x355_in,                      
			input    [width-1:0]    x356_in,                      
			input    [width-1:0]    x357_in,                      
			input    [width-1:0]    x358_in,                      
			input    [width-1:0]    x359_in,                      
			input    [width-1:0]    x360_in,                      
			input    [width-1:0]    x361_in,                      
			input    [width-1:0]    x362_in,                      
			input    [width-1:0]    x363_in,                      
			input    [width-1:0]    x364_in,                      
			input    [width-1:0]    x365_in,                      
			input    [width-1:0]    x366_in,                      
			input    [width-1:0]    x367_in,                      
			input    [width-1:0]    x368_in,                      
			input    [width-1:0]    x369_in,                      
			input    [width-1:0]    x370_in,                      
			input    [width-1:0]    x371_in,                      
			input    [width-1:0]    x372_in,                      
			input    [width-1:0]    x373_in,                      
			input    [width-1:0]    x374_in,                      
			input    [width-1:0]    x375_in,                      
			input    [width-1:0]    x376_in,                      
			input    [width-1:0]    x377_in,                      
			input    [width-1:0]    x378_in,                      
			input    [width-1:0]    x379_in,                      
			input    [width-1:0]    x380_in,                      
			input    [width-1:0]    x381_in,                      
			input    [width-1:0]    x382_in,                      
			input    [width-1:0]    x383_in,                      
			input    [width-1:0]    x384_in,                      
			input    [width-1:0]    x385_in,                      
			input    [width-1:0]    x386_in,                      
			input    [width-1:0]    x387_in,                      
			input    [width-1:0]    x388_in,                      
			input    [width-1:0]    x389_in,                      
			input    [width-1:0]    x390_in,                      
			input    [width-1:0]    x391_in,                      
			input    [width-1:0]    x392_in,                      
			input    [width-1:0]    x393_in,                      
			input    [width-1:0]    x394_in,                      
			input    [width-1:0]    x395_in,                      
			input    [width-1:0]    x396_in,                      
			input    [width-1:0]    x397_in,                      
			input    [width-1:0]    x398_in,                      
			input    [width-1:0]    x399_in,                      
			input    [width-1:0]    x400_in,                      
			input    [width-1:0]    x401_in,                      
			input    [width-1:0]    x402_in,                      
			input    [width-1:0]    x403_in,                      
			input    [width-1:0]    x404_in,                      
			input    [width-1:0]    x405_in,                      
			input    [width-1:0]    x406_in,                      
			input    [width-1:0]    x407_in,                      
			input    [width-1:0]    x408_in,                      
			input    [width-1:0]    x409_in,                      
			input    [width-1:0]    x410_in,                      
			input    [width-1:0]    x411_in,                      
			input    [width-1:0]    x412_in,                      
			input    [width-1:0]    x413_in,                      
			input    [width-1:0]    x414_in,                      
			input    [width-1:0]    x415_in,                      
			input    [width-1:0]    x416_in,                      
			input    [width-1:0]    x417_in,                      
			input    [width-1:0]    x418_in,                      
			input    [width-1:0]    x419_in,                      
			input    [width-1:0]    x420_in,                      
			input    [width-1:0]    x421_in,                      
			input    [width-1:0]    x422_in,                      
			input    [width-1:0]    x423_in,                      
			input    [width-1:0]    x424_in,                      
			input    [width-1:0]    x425_in,                      
			input    [width-1:0]    x426_in,                      
			input    [width-1:0]    x427_in,                      
			input    [width-1:0]    x428_in,                      
			input    [width-1:0]    x429_in,                      
			input    [width-1:0]    x430_in,                      
			input    [width-1:0]    x431_in,                      
			input    [width-1:0]    x432_in,                      
			input    [width-1:0]    x433_in,                      
			input    [width-1:0]    x434_in,                      
			input    [width-1:0]    x435_in,                      
			input    [width-1:0]    x436_in,                      
			input    [width-1:0]    x437_in,                      
			input    [width-1:0]    x438_in,                      
			input    [width-1:0]    x439_in,                      
			input    [width-1:0]    x440_in,                      
			input    [width-1:0]    x441_in,                      
			input    [width-1:0]    x442_in,                      
			input    [width-1:0]    x443_in,                      
			input    [width-1:0]    x444_in,                      
			input    [width-1:0]    x445_in,                      
			input    [width-1:0]    x446_in,                      
			input    [width-1:0]    x447_in,                      
			input    [width-1:0]    x448_in,                      
			input    [width-1:0]    x449_in,                      
			input    [width-1:0]    x450_in,                      
			input    [width-1:0]    x451_in,                      
			input    [width-1:0]    x452_in,                      
			input    [width-1:0]    x453_in,                      
			input    [width-1:0]    x454_in,                      
			input    [width-1:0]    x455_in,                      
			input    [width-1:0]    x456_in,                      
			input    [width-1:0]    x457_in,                      
			input    [width-1:0]    x458_in,                      
			input    [width-1:0]    x459_in,                      
			input    [width-1:0]    x460_in,                      
			input    [width-1:0]    x461_in,                      
			input    [width-1:0]    x462_in,                      
			input    [width-1:0]    x463_in,                      
			input    [width-1:0]    x464_in,                      
			input    [width-1:0]    x465_in,                      
			input    [width-1:0]    x466_in,                      
			input    [width-1:0]    x467_in,                      
			input    [width-1:0]    x468_in,                      
			input    [width-1:0]    x469_in,                      
			input    [width-1:0]    x470_in,                      
			input    [width-1:0]    x471_in,                      
			input    [width-1:0]    x472_in,                      
			input    [width-1:0]    x473_in,                      
			input    [width-1:0]    x474_in,                      
			input    [width-1:0]    x475_in,                      
			input    [width-1:0]    x476_in,                      
			input    [width-1:0]    x477_in,                      
			input    [width-1:0]    x478_in,                      
			input    [width-1:0]    x479_in,                      
			input    [width-1:0]    x480_in,                      
			input    [width-1:0]    x481_in,                      
			input    [width-1:0]    x482_in,                      
			input    [width-1:0]    x483_in,                      
			input    [width-1:0]    x484_in,                      
			input    [width-1:0]    x485_in,                      
			input    [width-1:0]    x486_in,                      
			input    [width-1:0]    x487_in,                      
			input    [width-1:0]    x488_in,                      
			input    [width-1:0]    x489_in,                      
			input    [width-1:0]    x490_in,                      
			input    [width-1:0]    x491_in,                      
			input    [width-1:0]    x492_in,                      
			input    [width-1:0]    x493_in,                      
			input    [width-1:0]    x494_in,                      
			input    [width-1:0]    x495_in,                      
			input    [width-1:0]    x496_in,                      
			input    [width-1:0]    x497_in,                      
			input    [width-1:0]    x498_in,                      
			input    [width-1:0]    x499_in,                      
			input    [width-1:0]    x500_in,                      
			input    [width-1:0]    x501_in,                      
			input    [width-1:0]    x502_in,                      
			input    [width-1:0]    x503_in,                      
			input    [width-1:0]    x504_in,                      
			input    [width-1:0]    x505_in,                      
			input    [width-1:0]    x506_in,                      
			input    [width-1:0]    x507_in,                      
			input    [width-1:0]    x508_in,                      
			input    [width-1:0]    x509_in,                      
			input    [width-1:0]    x510_in,                      
			input    [width-1:0]    x511_in,                      
			input    [width-1:0]    x512_in,                      
			input    [width-1:0]    x513_in,                      
			input    [width-1:0]    x514_in,                      
			input    [width-1:0]    x515_in,                      
			input    [width-1:0]    x516_in,                      
			input    [width-1:0]    x517_in,                      
			input    [width-1:0]    x518_in,                      
			input    [width-1:0]    x519_in,                      
			input    [width-1:0]    x520_in,                      
			input    [width-1:0]    x521_in,                      
			input    [width-1:0]    x522_in,                      
			input    [width-1:0]    x523_in,                      
			input    [width-1:0]    x524_in,                      
			input    [width-1:0]    x525_in,                      
			input    [width-1:0]    x526_in,                      
			input    [width-1:0]    x527_in,                      
			input    [width-1:0]    x528_in,                      
			input    [width-1:0]    x529_in,                      
			input    [width-1:0]    x530_in,                      
			input    [width-1:0]    x531_in,                      
			input    [width-1:0]    x532_in,                      
			input    [width-1:0]    x533_in,                      
			input    [width-1:0]    x534_in,                      
			input    [width-1:0]    x535_in,                      
			input    [width-1:0]    x536_in,                      
			input    [width-1:0]    x537_in,                      
			input    [width-1:0]    x538_in,                      
			input    [width-1:0]    x539_in,                      
			input    [width-1:0]    x540_in,                      
			input    [width-1:0]    x541_in,                      
			input    [width-1:0]    x542_in,                      
			input    [width-1:0]    x543_in,                      
			input    [width-1:0]    x544_in,                      
			input    [width-1:0]    x545_in,                      
			input    [width-1:0]    x546_in,                      
			input    [width-1:0]    x547_in,                      
			input    [width-1:0]    x548_in,                      
			input    [width-1:0]    x549_in,                      
			input    [width-1:0]    x550_in,                      
			input    [width-1:0]    x551_in,                      
			input    [width-1:0]    x552_in,                      
			input    [width-1:0]    x553_in,                      
			input    [width-1:0]    x554_in,                      
			input    [width-1:0]    x555_in,                      
			input    [width-1:0]    x556_in,                      
			input    [width-1:0]    x557_in,                      
			input    [width-1:0]    x558_in,                      
			input    [width-1:0]    x559_in,                      
			input    [width-1:0]    x560_in,                      
			input    [width-1:0]    x561_in,                      
			input    [width-1:0]    x562_in,                      
			input    [width-1:0]    x563_in,                      
			input    [width-1:0]    x564_in,                      
			input    [width-1:0]    x565_in,                      
			input    [width-1:0]    x566_in,                      
			input    [width-1:0]    x567_in,                      
			input    [width-1:0]    x568_in,                      
			input    [width-1:0]    x569_in,                      
			input    [width-1:0]    x570_in,                      
			input    [width-1:0]    x571_in,                      
			input    [width-1:0]    x572_in,                      
			input    [width-1:0]    x573_in,                      
			input    [width-1:0]    x574_in,                      
			input    [width-1:0]    x575_in,                      
			input    [width-1:0]    x576_in,                      
			input    [width-1:0]    x577_in,                      
			input    [width-1:0]    x578_in,                      
			input    [width-1:0]    x579_in,                      
			input    [width-1:0]    x580_in,                      
			input    [width-1:0]    x581_in,                      
			input    [width-1:0]    x582_in,                      
			input    [width-1:0]    x583_in,                      
			input    [width-1:0]    x584_in,                      
			input    [width-1:0]    x585_in,                      
			input    [width-1:0]    x586_in,                      
			input    [width-1:0]    x587_in,                      
			input    [width-1:0]    x588_in,                      
			input    [width-1:0]    x589_in,                      
			input    [width-1:0]    x590_in,                      
			input    [width-1:0]    x591_in,                      
			input    [width-1:0]    x592_in,                      
			input    [width-1:0]    x593_in,                      
			input    [width-1:0]    x594_in,                      
			input    [width-1:0]    x595_in,                      
			input    [width-1:0]    x596_in,                      
			input    [width-1:0]    x597_in,                      
			input    [width-1:0]    x598_in,                      
			input    [width-1:0]    x599_in,                      
			input    [width-1:0]    x600_in,                      
			input    [width-1:0]    x601_in,                      
			input    [width-1:0]    x602_in,                      
			input    [width-1:0]    x603_in,                      
			input    [width-1:0]    x604_in,                      
			input    [width-1:0]    x605_in,                      
			input    [width-1:0]    x606_in,                      
			input    [width-1:0]    x607_in,                      
			input    [width-1:0]    x608_in,                      
			input    [width-1:0]    x609_in,                      
			input    [width-1:0]    x610_in,                      
			input    [width-1:0]    x611_in,                      
			input    [width-1:0]    x612_in,                      
			input    [width-1:0]    x613_in,                      
			input    [width-1:0]    x614_in,                      
			input    [width-1:0]    x615_in,                      
			input    [width-1:0]    x616_in,                      
			input    [width-1:0]    x617_in,                      
			input    [width-1:0]    x618_in,                      
			input    [width-1:0]    x619_in,                      
			input    [width-1:0]    x620_in,                      
			input    [width-1:0]    x621_in,                      
			input    [width-1:0]    x622_in,                      
			input    [width-1:0]    x623_in,                      
			input    [width-1:0]    x624_in,                      
			input    [width-1:0]    x625_in,                      
			input    [width-1:0]    x626_in,                      
			input    [width-1:0]    x627_in,                      
			input    [width-1:0]    x628_in,                      
			input    [width-1:0]    x629_in,                      
			input    [width-1:0]    x630_in,                      
			input    [width-1:0]    x631_in,                      
			input    [width-1:0]    x632_in,                      
			input    [width-1:0]    x633_in,                      
			input    [width-1:0]    x634_in,                      
			input    [width-1:0]    x635_in,                      
			input    [width-1:0]    x636_in,                      
			input    [width-1:0]    x637_in,                      
			input    [width-1:0]    x638_in,                      
			input    [width-1:0]    x639_in,                      
			input    [width-1:0]    x640_in,                      
			input    [width-1:0]    x641_in,                      
			input    [width-1:0]    x642_in,                      
			input    [width-1:0]    x643_in,                      
			input    [width-1:0]    x644_in,                      
			input    [width-1:0]    x645_in,                      
			input    [width-1:0]    x646_in,                      
			input    [width-1:0]    x647_in,                      
			input    [width-1:0]    x648_in,                      
			input    [width-1:0]    x649_in,                      
			input    [width-1:0]    x650_in,                      
			input    [width-1:0]    x651_in,                      
			input    [width-1:0]    x652_in,                      
			input    [width-1:0]    x653_in,                      
			input    [width-1:0]    x654_in,                      
			input    [width-1:0]    x655_in,                      
			input    [width-1:0]    x656_in,                      
			input    [width-1:0]    x657_in,                      
			input    [width-1:0]    x658_in,                      
			input    [width-1:0]    x659_in,                      
			input    [width-1:0]    x660_in,                      
			input    [width-1:0]    x661_in,                      
			input    [width-1:0]    x662_in,                      
			input    [width-1:0]    x663_in,                      
			input    [width-1:0]    x664_in,                      
			input    [width-1:0]    x665_in,                      
			input    [width-1:0]    x666_in,                      
			input    [width-1:0]    x667_in,                      
			input    [width-1:0]    x668_in,                      
			input    [width-1:0]    x669_in,                      
			input    [width-1:0]    x670_in,                      
			input    [width-1:0]    x671_in,                      
			input    [width-1:0]    x672_in,                      
			input    [width-1:0]    x673_in,                      
			input    [width-1:0]    x674_in,                      
			input    [width-1:0]    x675_in,                      
			input    [width-1:0]    x676_in,                      
			input    [width-1:0]    x677_in,                      
			input    [width-1:0]    x678_in,                      
			input    [width-1:0]    x679_in,                      
			input    [width-1:0]    x680_in,                      
			input    [width-1:0]    x681_in,                      
			input    [width-1:0]    x682_in,                      
			input    [width-1:0]    x683_in,                      
			input    [width-1:0]    x684_in,                      
			input    [width-1:0]    x685_in,                      
			input    [width-1:0]    x686_in,                      
			input    [width-1:0]    x687_in,                      
			input    [width-1:0]    x688_in,                      
			input    [width-1:0]    x689_in,                      
			input    [width-1:0]    x690_in,                      
			input    [width-1:0]    x691_in,                      
			input    [width-1:0]    x692_in,                      
			input    [width-1:0]    x693_in,                      
			input    [width-1:0]    x694_in,                      
			input    [width-1:0]    x695_in,                      
			input    [width-1:0]    x696_in,                      
			input    [width-1:0]    x697_in,                      
			input    [width-1:0]    x698_in,                      
			input    [width-1:0]    x699_in,                      
			input    [width-1:0]    x700_in,                      
			input    [width-1:0]    x701_in,                      
			input    [width-1:0]    x702_in,                      
			input    [width-1:0]    x703_in,                      
			input    [width-1:0]    x704_in,                      
			input    [width-1:0]    x705_in,                      
			input    [width-1:0]    x706_in,                      
			input    [width-1:0]    x707_in,                      
			input    [width-1:0]    x708_in,                      
			input    [width-1:0]    x709_in,                      
			input    [width-1:0]    x710_in,                      
			input    [width-1:0]    x711_in,                      
			input    [width-1:0]    x712_in,                      
			input    [width-1:0]    x713_in,                      
			input    [width-1:0]    x714_in,                      
			input    [width-1:0]    x715_in,                      
			input    [width-1:0]    x716_in,                      
			input    [width-1:0]    x717_in,                      
			input    [width-1:0]    x718_in,                      
			input    [width-1:0]    x719_in,                      
			input    [width-1:0]    x720_in,                      
			input    [width-1:0]    x721_in,                      
			input    [width-1:0]    x722_in,                      
			input    [width-1:0]    x723_in,                      
			input    [width-1:0]    x724_in,                      
			input    [width-1:0]    x725_in,                      
			input    [width-1:0]    x726_in,                      
			input    [width-1:0]    x727_in,                      
			input    [width-1:0]    x728_in,                      
			input    [width-1:0]    x729_in,                      
			input    [width-1:0]    x730_in,                      
			input    [width-1:0]    x731_in,                      
			input    [width-1:0]    x732_in,                      
			input    [width-1:0]    x733_in,                      
			input    [width-1:0]    x734_in,                      
			input    [width-1:0]    x735_in,                      
			input    [width-1:0]    x736_in,                      
			input    [width-1:0]    x737_in,                      
			input    [width-1:0]    x738_in,                      
			input    [width-1:0]    x739_in,                      
			input    [width-1:0]    x740_in,                      
			input    [width-1:0]    x741_in,                      
			input    [width-1:0]    x742_in,                      
			input    [width-1:0]    x743_in,                      
			input    [width-1:0]    x744_in,                      
			input    [width-1:0]    x745_in,                      
			input    [width-1:0]    x746_in,                      
			input    [width-1:0]    x747_in,                      
			input    [width-1:0]    x748_in,                      
			input    [width-1:0]    x749_in,                      
			input    [width-1:0]    x750_in,                      
			input    [width-1:0]    x751_in,                      
			input    [width-1:0]    x752_in,                      
			input    [width-1:0]    x753_in,                      
			input    [width-1:0]    x754_in,                      
			input    [width-1:0]    x755_in,                      
			input    [width-1:0]    x756_in,                      
			input    [width-1:0]    x757_in,                      
			input    [width-1:0]    x758_in,                      
			input    [width-1:0]    x759_in,                      
			input    [width-1:0]    x760_in,                      
			input    [width-1:0]    x761_in,                      
			input    [width-1:0]    x762_in,                      
			input    [width-1:0]    x763_in,                      
			input    [width-1:0]    x764_in,                      
			input    [width-1:0]    x765_in,                      
			input    [width-1:0]    x766_in,                      
			input    [width-1:0]    x767_in,                      
			input    [width-1:0]    x768_in,                      
			input    [width-1:0]    x769_in,                      
			input    [width-1:0]    x770_in,                      
			input    [width-1:0]    x771_in,                      
			input    [width-1:0]    x772_in,                      
			input    [width-1:0]    x773_in,                      
			input    [width-1:0]    x774_in,                      
			input    [width-1:0]    x775_in,                      
			input    [width-1:0]    x776_in,                      
			input    [width-1:0]    x777_in,                      
			input    [width-1:0]    x778_in,                      
			input    [width-1:0]    x779_in,                      
			input    [width-1:0]    x780_in,                      
			input    [width-1:0]    x781_in,                      
			input    [width-1:0]    x782_in,                      
			input    [width-1:0]    x783_in,                      
			input    [width-1:0]    x784_in,                      
			input    [width-1:0]    x785_in,                      
			input    [width-1:0]    x786_in,                      
			input    [width-1:0]    x787_in,                      
			input    [width-1:0]    x788_in,                      
			input    [width-1:0]    x789_in,                      
			input    [width-1:0]    x790_in,                      
			input    [width-1:0]    x791_in,                      
			input    [width-1:0]    x792_in,                      
			input    [width-1:0]    x793_in,                      
			input    [width-1:0]    x794_in,                      
			input    [width-1:0]    x795_in,                      
			input    [width-1:0]    x796_in,                      
			input    [width-1:0]    x797_in,                      
			input    [width-1:0]    x798_in,                      
			input    [width-1:0]    x799_in,                      
			input    [width-1:0]    x800_in,                      
			input    [width-1:0]    x801_in,                      
			input    [width-1:0]    x802_in,                      
			input    [width-1:0]    x803_in,                      
			input    [width-1:0]    x804_in,                      
			input    [width-1:0]    x805_in,                      
			input    [width-1:0]    x806_in,                      
			input    [width-1:0]    x807_in,                      
			input    [width-1:0]    x808_in,                      
			input    [width-1:0]    x809_in,                      
			input    [width-1:0]    x810_in,                      
			input    [width-1:0]    x811_in,                      
			input    [width-1:0]    x812_in,                      
			input    [width-1:0]    x813_in,                      
			input    [width-1:0]    x814_in,                      
			input    [width-1:0]    x815_in,                      
			input    [width-1:0]    x816_in,                      
			input    [width-1:0]    x817_in,                      
			input    [width-1:0]    x818_in,                      
			input    [width-1:0]    x819_in,                      
			input    [width-1:0]    x820_in,                      
			input    [width-1:0]    x821_in,                      
			input    [width-1:0]    x822_in,                      
			input    [width-1:0]    x823_in,                      
			input    [width-1:0]    x824_in,                      
			input    [width-1:0]    x825_in,                      
			input    [width-1:0]    x826_in,                      
			input    [width-1:0]    x827_in,                      
			input    [width-1:0]    x828_in,                      
			input    [width-1:0]    x829_in,                      
			input    [width-1:0]    x830_in,                      
			input    [width-1:0]    x831_in,                      
			input    [width-1:0]    x832_in,                      
			input    [width-1:0]    x833_in,                      
			input    [width-1:0]    x834_in,                      
			input    [width-1:0]    x835_in,                      
			input    [width-1:0]    x836_in,                      
			input    [width-1:0]    x837_in,                      
			input    [width-1:0]    x838_in,                      
			input    [width-1:0]    x839_in,                      
			input    [width-1:0]    x840_in,                      
			input    [width-1:0]    x841_in,                      
			input    [width-1:0]    x842_in,                      
			input    [width-1:0]    x843_in,                      
			input    [width-1:0]    x844_in,                      
			input    [width-1:0]    x845_in,                      
			input    [width-1:0]    x846_in,                      
			input    [width-1:0]    x847_in,                      
			input    [width-1:0]    x848_in,                      
			input    [width-1:0]    x849_in,                      
			input    [width-1:0]    x850_in,                      
			input    [width-1:0]    x851_in,                      
			input    [width-1:0]    x852_in,                      
			input    [width-1:0]    x853_in,                      
			input    [width-1:0]    x854_in,                      
			input    [width-1:0]    x855_in,                      
			input    [width-1:0]    x856_in,                      
			input    [width-1:0]    x857_in,                      
			input    [width-1:0]    x858_in,                      
			input    [width-1:0]    x859_in,                      
			input    [width-1:0]    x860_in,                      
			input    [width-1:0]    x861_in,                      
			input    [width-1:0]    x862_in,                      
			input    [width-1:0]    x863_in,                      
			input    [width-1:0]    x864_in,                      
			input    [width-1:0]    x865_in,                      
			input    [width-1:0]    x866_in,                      
			input    [width-1:0]    x867_in,                      
			input    [width-1:0]    x868_in,                      
			input    [width-1:0]    x869_in,                      
			input    [width-1:0]    x870_in,                      
			input    [width-1:0]    x871_in,                      
			input    [width-1:0]    x872_in,                      
			input    [width-1:0]    x873_in,                      
			input    [width-1:0]    x874_in,                      
			input    [width-1:0]    x875_in,                      
			input    [width-1:0]    x876_in,                      
			input    [width-1:0]    x877_in,                      
			input    [width-1:0]    x878_in,                      
			input    [width-1:0]    x879_in,                      
			input    [width-1:0]    x880_in,                      
			input    [width-1:0]    x881_in,                      
			input    [width-1:0]    x882_in,                      
			input    [width-1:0]    x883_in,                      
			input    [width-1:0]    x884_in,                      
			input    [width-1:0]    x885_in,                      
			input    [width-1:0]    x886_in,                      
			input    [width-1:0]    x887_in,                      
			input    [width-1:0]    x888_in,                      
			input    [width-1:0]    x889_in,                      
			input    [width-1:0]    x890_in,                      
			input    [width-1:0]    x891_in,                      
			input    [width-1:0]    x892_in,                      
			input    [width-1:0]    x893_in,                      
			input    [width-1:0]    x894_in,                      
			input    [width-1:0]    x895_in,                      
			input    [width-1:0]    x896_in,                      
			input    [width-1:0]    x897_in,                      
			input    [width-1:0]    x898_in,                      
			input    [width-1:0]    x899_in,                      
			input    [width-1:0]    x900_in,                      
			input    [width-1:0]    x901_in,                      
			input    [width-1:0]    x902_in,                      
			input    [width-1:0]    x903_in,                      
			input    [width-1:0]    x904_in,                      
			input    [width-1:0]    x905_in,                      
			input    [width-1:0]    x906_in,                      
			input    [width-1:0]    x907_in,                      
			input    [width-1:0]    x908_in,                      
			input    [width-1:0]    x909_in,                      
			input    [width-1:0]    x910_in,                      
			input    [width-1:0]    x911_in,                      
			input    [width-1:0]    x912_in,                      
			input    [width-1:0]    x913_in,                      
			input    [width-1:0]    x914_in,                      
			input    [width-1:0]    x915_in,                      
			input    [width-1:0]    x916_in,                      
			input    [width-1:0]    x917_in,                      
			input    [width-1:0]    x918_in,                      
			input    [width-1:0]    x919_in,                      
			input    [width-1:0]    x920_in,                      
			input    [width-1:0]    x921_in,                      
			input    [width-1:0]    x922_in,                      
			input    [width-1:0]    x923_in,                      
			input    [width-1:0]    x924_in,                      
			input    [width-1:0]    x925_in,                      
			input    [width-1:0]    x926_in,                      
			input    [width-1:0]    x927_in,                      
			input    [width-1:0]    x928_in,                      
			input    [width-1:0]    x929_in,                      
			input    [width-1:0]    x930_in,                      
			input    [width-1:0]    x931_in,                      
			input    [width-1:0]    x932_in,                      
			input    [width-1:0]    x933_in,                      
			input    [width-1:0]    x934_in,                      
			input    [width-1:0]    x935_in,                      
			input    [width-1:0]    x936_in,                      
			input    [width-1:0]    x937_in,                      
			input    [width-1:0]    x938_in,                      
			input    [width-1:0]    x939_in,                      
			input    [width-1:0]    x940_in,                      
			input    [width-1:0]    x941_in,                      
			input    [width-1:0]    x942_in,                      
			input    [width-1:0]    x943_in,                      
			input    [width-1:0]    x944_in,                      
			input    [width-1:0]    x945_in,                      
			input    [width-1:0]    x946_in,                      
			input    [width-1:0]    x947_in,                      
			input    [width-1:0]    x948_in,                      
			input    [width-1:0]    x949_in,                      
			input    [width-1:0]    x950_in,                      
			input    [width-1:0]    x951_in,                      
			input    [width-1:0]    x952_in,                      
			input    [width-1:0]    x953_in,                      
			input    [width-1:0]    x954_in,                      
			input    [width-1:0]    x955_in,                      
			input    [width-1:0]    x956_in,                      
			input    [width-1:0]    x957_in,                      
			input    [width-1:0]    x958_in,                      
			input    [width-1:0]    x959_in,                      
			input    [width-1:0]    x960_in,                      
			input    [width-1:0]    x961_in,                      
			input    [width-1:0]    x962_in,                      
			input    [width-1:0]    x963_in,                      
			input    [width-1:0]    x964_in,                      
			input    [width-1:0]    x965_in,                      
			input    [width-1:0]    x966_in,                      
			input    [width-1:0]    x967_in,                      
			input    [width-1:0]    x968_in,                      
			input    [width-1:0]    x969_in,                      
			input    [width-1:0]    x970_in,                      
			input    [width-1:0]    x971_in,                      
			input    [width-1:0]    x972_in,                      
			input    [width-1:0]    x973_in,                      
			input    [width-1:0]    x974_in,                      
			input    [width-1:0]    x975_in,                      
			input    [width-1:0]    x976_in,                      
			input    [width-1:0]    x977_in,                      
			input    [width-1:0]    x978_in,                      
			input    [width-1:0]    x979_in,                      
			input    [width-1:0]    x980_in,                      
			input    [width-1:0]    x981_in,                      
			input    [width-1:0]    x982_in,                      
			input    [width-1:0]    x983_in,                      
			input    [width-1:0]    x984_in,                      
			input    [width-1:0]    x985_in,                      
			input    [width-1:0]    x986_in,                      
			input    [width-1:0]    x987_in,                      
			input    [width-1:0]    x988_in,                      
			input    [width-1:0]    x989_in,                      
			input    [width-1:0]    x990_in,                      
			input    [width-1:0]    x991_in,                      
			input    [width-1:0]    x992_in,                      
			input    [width-1:0]    x993_in,                      
			input    [width-1:0]    x994_in,                      
			input    [width-1:0]    x995_in,                      
			input    [width-1:0]    x996_in,                      
			input    [width-1:0]    x997_in,                      
			input    [width-1:0]    x998_in,                      
			input    [width-1:0]    x999_in,                      
			input    [width-1:0]    x1000_in,                     
			input    [width-1:0]    x1001_in,                     
			input    [width-1:0]    x1002_in,                     
			input    [width-1:0]    x1003_in,                     
			input    [width-1:0]    x1004_in,                     
			input    [width-1:0]    x1005_in,                     
			input    [width-1:0]    x1006_in,                     
			input    [width-1:0]    x1007_in,                     
			input    [width-1:0]    x1008_in,                     
			input    [width-1:0]    x1009_in,                     
			input    [width-1:0]    x1010_in,                     
			input    [width-1:0]    x1011_in,                     
			input    [width-1:0]    x1012_in,                     
			input    [width-1:0]    x1013_in,                     
			input    [width-1:0]    x1014_in,                     
			input    [width-1:0]    x1015_in,                     
			input    [width-1:0]    x1016_in,                     
			input    [width-1:0]    x1017_in,                     
			input    [width-1:0]    x1018_in,                     
			input    [width-1:0]    x1019_in,                     
			input    [width-1:0]    x1020_in,                     
			input    [width-1:0]    x1021_in,                     
			input    [width-1:0]    x1022_in,                     
			input    [width-1:0]    x1023_in,                     
		//--- outputs
			output                  stall_out,                    
			output   [width-1:0]    x0_out,                       
			output   [width-1:0]    x1_out,                       
			output   [width-1:0]    x2_out,                       
			output   [width-1:0]    x3_out,                       
			output   [width-1:0]    x4_out,                       
			output   [width-1:0]    x5_out,                       
			output   [width-1:0]    x6_out,                       
			output   [width-1:0]    x7_out,                       
			output   [width-1:0]    x8_out,                       
			output   [width-1:0]    x9_out,                       
			output   [width-1:0]    x10_out,                      
			output   [width-1:0]    x11_out,                      
			output   [width-1:0]    x12_out,                      
			output   [width-1:0]    x13_out,                      
			output   [width-1:0]    x14_out,                      
			output   [width-1:0]    x15_out,                      
			output   [width-1:0]    x16_out,                      
			output   [width-1:0]    x17_out,                      
			output   [width-1:0]    x18_out,                      
			output   [width-1:0]    x19_out,                      
			output   [width-1:0]    x20_out,                      
			output   [width-1:0]    x21_out,                      
			output   [width-1:0]    x22_out,                      
			output   [width-1:0]    x23_out,                      
			output   [width-1:0]    x24_out,                      
			output   [width-1:0]    x25_out,                      
			output   [width-1:0]    x26_out,                      
			output   [width-1:0]    x27_out,                      
			output   [width-1:0]    x28_out,                      
			output   [width-1:0]    x29_out,                      
			output   [width-1:0]    x30_out,                      
			output   [width-1:0]    x31_out,                      
			output   [width-1:0]    x32_out,                      
			output   [width-1:0]    x33_out,                      
			output   [width-1:0]    x34_out,                      
			output   [width-1:0]    x35_out,                      
			output   [width-1:0]    x36_out,                      
			output   [width-1:0]    x37_out,                      
			output   [width-1:0]    x38_out,                      
			output   [width-1:0]    x39_out,                      
			output   [width-1:0]    x40_out,                      
			output   [width-1:0]    x41_out,                      
			output   [width-1:0]    x42_out,                      
			output   [width-1:0]    x43_out,                      
			output   [width-1:0]    x44_out,                      
			output   [width-1:0]    x45_out,                      
			output   [width-1:0]    x46_out,                      
			output   [width-1:0]    x47_out,                      
			output   [width-1:0]    x48_out,                      
			output   [width-1:0]    x49_out,                      
			output   [width-1:0]    x50_out,                      
			output   [width-1:0]    x51_out,                      
			output   [width-1:0]    x52_out,                      
			output   [width-1:0]    x53_out,                      
			output   [width-1:0]    x54_out,                      
			output   [width-1:0]    x55_out,                      
			output   [width-1:0]    x56_out,                      
			output   [width-1:0]    x57_out,                      
			output   [width-1:0]    x58_out,                      
			output   [width-1:0]    x59_out,                      
			output   [width-1:0]    x60_out,                      
			output   [width-1:0]    x61_out,                      
			output   [width-1:0]    x62_out,                      
			output   [width-1:0]    x63_out,                      
			output   [width-1:0]    x64_out,                      
			output   [width-1:0]    x65_out,                      
			output   [width-1:0]    x66_out,                      
			output   [width-1:0]    x67_out,                      
			output   [width-1:0]    x68_out,                      
			output   [width-1:0]    x69_out,                      
			output   [width-1:0]    x70_out,                      
			output   [width-1:0]    x71_out,                      
			output   [width-1:0]    x72_out,                      
			output   [width-1:0]    x73_out,                      
			output   [width-1:0]    x74_out,                      
			output   [width-1:0]    x75_out,                      
			output   [width-1:0]    x76_out,                      
			output   [width-1:0]    x77_out,                      
			output   [width-1:0]    x78_out,                      
			output   [width-1:0]    x79_out,                      
			output   [width-1:0]    x80_out,                      
			output   [width-1:0]    x81_out,                      
			output   [width-1:0]    x82_out,                      
			output   [width-1:0]    x83_out,                      
			output   [width-1:0]    x84_out,                      
			output   [width-1:0]    x85_out,                      
			output   [width-1:0]    x86_out,                      
			output   [width-1:0]    x87_out,                      
			output   [width-1:0]    x88_out,                      
			output   [width-1:0]    x89_out,                      
			output   [width-1:0]    x90_out,                      
			output   [width-1:0]    x91_out,                      
			output   [width-1:0]    x92_out,                      
			output   [width-1:0]    x93_out,                      
			output   [width-1:0]    x94_out,                      
			output   [width-1:0]    x95_out,                      
			output   [width-1:0]    x96_out,                      
			output   [width-1:0]    x97_out,                      
			output   [width-1:0]    x98_out,                      
			output   [width-1:0]    x99_out,                      
			output   [width-1:0]    x100_out,                     
			output   [width-1:0]    x101_out,                     
			output   [width-1:0]    x102_out,                     
			output   [width-1:0]    x103_out,                     
			output   [width-1:0]    x104_out,                     
			output   [width-1:0]    x105_out,                     
			output   [width-1:0]    x106_out,                     
			output   [width-1:0]    x107_out,                     
			output   [width-1:0]    x108_out,                     
			output   [width-1:0]    x109_out,                     
			output   [width-1:0]    x110_out,                     
			output   [width-1:0]    x111_out,                     
			output   [width-1:0]    x112_out,                     
			output   [width-1:0]    x113_out,                     
			output   [width-1:0]    x114_out,                     
			output   [width-1:0]    x115_out,                     
			output   [width-1:0]    x116_out,                     
			output   [width-1:0]    x117_out,                     
			output   [width-1:0]    x118_out,                     
			output   [width-1:0]    x119_out,                     
			output   [width-1:0]    x120_out,                     
			output   [width-1:0]    x121_out,                     
			output   [width-1:0]    x122_out,                     
			output   [width-1:0]    x123_out,                     
			output   [width-1:0]    x124_out,                     
			output   [width-1:0]    x125_out,                     
			output   [width-1:0]    x126_out,                     
			output   [width-1:0]    x127_out,                     
			output   [width-1:0]    x128_out,                     
			output   [width-1:0]    x129_out,                     
			output   [width-1:0]    x130_out,                     
			output   [width-1:0]    x131_out,                     
			output   [width-1:0]    x132_out,                     
			output   [width-1:0]    x133_out,                     
			output   [width-1:0]    x134_out,                     
			output   [width-1:0]    x135_out,                     
			output   [width-1:0]    x136_out,                     
			output   [width-1:0]    x137_out,                     
			output   [width-1:0]    x138_out,                     
			output   [width-1:0]    x139_out,                     
			output   [width-1:0]    x140_out,                     
			output   [width-1:0]    x141_out,                     
			output   [width-1:0]    x142_out,                     
			output   [width-1:0]    x143_out,                     
			output   [width-1:0]    x144_out,                     
			output   [width-1:0]    x145_out,                     
			output   [width-1:0]    x146_out,                     
			output   [width-1:0]    x147_out,                     
			output   [width-1:0]    x148_out,                     
			output   [width-1:0]    x149_out,                     
			output   [width-1:0]    x150_out,                     
			output   [width-1:0]    x151_out,                     
			output   [width-1:0]    x152_out,                     
			output   [width-1:0]    x153_out,                     
			output   [width-1:0]    x154_out,                     
			output   [width-1:0]    x155_out,                     
			output   [width-1:0]    x156_out,                     
			output   [width-1:0]    x157_out,                     
			output   [width-1:0]    x158_out,                     
			output   [width-1:0]    x159_out,                     
			output   [width-1:0]    x160_out,                     
			output   [width-1:0]    x161_out,                     
			output   [width-1:0]    x162_out,                     
			output   [width-1:0]    x163_out,                     
			output   [width-1:0]    x164_out,                     
			output   [width-1:0]    x165_out,                     
			output   [width-1:0]    x166_out,                     
			output   [width-1:0]    x167_out,                     
			output   [width-1:0]    x168_out,                     
			output   [width-1:0]    x169_out,                     
			output   [width-1:0]    x170_out,                     
			output   [width-1:0]    x171_out,                     
			output   [width-1:0]    x172_out,                     
			output   [width-1:0]    x173_out,                     
			output   [width-1:0]    x174_out,                     
			output   [width-1:0]    x175_out,                     
			output   [width-1:0]    x176_out,                     
			output   [width-1:0]    x177_out,                     
			output   [width-1:0]    x178_out,                     
			output   [width-1:0]    x179_out,                     
			output   [width-1:0]    x180_out,                     
			output   [width-1:0]    x181_out,                     
			output   [width-1:0]    x182_out,                     
			output   [width-1:0]    x183_out,                     
			output   [width-1:0]    x184_out,                     
			output   [width-1:0]    x185_out,                     
			output   [width-1:0]    x186_out,                     
			output   [width-1:0]    x187_out,                     
			output   [width-1:0]    x188_out,                     
			output   [width-1:0]    x189_out,                     
			output   [width-1:0]    x190_out,                     
			output   [width-1:0]    x191_out,                     
			output   [width-1:0]    x192_out,                     
			output   [width-1:0]    x193_out,                     
			output   [width-1:0]    x194_out,                     
			output   [width-1:0]    x195_out,                     
			output   [width-1:0]    x196_out,                     
			output   [width-1:0]    x197_out,                     
			output   [width-1:0]    x198_out,                     
			output   [width-1:0]    x199_out,                     
			output   [width-1:0]    x200_out,                     
			output   [width-1:0]    x201_out,                     
			output   [width-1:0]    x202_out,                     
			output   [width-1:0]    x203_out,                     
			output   [width-1:0]    x204_out,                     
			output   [width-1:0]    x205_out,                     
			output   [width-1:0]    x206_out,                     
			output   [width-1:0]    x207_out,                     
			output   [width-1:0]    x208_out,                     
			output   [width-1:0]    x209_out,                     
			output   [width-1:0]    x210_out,                     
			output   [width-1:0]    x211_out,                     
			output   [width-1:0]    x212_out,                     
			output   [width-1:0]    x213_out,                     
			output   [width-1:0]    x214_out,                     
			output   [width-1:0]    x215_out,                     
			output   [width-1:0]    x216_out,                     
			output   [width-1:0]    x217_out,                     
			output   [width-1:0]    x218_out,                     
			output   [width-1:0]    x219_out,                     
			output   [width-1:0]    x220_out,                     
			output   [width-1:0]    x221_out,                     
			output   [width-1:0]    x222_out,                     
			output   [width-1:0]    x223_out,                     
			output   [width-1:0]    x224_out,                     
			output   [width-1:0]    x225_out,                     
			output   [width-1:0]    x226_out,                     
			output   [width-1:0]    x227_out,                     
			output   [width-1:0]    x228_out,                     
			output   [width-1:0]    x229_out,                     
			output   [width-1:0]    x230_out,                     
			output   [width-1:0]    x231_out,                     
			output   [width-1:0]    x232_out,                     
			output   [width-1:0]    x233_out,                     
			output   [width-1:0]    x234_out,                     
			output   [width-1:0]    x235_out,                     
			output   [width-1:0]    x236_out,                     
			output   [width-1:0]    x237_out,                     
			output   [width-1:0]    x238_out,                     
			output   [width-1:0]    x239_out,                     
			output   [width-1:0]    x240_out,                     
			output   [width-1:0]    x241_out,                     
			output   [width-1:0]    x242_out,                     
			output   [width-1:0]    x243_out,                     
			output   [width-1:0]    x244_out,                     
			output   [width-1:0]    x245_out,                     
			output   [width-1:0]    x246_out,                     
			output   [width-1:0]    x247_out,                     
			output   [width-1:0]    x248_out,                     
			output   [width-1:0]    x249_out,                     
			output   [width-1:0]    x250_out,                     
			output   [width-1:0]    x251_out,                     
			output   [width-1:0]    x252_out,                     
			output   [width-1:0]    x253_out,                     
			output   [width-1:0]    x254_out,                     
			output   [width-1:0]    x255_out,                     
			output   [width-1:0]    x256_out,                     
			output   [width-1:0]    x257_out,                     
			output   [width-1:0]    x258_out,                     
			output   [width-1:0]    x259_out,                     
			output   [width-1:0]    x260_out,                     
			output   [width-1:0]    x261_out,                     
			output   [width-1:0]    x262_out,                     
			output   [width-1:0]    x263_out,                     
			output   [width-1:0]    x264_out,                     
			output   [width-1:0]    x265_out,                     
			output   [width-1:0]    x266_out,                     
			output   [width-1:0]    x267_out,                     
			output   [width-1:0]    x268_out,                     
			output   [width-1:0]    x269_out,                     
			output   [width-1:0]    x270_out,                     
			output   [width-1:0]    x271_out,                     
			output   [width-1:0]    x272_out,                     
			output   [width-1:0]    x273_out,                     
			output   [width-1:0]    x274_out,                     
			output   [width-1:0]    x275_out,                     
			output   [width-1:0]    x276_out,                     
			output   [width-1:0]    x277_out,                     
			output   [width-1:0]    x278_out,                     
			output   [width-1:0]    x279_out,                     
			output   [width-1:0]    x280_out,                     
			output   [width-1:0]    x281_out,                     
			output   [width-1:0]    x282_out,                     
			output   [width-1:0]    x283_out,                     
			output   [width-1:0]    x284_out,                     
			output   [width-1:0]    x285_out,                     
			output   [width-1:0]    x286_out,                     
			output   [width-1:0]    x287_out,                     
			output   [width-1:0]    x288_out,                     
			output   [width-1:0]    x289_out,                     
			output   [width-1:0]    x290_out,                     
			output   [width-1:0]    x291_out,                     
			output   [width-1:0]    x292_out,                     
			output   [width-1:0]    x293_out,                     
			output   [width-1:0]    x294_out,                     
			output   [width-1:0]    x295_out,                     
			output   [width-1:0]    x296_out,                     
			output   [width-1:0]    x297_out,                     
			output   [width-1:0]    x298_out,                     
			output   [width-1:0]    x299_out,                     
			output   [width-1:0]    x300_out,                     
			output   [width-1:0]    x301_out,                     
			output   [width-1:0]    x302_out,                     
			output   [width-1:0]    x303_out,                     
			output   [width-1:0]    x304_out,                     
			output   [width-1:0]    x305_out,                     
			output   [width-1:0]    x306_out,                     
			output   [width-1:0]    x307_out,                     
			output   [width-1:0]    x308_out,                     
			output   [width-1:0]    x309_out,                     
			output   [width-1:0]    x310_out,                     
			output   [width-1:0]    x311_out,                     
			output   [width-1:0]    x312_out,                     
			output   [width-1:0]    x313_out,                     
			output   [width-1:0]    x314_out,                     
			output   [width-1:0]    x315_out,                     
			output   [width-1:0]    x316_out,                     
			output   [width-1:0]    x317_out,                     
			output   [width-1:0]    x318_out,                     
			output   [width-1:0]    x319_out,                     
			output   [width-1:0]    x320_out,                     
			output   [width-1:0]    x321_out,                     
			output   [width-1:0]    x322_out,                     
			output   [width-1:0]    x323_out,                     
			output   [width-1:0]    x324_out,                     
			output   [width-1:0]    x325_out,                     
			output   [width-1:0]    x326_out,                     
			output   [width-1:0]    x327_out,                     
			output   [width-1:0]    x328_out,                     
			output   [width-1:0]    x329_out,                     
			output   [width-1:0]    x330_out,                     
			output   [width-1:0]    x331_out,                     
			output   [width-1:0]    x332_out,                     
			output   [width-1:0]    x333_out,                     
			output   [width-1:0]    x334_out,                     
			output   [width-1:0]    x335_out,                     
			output   [width-1:0]    x336_out,                     
			output   [width-1:0]    x337_out,                     
			output   [width-1:0]    x338_out,                     
			output   [width-1:0]    x339_out,                     
			output   [width-1:0]    x340_out,                     
			output   [width-1:0]    x341_out,                     
			output   [width-1:0]    x342_out,                     
			output   [width-1:0]    x343_out,                     
			output   [width-1:0]    x344_out,                     
			output   [width-1:0]    x345_out,                     
			output   [width-1:0]    x346_out,                     
			output   [width-1:0]    x347_out,                     
			output   [width-1:0]    x348_out,                     
			output   [width-1:0]    x349_out,                     
			output   [width-1:0]    x350_out,                     
			output   [width-1:0]    x351_out,                     
			output   [width-1:0]    x352_out,                     
			output   [width-1:0]    x353_out,                     
			output   [width-1:0]    x354_out,                     
			output   [width-1:0]    x355_out,                     
			output   [width-1:0]    x356_out,                     
			output   [width-1:0]    x357_out,                     
			output   [width-1:0]    x358_out,                     
			output   [width-1:0]    x359_out,                     
			output   [width-1:0]    x360_out,                     
			output   [width-1:0]    x361_out,                     
			output   [width-1:0]    x362_out,                     
			output   [width-1:0]    x363_out,                     
			output   [width-1:0]    x364_out,                     
			output   [width-1:0]    x365_out,                     
			output   [width-1:0]    x366_out,                     
			output   [width-1:0]    x367_out,                     
			output   [width-1:0]    x368_out,                     
			output   [width-1:0]    x369_out,                     
			output   [width-1:0]    x370_out,                     
			output   [width-1:0]    x371_out,                     
			output   [width-1:0]    x372_out,                     
			output   [width-1:0]    x373_out,                     
			output   [width-1:0]    x374_out,                     
			output   [width-1:0]    x375_out,                     
			output   [width-1:0]    x376_out,                     
			output   [width-1:0]    x377_out,                     
			output   [width-1:0]    x378_out,                     
			output   [width-1:0]    x379_out,                     
			output   [width-1:0]    x380_out,                     
			output   [width-1:0]    x381_out,                     
			output   [width-1:0]    x382_out,                     
			output   [width-1:0]    x383_out,                     
			output   [width-1:0]    x384_out,                     
			output   [width-1:0]    x385_out,                     
			output   [width-1:0]    x386_out,                     
			output   [width-1:0]    x387_out,                     
			output   [width-1:0]    x388_out,                     
			output   [width-1:0]    x389_out,                     
			output   [width-1:0]    x390_out,                     
			output   [width-1:0]    x391_out,                     
			output   [width-1:0]    x392_out,                     
			output   [width-1:0]    x393_out,                     
			output   [width-1:0]    x394_out,                     
			output   [width-1:0]    x395_out,                     
			output   [width-1:0]    x396_out,                     
			output   [width-1:0]    x397_out,                     
			output   [width-1:0]    x398_out,                     
			output   [width-1:0]    x399_out,                     
			output   [width-1:0]    x400_out,                     
			output   [width-1:0]    x401_out,                     
			output   [width-1:0]    x402_out,                     
			output   [width-1:0]    x403_out,                     
			output   [width-1:0]    x404_out,                     
			output   [width-1:0]    x405_out,                     
			output   [width-1:0]    x406_out,                     
			output   [width-1:0]    x407_out,                     
			output   [width-1:0]    x408_out,                     
			output   [width-1:0]    x409_out,                     
			output   [width-1:0]    x410_out,                     
			output   [width-1:0]    x411_out,                     
			output   [width-1:0]    x412_out,                     
			output   [width-1:0]    x413_out,                     
			output   [width-1:0]    x414_out,                     
			output   [width-1:0]    x415_out,                     
			output   [width-1:0]    x416_out,                     
			output   [width-1:0]    x417_out,                     
			output   [width-1:0]    x418_out,                     
			output   [width-1:0]    x419_out,                     
			output   [width-1:0]    x420_out,                     
			output   [width-1:0]    x421_out,                     
			output   [width-1:0]    x422_out,                     
			output   [width-1:0]    x423_out,                     
			output   [width-1:0]    x424_out,                     
			output   [width-1:0]    x425_out,                     
			output   [width-1:0]    x426_out,                     
			output   [width-1:0]    x427_out,                     
			output   [width-1:0]    x428_out,                     
			output   [width-1:0]    x429_out,                     
			output   [width-1:0]    x430_out,                     
			output   [width-1:0]    x431_out,                     
			output   [width-1:0]    x432_out,                     
			output   [width-1:0]    x433_out,                     
			output   [width-1:0]    x434_out,                     
			output   [width-1:0]    x435_out,                     
			output   [width-1:0]    x436_out,                     
			output   [width-1:0]    x437_out,                     
			output   [width-1:0]    x438_out,                     
			output   [width-1:0]    x439_out,                     
			output   [width-1:0]    x440_out,                     
			output   [width-1:0]    x441_out,                     
			output   [width-1:0]    x442_out,                     
			output   [width-1:0]    x443_out,                     
			output   [width-1:0]    x444_out,                     
			output   [width-1:0]    x445_out,                     
			output   [width-1:0]    x446_out,                     
			output   [width-1:0]    x447_out,                     
			output   [width-1:0]    x448_out,                     
			output   [width-1:0]    x449_out,                     
			output   [width-1:0]    x450_out,                     
			output   [width-1:0]    x451_out,                     
			output   [width-1:0]    x452_out,                     
			output   [width-1:0]    x453_out,                     
			output   [width-1:0]    x454_out,                     
			output   [width-1:0]    x455_out,                     
			output   [width-1:0]    x456_out,                     
			output   [width-1:0]    x457_out,                     
			output   [width-1:0]    x458_out,                     
			output   [width-1:0]    x459_out,                     
			output   [width-1:0]    x460_out,                     
			output   [width-1:0]    x461_out,                     
			output   [width-1:0]    x462_out,                     
			output   [width-1:0]    x463_out,                     
			output   [width-1:0]    x464_out,                     
			output   [width-1:0]    x465_out,                     
			output   [width-1:0]    x466_out,                     
			output   [width-1:0]    x467_out,                     
			output   [width-1:0]    x468_out,                     
			output   [width-1:0]    x469_out,                     
			output   [width-1:0]    x470_out,                     
			output   [width-1:0]    x471_out,                     
			output   [width-1:0]    x472_out,                     
			output   [width-1:0]    x473_out,                     
			output   [width-1:0]    x474_out,                     
			output   [width-1:0]    x475_out,                     
			output   [width-1:0]    x476_out,                     
			output   [width-1:0]    x477_out,                     
			output   [width-1:0]    x478_out,                     
			output   [width-1:0]    x479_out,                     
			output   [width-1:0]    x480_out,                     
			output   [width-1:0]    x481_out,                     
			output   [width-1:0]    x482_out,                     
			output   [width-1:0]    x483_out,                     
			output   [width-1:0]    x484_out,                     
			output   [width-1:0]    x485_out,                     
			output   [width-1:0]    x486_out,                     
			output   [width-1:0]    x487_out,                     
			output   [width-1:0]    x488_out,                     
			output   [width-1:0]    x489_out,                     
			output   [width-1:0]    x490_out,                     
			output   [width-1:0]    x491_out,                     
			output   [width-1:0]    x492_out,                     
			output   [width-1:0]    x493_out,                     
			output   [width-1:0]    x494_out,                     
			output   [width-1:0]    x495_out,                     
			output   [width-1:0]    x496_out,                     
			output   [width-1:0]    x497_out,                     
			output   [width-1:0]    x498_out,                     
			output   [width-1:0]    x499_out,                     
			output   [width-1:0]    x500_out,                     
			output   [width-1:0]    x501_out,                     
			output   [width-1:0]    x502_out,                     
			output   [width-1:0]    x503_out,                     
			output   [width-1:0]    x504_out,                     
			output   [width-1:0]    x505_out,                     
			output   [width-1:0]    x506_out,                     
			output   [width-1:0]    x507_out,                     
			output   [width-1:0]    x508_out,                     
			output   [width-1:0]    x509_out,                     
			output   [width-1:0]    x510_out,                     
			output   [width-1:0]    x511_out,                     
			output   [width-1:0]    x512_out,                     
			output   [width-1:0]    x513_out,                     
			output   [width-1:0]    x514_out,                     
			output   [width-1:0]    x515_out,                     
			output   [width-1:0]    x516_out,                     
			output   [width-1:0]    x517_out,                     
			output   [width-1:0]    x518_out,                     
			output   [width-1:0]    x519_out,                     
			output   [width-1:0]    x520_out,                     
			output   [width-1:0]    x521_out,                     
			output   [width-1:0]    x522_out,                     
			output   [width-1:0]    x523_out,                     
			output   [width-1:0]    x524_out,                     
			output   [width-1:0]    x525_out,                     
			output   [width-1:0]    x526_out,                     
			output   [width-1:0]    x527_out,                     
			output   [width-1:0]    x528_out,                     
			output   [width-1:0]    x529_out,                     
			output   [width-1:0]    x530_out,                     
			output   [width-1:0]    x531_out,                     
			output   [width-1:0]    x532_out,                     
			output   [width-1:0]    x533_out,                     
			output   [width-1:0]    x534_out,                     
			output   [width-1:0]    x535_out,                     
			output   [width-1:0]    x536_out,                     
			output   [width-1:0]    x537_out,                     
			output   [width-1:0]    x538_out,                     
			output   [width-1:0]    x539_out,                     
			output   [width-1:0]    x540_out,                     
			output   [width-1:0]    x541_out,                     
			output   [width-1:0]    x542_out,                     
			output   [width-1:0]    x543_out,                     
			output   [width-1:0]    x544_out,                     
			output   [width-1:0]    x545_out,                     
			output   [width-1:0]    x546_out,                     
			output   [width-1:0]    x547_out,                     
			output   [width-1:0]    x548_out,                     
			output   [width-1:0]    x549_out,                     
			output   [width-1:0]    x550_out,                     
			output   [width-1:0]    x551_out,                     
			output   [width-1:0]    x552_out,                     
			output   [width-1:0]    x553_out,                     
			output   [width-1:0]    x554_out,                     
			output   [width-1:0]    x555_out,                     
			output   [width-1:0]    x556_out,                     
			output   [width-1:0]    x557_out,                     
			output   [width-1:0]    x558_out,                     
			output   [width-1:0]    x559_out,                     
			output   [width-1:0]    x560_out,                     
			output   [width-1:0]    x561_out,                     
			output   [width-1:0]    x562_out,                     
			output   [width-1:0]    x563_out,                     
			output   [width-1:0]    x564_out,                     
			output   [width-1:0]    x565_out,                     
			output   [width-1:0]    x566_out,                     
			output   [width-1:0]    x567_out,                     
			output   [width-1:0]    x568_out,                     
			output   [width-1:0]    x569_out,                     
			output   [width-1:0]    x570_out,                     
			output   [width-1:0]    x571_out,                     
			output   [width-1:0]    x572_out,                     
			output   [width-1:0]    x573_out,                     
			output   [width-1:0]    x574_out,                     
			output   [width-1:0]    x575_out,                     
			output   [width-1:0]    x576_out,                     
			output   [width-1:0]    x577_out,                     
			output   [width-1:0]    x578_out,                     
			output   [width-1:0]    x579_out,                     
			output   [width-1:0]    x580_out,                     
			output   [width-1:0]    x581_out,                     
			output   [width-1:0]    x582_out,                     
			output   [width-1:0]    x583_out,                     
			output   [width-1:0]    x584_out,                     
			output   [width-1:0]    x585_out,                     
			output   [width-1:0]    x586_out,                     
			output   [width-1:0]    x587_out,                     
			output   [width-1:0]    x588_out,                     
			output   [width-1:0]    x589_out,                     
			output   [width-1:0]    x590_out,                     
			output   [width-1:0]    x591_out,                     
			output   [width-1:0]    x592_out,                     
			output   [width-1:0]    x593_out,                     
			output   [width-1:0]    x594_out,                     
			output   [width-1:0]    x595_out,                     
			output   [width-1:0]    x596_out,                     
			output   [width-1:0]    x597_out,                     
			output   [width-1:0]    x598_out,                     
			output   [width-1:0]    x599_out,                     
			output   [width-1:0]    x600_out,                     
			output   [width-1:0]    x601_out,                     
			output   [width-1:0]    x602_out,                     
			output   [width-1:0]    x603_out,                     
			output   [width-1:0]    x604_out,                     
			output   [width-1:0]    x605_out,                     
			output   [width-1:0]    x606_out,                     
			output   [width-1:0]    x607_out,                     
			output   [width-1:0]    x608_out,                     
			output   [width-1:0]    x609_out,                     
			output   [width-1:0]    x610_out,                     
			output   [width-1:0]    x611_out,                     
			output   [width-1:0]    x612_out,                     
			output   [width-1:0]    x613_out,                     
			output   [width-1:0]    x614_out,                     
			output   [width-1:0]    x615_out,                     
			output   [width-1:0]    x616_out,                     
			output   [width-1:0]    x617_out,                     
			output   [width-1:0]    x618_out,                     
			output   [width-1:0]    x619_out,                     
			output   [width-1:0]    x620_out,                     
			output   [width-1:0]    x621_out,                     
			output   [width-1:0]    x622_out,                     
			output   [width-1:0]    x623_out,                     
			output   [width-1:0]    x624_out,                     
			output   [width-1:0]    x625_out,                     
			output   [width-1:0]    x626_out,                     
			output   [width-1:0]    x627_out,                     
			output   [width-1:0]    x628_out,                     
			output   [width-1:0]    x629_out,                     
			output   [width-1:0]    x630_out,                     
			output   [width-1:0]    x631_out,                     
			output   [width-1:0]    x632_out,                     
			output   [width-1:0]    x633_out,                     
			output   [width-1:0]    x634_out,                     
			output   [width-1:0]    x635_out,                     
			output   [width-1:0]    x636_out,                     
			output   [width-1:0]    x637_out,                     
			output   [width-1:0]    x638_out,                     
			output   [width-1:0]    x639_out,                     
			output   [width-1:0]    x640_out,                     
			output   [width-1:0]    x641_out,                     
			output   [width-1:0]    x642_out,                     
			output   [width-1:0]    x643_out,                     
			output   [width-1:0]    x644_out,                     
			output   [width-1:0]    x645_out,                     
			output   [width-1:0]    x646_out,                     
			output   [width-1:0]    x647_out,                     
			output   [width-1:0]    x648_out,                     
			output   [width-1:0]    x649_out,                     
			output   [width-1:0]    x650_out,                     
			output   [width-1:0]    x651_out,                     
			output   [width-1:0]    x652_out,                     
			output   [width-1:0]    x653_out,                     
			output   [width-1:0]    x654_out,                     
			output   [width-1:0]    x655_out,                     
			output   [width-1:0]    x656_out,                     
			output   [width-1:0]    x657_out,                     
			output   [width-1:0]    x658_out,                     
			output   [width-1:0]    x659_out,                     
			output   [width-1:0]    x660_out,                     
			output   [width-1:0]    x661_out,                     
			output   [width-1:0]    x662_out,                     
			output   [width-1:0]    x663_out,                     
			output   [width-1:0]    x664_out,                     
			output   [width-1:0]    x665_out,                     
			output   [width-1:0]    x666_out,                     
			output   [width-1:0]    x667_out,                     
			output   [width-1:0]    x668_out,                     
			output   [width-1:0]    x669_out,                     
			output   [width-1:0]    x670_out,                     
			output   [width-1:0]    x671_out,                     
			output   [width-1:0]    x672_out,                     
			output   [width-1:0]    x673_out,                     
			output   [width-1:0]    x674_out,                     
			output   [width-1:0]    x675_out,                     
			output   [width-1:0]    x676_out,                     
			output   [width-1:0]    x677_out,                     
			output   [width-1:0]    x678_out,                     
			output   [width-1:0]    x679_out,                     
			output   [width-1:0]    x680_out,                     
			output   [width-1:0]    x681_out,                     
			output   [width-1:0]    x682_out,                     
			output   [width-1:0]    x683_out,                     
			output   [width-1:0]    x684_out,                     
			output   [width-1:0]    x685_out,                     
			output   [width-1:0]    x686_out,                     
			output   [width-1:0]    x687_out,                     
			output   [width-1:0]    x688_out,                     
			output   [width-1:0]    x689_out,                     
			output   [width-1:0]    x690_out,                     
			output   [width-1:0]    x691_out,                     
			output   [width-1:0]    x692_out,                     
			output   [width-1:0]    x693_out,                     
			output   [width-1:0]    x694_out,                     
			output   [width-1:0]    x695_out,                     
			output   [width-1:0]    x696_out,                     
			output   [width-1:0]    x697_out,                     
			output   [width-1:0]    x698_out,                     
			output   [width-1:0]    x699_out,                     
			output   [width-1:0]    x700_out,                     
			output   [width-1:0]    x701_out,                     
			output   [width-1:0]    x702_out,                     
			output   [width-1:0]    x703_out,                     
			output   [width-1:0]    x704_out,                     
			output   [width-1:0]    x705_out,                     
			output   [width-1:0]    x706_out,                     
			output   [width-1:0]    x707_out,                     
			output   [width-1:0]    x708_out,                     
			output   [width-1:0]    x709_out,                     
			output   [width-1:0]    x710_out,                     
			output   [width-1:0]    x711_out,                     
			output   [width-1:0]    x712_out,                     
			output   [width-1:0]    x713_out,                     
			output   [width-1:0]    x714_out,                     
			output   [width-1:0]    x715_out,                     
			output   [width-1:0]    x716_out,                     
			output   [width-1:0]    x717_out,                     
			output   [width-1:0]    x718_out,                     
			output   [width-1:0]    x719_out,                     
			output   [width-1:0]    x720_out,                     
			output   [width-1:0]    x721_out,                     
			output   [width-1:0]    x722_out,                     
			output   [width-1:0]    x723_out,                     
			output   [width-1:0]    x724_out,                     
			output   [width-1:0]    x725_out,                     
			output   [width-1:0]    x726_out,                     
			output   [width-1:0]    x727_out,                     
			output   [width-1:0]    x728_out,                     
			output   [width-1:0]    x729_out,                     
			output   [width-1:0]    x730_out,                     
			output   [width-1:0]    x731_out,                     
			output   [width-1:0]    x732_out,                     
			output   [width-1:0]    x733_out,                     
			output   [width-1:0]    x734_out,                     
			output   [width-1:0]    x735_out,                     
			output   [width-1:0]    x736_out,                     
			output   [width-1:0]    x737_out,                     
			output   [width-1:0]    x738_out,                     
			output   [width-1:0]    x739_out,                     
			output   [width-1:0]    x740_out,                     
			output   [width-1:0]    x741_out,                     
			output   [width-1:0]    x742_out,                     
			output   [width-1:0]    x743_out,                     
			output   [width-1:0]    x744_out,                     
			output   [width-1:0]    x745_out,                     
			output   [width-1:0]    x746_out,                     
			output   [width-1:0]    x747_out,                     
			output   [width-1:0]    x748_out,                     
			output   [width-1:0]    x749_out,                     
			output   [width-1:0]    x750_out,                     
			output   [width-1:0]    x751_out,                     
			output   [width-1:0]    x752_out,                     
			output   [width-1:0]    x753_out,                     
			output   [width-1:0]    x754_out,                     
			output   [width-1:0]    x755_out,                     
			output   [width-1:0]    x756_out,                     
			output   [width-1:0]    x757_out,                     
			output   [width-1:0]    x758_out,                     
			output   [width-1:0]    x759_out,                     
			output   [width-1:0]    x760_out,                     
			output   [width-1:0]    x761_out,                     
			output   [width-1:0]    x762_out,                     
			output   [width-1:0]    x763_out,                     
			output   [width-1:0]    x764_out,                     
			output   [width-1:0]    x765_out,                     
			output   [width-1:0]    x766_out,                     
			output   [width-1:0]    x767_out,                     
			output   [width-1:0]    x768_out,                     
			output   [width-1:0]    x769_out,                     
			output   [width-1:0]    x770_out,                     
			output   [width-1:0]    x771_out,                     
			output   [width-1:0]    x772_out,                     
			output   [width-1:0]    x773_out,                     
			output   [width-1:0]    x774_out,                     
			output   [width-1:0]    x775_out,                     
			output   [width-1:0]    x776_out,                     
			output   [width-1:0]    x777_out,                     
			output   [width-1:0]    x778_out,                     
			output   [width-1:0]    x779_out,                     
			output   [width-1:0]    x780_out,                     
			output   [width-1:0]    x781_out,                     
			output   [width-1:0]    x782_out,                     
			output   [width-1:0]    x783_out,                     
			output   [width-1:0]    x784_out,                     
			output   [width-1:0]    x785_out,                     
			output   [width-1:0]    x786_out,                     
			output   [width-1:0]    x787_out,                     
			output   [width-1:0]    x788_out,                     
			output   [width-1:0]    x789_out,                     
			output   [width-1:0]    x790_out,                     
			output   [width-1:0]    x791_out,                     
			output   [width-1:0]    x792_out,                     
			output   [width-1:0]    x793_out,                     
			output   [width-1:0]    x794_out,                     
			output   [width-1:0]    x795_out,                     
			output   [width-1:0]    x796_out,                     
			output   [width-1:0]    x797_out,                     
			output   [width-1:0]    x798_out,                     
			output   [width-1:0]    x799_out,                     
			output   [width-1:0]    x800_out,                     
			output   [width-1:0]    x801_out,                     
			output   [width-1:0]    x802_out,                     
			output   [width-1:0]    x803_out,                     
			output   [width-1:0]    x804_out,                     
			output   [width-1:0]    x805_out,                     
			output   [width-1:0]    x806_out,                     
			output   [width-1:0]    x807_out,                     
			output   [width-1:0]    x808_out,                     
			output   [width-1:0]    x809_out,                     
			output   [width-1:0]    x810_out,                     
			output   [width-1:0]    x811_out,                     
			output   [width-1:0]    x812_out,                     
			output   [width-1:0]    x813_out,                     
			output   [width-1:0]    x814_out,                     
			output   [width-1:0]    x815_out,                     
			output   [width-1:0]    x816_out,                     
			output   [width-1:0]    x817_out,                     
			output   [width-1:0]    x818_out,                     
			output   [width-1:0]    x819_out,                     
			output   [width-1:0]    x820_out,                     
			output   [width-1:0]    x821_out,                     
			output   [width-1:0]    x822_out,                     
			output   [width-1:0]    x823_out,                     
			output   [width-1:0]    x824_out,                     
			output   [width-1:0]    x825_out,                     
			output   [width-1:0]    x826_out,                     
			output   [width-1:0]    x827_out,                     
			output   [width-1:0]    x828_out,                     
			output   [width-1:0]    x829_out,                     
			output   [width-1:0]    x830_out,                     
			output   [width-1:0]    x831_out,                     
			output   [width-1:0]    x832_out,                     
			output   [width-1:0]    x833_out,                     
			output   [width-1:0]    x834_out,                     
			output   [width-1:0]    x835_out,                     
			output   [width-1:0]    x836_out,                     
			output   [width-1:0]    x837_out,                     
			output   [width-1:0]    x838_out,                     
			output   [width-1:0]    x839_out,                     
			output   [width-1:0]    x840_out,                     
			output   [width-1:0]    x841_out,                     
			output   [width-1:0]    x842_out,                     
			output   [width-1:0]    x843_out,                     
			output   [width-1:0]    x844_out,                     
			output   [width-1:0]    x845_out,                     
			output   [width-1:0]    x846_out,                     
			output   [width-1:0]    x847_out,                     
			output   [width-1:0]    x848_out,                     
			output   [width-1:0]    x849_out,                     
			output   [width-1:0]    x850_out,                     
			output   [width-1:0]    x851_out,                     
			output   [width-1:0]    x852_out,                     
			output   [width-1:0]    x853_out,                     
			output   [width-1:0]    x854_out,                     
			output   [width-1:0]    x855_out,                     
			output   [width-1:0]    x856_out,                     
			output   [width-1:0]    x857_out,                     
			output   [width-1:0]    x858_out,                     
			output   [width-1:0]    x859_out,                     
			output   [width-1:0]    x860_out,                     
			output   [width-1:0]    x861_out,                     
			output   [width-1:0]    x862_out,                     
			output   [width-1:0]    x863_out,                     
			output   [width-1:0]    x864_out,                     
			output   [width-1:0]    x865_out,                     
			output   [width-1:0]    x866_out,                     
			output   [width-1:0]    x867_out,                     
			output   [width-1:0]    x868_out,                     
			output   [width-1:0]    x869_out,                     
			output   [width-1:0]    x870_out,                     
			output   [width-1:0]    x871_out,                     
			output   [width-1:0]    x872_out,                     
			output   [width-1:0]    x873_out,                     
			output   [width-1:0]    x874_out,                     
			output   [width-1:0]    x875_out,                     
			output   [width-1:0]    x876_out,                     
			output   [width-1:0]    x877_out,                     
			output   [width-1:0]    x878_out,                     
			output   [width-1:0]    x879_out,                     
			output   [width-1:0]    x880_out,                     
			output   [width-1:0]    x881_out,                     
			output   [width-1:0]    x882_out,                     
			output   [width-1:0]    x883_out,                     
			output   [width-1:0]    x884_out,                     
			output   [width-1:0]    x885_out,                     
			output   [width-1:0]    x886_out,                     
			output   [width-1:0]    x887_out,                     
			output   [width-1:0]    x888_out,                     
			output   [width-1:0]    x889_out,                     
			output   [width-1:0]    x890_out,                     
			output   [width-1:0]    x891_out,                     
			output   [width-1:0]    x892_out,                     
			output   [width-1:0]    x893_out,                     
			output   [width-1:0]    x894_out,                     
			output   [width-1:0]    x895_out,                     
			output   [width-1:0]    x896_out,                     
			output   [width-1:0]    x897_out,                     
			output   [width-1:0]    x898_out,                     
			output   [width-1:0]    x899_out,                     
			output   [width-1:0]    x900_out,                     
			output   [width-1:0]    x901_out,                     
			output   [width-1:0]    x902_out,                     
			output   [width-1:0]    x903_out,                     
			output   [width-1:0]    x904_out,                     
			output   [width-1:0]    x905_out,                     
			output   [width-1:0]    x906_out,                     
			output   [width-1:0]    x907_out,                     
			output   [width-1:0]    x908_out,                     
			output   [width-1:0]    x909_out,                     
			output   [width-1:0]    x910_out,                     
			output   [width-1:0]    x911_out,                     
			output   [width-1:0]    x912_out,                     
			output   [width-1:0]    x913_out,                     
			output   [width-1:0]    x914_out,                     
			output   [width-1:0]    x915_out,                     
			output   [width-1:0]    x916_out,                     
			output   [width-1:0]    x917_out,                     
			output   [width-1:0]    x918_out,                     
			output   [width-1:0]    x919_out,                     
			output   [width-1:0]    x920_out,                     
			output   [width-1:0]    x921_out,                     
			output   [width-1:0]    x922_out,                     
			output   [width-1:0]    x923_out,                     
			output   [width-1:0]    x924_out,                     
			output   [width-1:0]    x925_out,                     
			output   [width-1:0]    x926_out,                     
			output   [width-1:0]    x927_out,                     
			output   [width-1:0]    x928_out,                     
			output   [width-1:0]    x929_out,                     
			output   [width-1:0]    x930_out,                     
			output   [width-1:0]    x931_out,                     
			output   [width-1:0]    x932_out,                     
			output   [width-1:0]    x933_out,                     
			output   [width-1:0]    x934_out,                     
			output   [width-1:0]    x935_out,                     
			output   [width-1:0]    x936_out,                     
			output   [width-1:0]    x937_out,                     
			output   [width-1:0]    x938_out,                     
			output   [width-1:0]    x939_out,                     
			output   [width-1:0]    x940_out,                     
			output   [width-1:0]    x941_out,                     
			output   [width-1:0]    x942_out,                     
			output   [width-1:0]    x943_out,                     
			output   [width-1:0]    x944_out,                     
			output   [width-1:0]    x945_out,                     
			output   [width-1:0]    x946_out,                     
			output   [width-1:0]    x947_out,                     
			output   [width-1:0]    x948_out,                     
			output   [width-1:0]    x949_out,                     
			output   [width-1:0]    x950_out,                     
			output   [width-1:0]    x951_out,                     
			output   [width-1:0]    x952_out,                     
			output   [width-1:0]    x953_out,                     
			output   [width-1:0]    x954_out,                     
			output   [width-1:0]    x955_out,                     
			output   [width-1:0]    x956_out,                     
			output   [width-1:0]    x957_out,                     
			output   [width-1:0]    x958_out,                     
			output   [width-1:0]    x959_out,                     
			output   [width-1:0]    x960_out,                     
			output   [width-1:0]    x961_out,                     
			output   [width-1:0]    x962_out,                     
			output   [width-1:0]    x963_out,                     
			output   [width-1:0]    x964_out,                     
			output   [width-1:0]    x965_out,                     
			output   [width-1:0]    x966_out,                     
			output   [width-1:0]    x967_out,                     
			output   [width-1:0]    x968_out,                     
			output   [width-1:0]    x969_out,                     
			output   [width-1:0]    x970_out,                     
			output   [width-1:0]    x971_out,                     
			output   [width-1:0]    x972_out,                     
			output   [width-1:0]    x973_out,                     
			output   [width-1:0]    x974_out,                     
			output   [width-1:0]    x975_out,                     
			output   [width-1:0]    x976_out,                     
			output   [width-1:0]    x977_out,                     
			output   [width-1:0]    x978_out,                     
			output   [width-1:0]    x979_out,                     
			output   [width-1:0]    x980_out,                     
			output   [width-1:0]    x981_out,                     
			output   [width-1:0]    x982_out,                     
			output   [width-1:0]    x983_out,                     
			output   [width-1:0]    x984_out,                     
			output   [width-1:0]    x985_out,                     
			output   [width-1:0]    x986_out,                     
			output   [width-1:0]    x987_out,                     
			output   [width-1:0]    x988_out,                     
			output   [width-1:0]    x989_out,                     
			output   [width-1:0]    x990_out,                     
			output   [width-1:0]    x991_out,                     
			output   [width-1:0]    x992_out,                     
			output   [width-1:0]    x993_out,                     
			output   [width-1:0]    x994_out,                     
			output   [width-1:0]    x995_out,                     
			output   [width-1:0]    x996_out,                     
			output   [width-1:0]    x997_out,                     
			output   [width-1:0]    x998_out,                     
			output   [width-1:0]    x999_out,                     
			output   [width-1:0]    x1000_out,                    
			output   [width-1:0]    x1001_out,                    
			output   [width-1:0]    x1002_out,                    
			output   [width-1:0]    x1003_out,                    
			output   [width-1:0]    x1004_out,                    
			output   [width-1:0]    x1005_out,                    
			output   [width-1:0]    x1006_out,                    
			output   [width-1:0]    x1007_out,                    
			output   [width-1:0]    x1008_out,                    
			output   [width-1:0]    x1009_out,                    
			output   [width-1:0]    x1010_out,                    
			output   [width-1:0]    x1011_out,                    
			output   [width-1:0]    x1012_out,                    
			output   [width-1:0]    x1013_out,                    
			output   [width-1:0]    x1014_out,                    
			output   [width-1:0]    x1015_out,                    
			output   [width-1:0]    x1016_out,                    
			output   [width-1:0]    x1017_out,                    
			output   [width-1:0]    x1018_out,                    
			output   [width-1:0]    x1019_out,                    
			output   [width-1:0]    x1020_out,                    
			output   [width-1:0]    x1021_out,                    
			output   [width-1:0]    x1022_out,                    
			output   [width-1:0]    x1023_out                     
);

		//--- signal definition
			wire  [width-1:0]        coef[size-1:0];

			reg   [width-1:0]        a0_wr[size-1:0];
			wire  [width-1:0]        a1_wr[size-1:0];
			wire  [width-1:0]        a2_wr[size-1:0];
			wire  [width-1:0]        a3_wr[size-1:0];
			wire  [width-1:0]        a4_wr[size-1:0];
			wire  [width-1:0]        a5_wr[size-1:0];
			wire  [width-1:0]        a6_wr[size-1:0];
			wire  [width-1:0]        a7_wr[size-1:0];
			wire  [width-1:0]        a8_wr[size-1:0];
			wire  [width-1:0]        a9_wr[size-1:0];
			wire  [width-1:0]        a10_wr[size-1:0];
			wire                     comb_stall;

		//--- cofficient assignment
			assign coef[0] =    {12'b011111111111, 12'b000000000000};
			assign coef[1] =    {12'b011111111111, 12'b111111110011};
			assign coef[2] =    {12'b011111111111, 12'b111111100111};
			assign coef[3] =    {12'b011111111111, 12'b111111011010};
			assign coef[4] =    {12'b011111111110, 12'b111111001110};
			assign coef[5] =    {12'b011111111110, 12'b111111000001};
			assign coef[6] =    {12'b011111111110, 12'b111110110101};
			assign coef[7] =    {12'b011111111101, 12'b111110101000};
			assign coef[8] =    {12'b011111111101, 12'b111110011100};
			assign coef[9] =    {12'b011111111100, 12'b111110001111};
			assign coef[10] =   {12'b011111111011, 12'b111110000010};
			assign coef[11] =   {12'b011111111010, 12'b111101110110};
			assign coef[12] =   {12'b011111111010, 12'b111101101001};
			assign coef[13] =   {12'b011111111001, 12'b111101011101};
			assign coef[14] =   {12'b011111111000, 12'b111101010000};
			assign coef[15] =   {12'b011111110110, 12'b111101000100};
			assign coef[16] =   {12'b011111110101, 12'b111100110111};
			assign coef[17] =   {12'b011111110100, 12'b111100101011};
			assign coef[18] =   {12'b011111110011, 12'b111100011110};
			assign coef[19] =   {12'b011111110001, 12'b111100010010};
			assign coef[20] =   {12'b011111110000, 12'b111100000101};
			assign coef[21] =   {12'b011111101110, 12'b111011111001};
			assign coef[22] =   {12'b011111101100, 12'b111011101100};
			assign coef[23] =   {12'b011111101011, 12'b111011100000};
			assign coef[24] =   {12'b011111101001, 12'b111011010100};
			assign coef[25] =   {12'b011111100111, 12'b111011000111};
			assign coef[26] =   {12'b011111100101, 12'b111010111011};
			assign coef[27] =   {12'b011111100011, 12'b111010101110};
			assign coef[28] =   {12'b011111100001, 12'b111010100010};
			assign coef[29] =   {12'b011111011111, 12'b111010010110};
			assign coef[30] =   {12'b011111011100, 12'b111010001001};
			assign coef[31] =   {12'b011111011010, 12'b111001111101};
			assign coef[32] =   {12'b011111011000, 12'b111001110001};
			assign coef[33] =   {12'b011111010101, 12'b111001100100};
			assign coef[34] =   {12'b011111010011, 12'b111001011000};
			assign coef[35] =   {12'b011111010000, 12'b111001001100};
			assign coef[36] =   {12'b011111001101, 12'b111000111111};
			assign coef[37] =   {12'b011111001011, 12'b111000110011};
			assign coef[38] =   {12'b011111001000, 12'b111000100111};
			assign coef[39] =   {12'b011111000101, 12'b111000011011};
			assign coef[40] =   {12'b011111000010, 12'b111000001111};
			assign coef[41] =   {12'b011110111111, 12'b111000000010};
			assign coef[42] =   {12'b011110111011, 12'b110111110110};
			assign coef[43] =   {12'b011110111000, 12'b110111101010};
			assign coef[44] =   {12'b011110110101, 12'b110111011110};
			assign coef[45] =   {12'b011110110010, 12'b110111010010};
			assign coef[46] =   {12'b011110101110, 12'b110111000110};
			assign coef[47] =   {12'b011110101011, 12'b110110111010};
			assign coef[48] =   {12'b011110100111, 12'b110110101110};
			assign coef[49] =   {12'b011110100011, 12'b110110100010};
			assign coef[50] =   {12'b011110011111, 12'b110110010110};
			assign coef[51] =   {12'b011110011100, 12'b110110001010};
			assign coef[52] =   {12'b011110011000, 12'b110101111110};
			assign coef[53] =   {12'b011110010100, 12'b110101110010};
			assign coef[54] =   {12'b011110010000, 12'b110101100110};
			assign coef[55] =   {12'b011110001100, 12'b110101011010};
			assign coef[56] =   {12'b011110000111, 12'b110101001110};
			assign coef[57] =   {12'b011110000011, 12'b110101000011};
			assign coef[58] =   {12'b011101111111, 12'b110100110111};
			assign coef[59] =   {12'b011101111010, 12'b110100101011};
			assign coef[60] =   {12'b011101110110, 12'b110100011111};
			assign coef[61] =   {12'b011101110001, 12'b110100010100};
			assign coef[62] =   {12'b011101101101, 12'b110100001000};
			assign coef[63] =   {12'b011101101000, 12'b110011111100};
			assign coef[64] =   {12'b011101100011, 12'b110011110001};
			assign coef[65] =   {12'b011101011110, 12'b110011100101};
			assign coef[66] =   {12'b011101011001, 12'b110011011001};
			assign coef[67] =   {12'b011101010100, 12'b110011001110};
			assign coef[68] =   {12'b011101001111, 12'b110011000010};
			assign coef[69] =   {12'b011101001010, 12'b110010110111};
			assign coef[70] =   {12'b011101000101, 12'b110010101100};
			assign coef[71] =   {12'b011101000000, 12'b110010100000};
			assign coef[72] =   {12'b011100111011, 12'b110010010101};
			assign coef[73] =   {12'b011100110101, 12'b110010001001};
			assign coef[74] =   {12'b011100110000, 12'b110001111110};
			assign coef[75] =   {12'b011100101010, 12'b110001110011};
			assign coef[76] =   {12'b011100100100, 12'b110001101000};
			assign coef[77] =   {12'b011100011111, 12'b110001011100};
			assign coef[78] =   {12'b011100011001, 12'b110001010001};
			assign coef[79] =   {12'b011100010011, 12'b110001000110};
			assign coef[80] =   {12'b011100001101, 12'b110000111011};
			assign coef[81] =   {12'b011100000111, 12'b110000110000};
			assign coef[82] =   {12'b011100000001, 12'b110000100101};
			assign coef[83] =   {12'b011011111011, 12'b110000011010};
			assign coef[84] =   {12'b011011110101, 12'b110000001111};
			assign coef[85] =   {12'b011011101111, 12'b110000000100};
			assign coef[86] =   {12'b011011101001, 12'b101111111001};
			assign coef[87] =   {12'b011011100010, 12'b101111101110};
			assign coef[88] =   {12'b011011011100, 12'b101111100100};
			assign coef[89] =   {12'b011011010101, 12'b101111011001};
			assign coef[90] =   {12'b011011001111, 12'b101111001110};
			assign coef[91] =   {12'b011011001000, 12'b101111000011};
			assign coef[92] =   {12'b011011000001, 12'b101110111001};
			assign coef[93] =   {12'b011010111011, 12'b101110101110};
			assign coef[94] =   {12'b011010110100, 12'b101110100100};
			assign coef[95] =   {12'b011010101101, 12'b101110011001};
			assign coef[96] =   {12'b011010100110, 12'b101110001111};
			assign coef[97] =   {12'b011010011111, 12'b101110000100};
			assign coef[98] =   {12'b011010011000, 12'b101101111010};
			assign coef[99] =   {12'b011010010001, 12'b101101110000};
			assign coef[100] =  {12'b011010001010, 12'b101101100101};
			assign coef[101] =  {12'b011010000010, 12'b101101011011};
			assign coef[102] =  {12'b011001111011, 12'b101101010001};
			assign coef[103] =  {12'b011001110100, 12'b101101000111};
			assign coef[104] =  {12'b011001101100, 12'b101100111101};
			assign coef[105] =  {12'b011001100101, 12'b101100110010};
			assign coef[106] =  {12'b011001011101, 12'b101100101000};
			assign coef[107] =  {12'b011001010101, 12'b101100011110};
			assign coef[108] =  {12'b011001001110, 12'b101100010101};
			assign coef[109] =  {12'b011001000110, 12'b101100001011};
			assign coef[110] =  {12'b011000111110, 12'b101100000001};
			assign coef[111] =  {12'b011000110110, 12'b101011110111};
			assign coef[112] =  {12'b011000101110, 12'b101011101101};
			assign coef[113] =  {12'b011000100110, 12'b101011100100};
			assign coef[114] =  {12'b011000011110, 12'b101011011010};
			assign coef[115] =  {12'b011000010110, 12'b101011010000};
			assign coef[116] =  {12'b011000001110, 12'b101011000111};
			assign coef[117] =  {12'b011000000110, 12'b101010111101};
			assign coef[118] =  {12'b010111111110, 12'b101010110100};
			assign coef[119] =  {12'b010111110101, 12'b101010101011};
			assign coef[120] =  {12'b010111101101, 12'b101010100001};
			assign coef[121] =  {12'b010111100100, 12'b101010011000};
			assign coef[122] =  {12'b010111011100, 12'b101010001111};
			assign coef[123] =  {12'b010111010011, 12'b101010000110};
			assign coef[124] =  {12'b010111001011, 12'b101001111100};
			assign coef[125] =  {12'b010111000010, 12'b101001110011};
			assign coef[126] =  {12'b010110111001, 12'b101001101010};
			assign coef[127] =  {12'b010110110000, 12'b101001100001};
			assign coef[128] =  {12'b010110100111, 12'b101001011001};
			assign coef[129] =  {12'b010110011111, 12'b101001010000};
			assign coef[130] =  {12'b010110010110, 12'b101001000111};
			assign coef[131] =  {12'b010110001101, 12'b101000111110};
			assign coef[132] =  {12'b010110000100, 12'b101000110101};
			assign coef[133] =  {12'b010101111010, 12'b101000101101};
			assign coef[134] =  {12'b010101110001, 12'b101000100100};
			assign coef[135] =  {12'b010101101000, 12'b101000011100};
			assign coef[136] =  {12'b010101011111, 12'b101000010011};
			assign coef[137] =  {12'b010101010101, 12'b101000001011};
			assign coef[138] =  {12'b010101001100, 12'b101000000010};
			assign coef[139] =  {12'b010101000011, 12'b100111111010};
			assign coef[140] =  {12'b010100111001, 12'b100111110010};
			assign coef[141] =  {12'b010100110000, 12'b100111101010};
			assign coef[142] =  {12'b010100100110, 12'b100111100010};
			assign coef[143] =  {12'b010100011100, 12'b100111011010};
			assign coef[144] =  {12'b010100010011, 12'b100111010010};
			assign coef[145] =  {12'b010100001001, 12'b100111001010};
			assign coef[146] =  {12'b010011111111, 12'b100111000010};
			assign coef[147] =  {12'b010011110101, 12'b100110111010};
			assign coef[148] =  {12'b010011101011, 12'b100110110010};
			assign coef[149] =  {12'b010011100010, 12'b100110101011};
			assign coef[150] =  {12'b010011011000, 12'b100110100011};
			assign coef[151] =  {12'b010011001110, 12'b100110011011};
			assign coef[152] =  {12'b010011000011, 12'b100110010100};
			assign coef[153] =  {12'b010010111001, 12'b100110001100};
			assign coef[154] =  {12'b010010101111, 12'b100110000101};
			assign coef[155] =  {12'b010010100101, 12'b100101111110};
			assign coef[156] =  {12'b010010011011, 12'b100101110110};
			assign coef[157] =  {12'b010010010000, 12'b100101101111};
			assign coef[158] =  {12'b010010000110, 12'b100101101000};
			assign coef[159] =  {12'b010001111100, 12'b100101100001};
			assign coef[160] =  {12'b010001110001, 12'b100101011010};
			assign coef[161] =  {12'b010001100111, 12'b100101010011};
			assign coef[162] =  {12'b010001011100, 12'b100101001100};
			assign coef[163] =  {12'b010001010010, 12'b100101000101};
			assign coef[164] =  {12'b010001000111, 12'b100100111111};
			assign coef[165] =  {12'b010000111101, 12'b100100111000};
			assign coef[166] =  {12'b010000110010, 12'b100100110001};
			assign coef[167] =  {12'b010000100111, 12'b100100101011};
			assign coef[168] =  {12'b010000011100, 12'b100100100100};
			assign coef[169] =  {12'b010000010010, 12'b100100011110};
			assign coef[170] =  {12'b010000000111, 12'b100100010111};
			assign coef[171] =  {12'b001111111100, 12'b100100010001};
			assign coef[172] =  {12'b001111110001, 12'b100100001011};
			assign coef[173] =  {12'b001111100110, 12'b100100000101};
			assign coef[174] =  {12'b001111011011, 12'b100011111111};
			assign coef[175] =  {12'b001111010000, 12'b100011111001};
			assign coef[176] =  {12'b001111000101, 12'b100011110011};
			assign coef[177] =  {12'b001110111010, 12'b100011101101};
			assign coef[178] =  {12'b001110101111, 12'b100011100111};
			assign coef[179] =  {12'b001110100100, 12'b100011100001};
			assign coef[180] =  {12'b001110011000, 12'b100011011100};
			assign coef[181] =  {12'b001110001101, 12'b100011010110};
			assign coef[182] =  {12'b001110000010, 12'b100011010000};
			assign coef[183] =  {12'b001101110111, 12'b100011001011};
			assign coef[184] =  {12'b001101101011, 12'b100011000101};
			assign coef[185] =  {12'b001101100000, 12'b100011000000};
			assign coef[186] =  {12'b001101010100, 12'b100010111011};
			assign coef[187] =  {12'b001101001001, 12'b100010110110};
			assign coef[188] =  {12'b001100111110, 12'b100010110001};
			assign coef[189] =  {12'b001100110010, 12'b100010101100};
			assign coef[190] =  {12'b001100100111, 12'b100010100111};
			assign coef[191] =  {12'b001100011011, 12'b100010100010};
			assign coef[192] =  {12'b001100001111, 12'b100010011101};
			assign coef[193] =  {12'b001100000100, 12'b100010011000};
			assign coef[194] =  {12'b001011111000, 12'b100010010011};
			assign coef[195] =  {12'b001011101100, 12'b100010001111};
			assign coef[196] =  {12'b001011100001, 12'b100010001010};
			assign coef[197] =  {12'b001011010101, 12'b100010000110};
			assign coef[198] =  {12'b001011001001, 12'b100010000001};
			assign coef[199] =  {12'b001010111101, 12'b100001111101};
			assign coef[200] =  {12'b001010110010, 12'b100001111001};
			assign coef[201] =  {12'b001010100110, 12'b100001110100};
			assign coef[202] =  {12'b001010011010, 12'b100001110000};
			assign coef[203] =  {12'b001010001110, 12'b100001101100};
			assign coef[204] =  {12'b001010000010, 12'b100001101000};
			assign coef[205] =  {12'b001001110110, 12'b100001100100};
			assign coef[206] =  {12'b001001101010, 12'b100001100001};
			assign coef[207] =  {12'b001001011110, 12'b100001011101};
			assign coef[208] =  {12'b001001010010, 12'b100001011001};
			assign coef[209] =  {12'b001001000110, 12'b100001010101};
			assign coef[210] =  {12'b001000111010, 12'b100001010010};
			assign coef[211] =  {12'b001000101110, 12'b100001001110};
			assign coef[212] =  {12'b001000100010, 12'b100001001011};
			assign coef[213] =  {12'b001000010110, 12'b100001001000};
			assign coef[214] =  {12'b001000001010, 12'b100001000101};
			assign coef[215] =  {12'b000111111110, 12'b100001000001};
			assign coef[216] =  {12'b000111110001, 12'b100000111110};
			assign coef[217] =  {12'b000111100101, 12'b100000111011};
			assign coef[218] =  {12'b000111011001, 12'b100000111000};
			assign coef[219] =  {12'b000111001101, 12'b100000110101};
			assign coef[220] =  {12'b000111000001, 12'b100000110011};
			assign coef[221] =  {12'b000110110100, 12'b100000110000};
			assign coef[222] =  {12'b000110101000, 12'b100000101101};
			assign coef[223] =  {12'b000110011100, 12'b100000101011};
			assign coef[224] =  {12'b000110001111, 12'b100000101000};
			assign coef[225] =  {12'b000110000011, 12'b100000100110};
			assign coef[226] =  {12'b000101110111, 12'b100000100100};
			assign coef[227] =  {12'b000101101010, 12'b100000100001};
			assign coef[228] =  {12'b000101011110, 12'b100000011111};
			assign coef[229] =  {12'b000101010010, 12'b100000011101};
			assign coef[230] =  {12'b000101000101, 12'b100000011011};
			assign coef[231] =  {12'b000100111001, 12'b100000011001};
			assign coef[232] =  {12'b000100101100, 12'b100000010111};
			assign coef[233] =  {12'b000100100000, 12'b100000010101};
			assign coef[234] =  {12'b000100010100, 12'b100000010100};
			assign coef[235] =  {12'b000100000111, 12'b100000010010};
			assign coef[236] =  {12'b000011111011, 12'b100000010000};
			assign coef[237] =  {12'b000011101110, 12'b100000001111};
			assign coef[238] =  {12'b000011100010, 12'b100000001101};
			assign coef[239] =  {12'b000011010101, 12'b100000001100};
			assign coef[240] =  {12'b000011001001, 12'b100000001011};
			assign coef[241] =  {12'b000010111100, 12'b100000001010};
			assign coef[242] =  {12'b000010110000, 12'b100000001000};
			assign coef[243] =  {12'b000010100011, 12'b100000000111};
			assign coef[244] =  {12'b000010010111, 12'b100000000110};
			assign coef[245] =  {12'b000010001010, 12'b100000000110};
			assign coef[246] =  {12'b000001111110, 12'b100000000101};
			assign coef[247] =  {12'b000001110001, 12'b100000000100};
			assign coef[248] =  {12'b000001100100, 12'b100000000011};
			assign coef[249] =  {12'b000001011000, 12'b100000000011};
			assign coef[250] =  {12'b000001001011, 12'b100000000010};
			assign coef[251] =  {12'b000000111111, 12'b100000000010};
			assign coef[252] =  {12'b000000110010, 12'b100000000010};
			assign coef[253] =  {12'b000000100110, 12'b100000000001};
			assign coef[254] =  {12'b000000011001, 12'b100000000001};
			assign coef[255] =  {12'b000000001101, 12'b100000000001};
			assign coef[256] =  {12'b000000000000, 12'b100000000001};
			assign coef[257] =  {12'b111111110011, 12'b100000000001};
			assign coef[258] =  {12'b111111100111, 12'b100000000001};
			assign coef[259] =  {12'b111111011010, 12'b100000000001};
			assign coef[260] =  {12'b111111001110, 12'b100000000010};
			assign coef[261] =  {12'b111111000001, 12'b100000000010};
			assign coef[262] =  {12'b111110110101, 12'b100000000010};
			assign coef[263] =  {12'b111110101000, 12'b100000000011};
			assign coef[264] =  {12'b111110011100, 12'b100000000011};
			assign coef[265] =  {12'b111110001111, 12'b100000000100};
			assign coef[266] =  {12'b111110000010, 12'b100000000101};
			assign coef[267] =  {12'b111101110110, 12'b100000000110};
			assign coef[268] =  {12'b111101101001, 12'b100000000110};
			assign coef[269] =  {12'b111101011101, 12'b100000000111};
			assign coef[270] =  {12'b111101010000, 12'b100000001000};
			assign coef[271] =  {12'b111101000100, 12'b100000001010};
			assign coef[272] =  {12'b111100110111, 12'b100000001011};
			assign coef[273] =  {12'b111100101011, 12'b100000001100};
			assign coef[274] =  {12'b111100011110, 12'b100000001101};
			assign coef[275] =  {12'b111100010010, 12'b100000001111};
			assign coef[276] =  {12'b111100000101, 12'b100000010000};
			assign coef[277] =  {12'b111011111001, 12'b100000010010};
			assign coef[278] =  {12'b111011101100, 12'b100000010100};
			assign coef[279] =  {12'b111011100000, 12'b100000010101};
			assign coef[280] =  {12'b111011010100, 12'b100000010111};
			assign coef[281] =  {12'b111011000111, 12'b100000011001};
			assign coef[282] =  {12'b111010111011, 12'b100000011011};
			assign coef[283] =  {12'b111010101110, 12'b100000011101};
			assign coef[284] =  {12'b111010100010, 12'b100000011111};
			assign coef[285] =  {12'b111010010110, 12'b100000100001};
			assign coef[286] =  {12'b111010001001, 12'b100000100100};
			assign coef[287] =  {12'b111001111101, 12'b100000100110};
			assign coef[288] =  {12'b111001110001, 12'b100000101000};
			assign coef[289] =  {12'b111001100100, 12'b100000101011};
			assign coef[290] =  {12'b111001011000, 12'b100000101101};
			assign coef[291] =  {12'b111001001100, 12'b100000110000};
			assign coef[292] =  {12'b111000111111, 12'b100000110011};
			assign coef[293] =  {12'b111000110011, 12'b100000110101};
			assign coef[294] =  {12'b111000100111, 12'b100000111000};
			assign coef[295] =  {12'b111000011011, 12'b100000111011};
			assign coef[296] =  {12'b111000001111, 12'b100000111110};
			assign coef[297] =  {12'b111000000010, 12'b100001000001};
			assign coef[298] =  {12'b110111110110, 12'b100001000101};
			assign coef[299] =  {12'b110111101010, 12'b100001001000};
			assign coef[300] =  {12'b110111011110, 12'b100001001011};
			assign coef[301] =  {12'b110111010010, 12'b100001001110};
			assign coef[302] =  {12'b110111000110, 12'b100001010010};
			assign coef[303] =  {12'b110110111010, 12'b100001010101};
			assign coef[304] =  {12'b110110101110, 12'b100001011001};
			assign coef[305] =  {12'b110110100010, 12'b100001011101};
			assign coef[306] =  {12'b110110010110, 12'b100001100001};
			assign coef[307] =  {12'b110110001010, 12'b100001100100};
			assign coef[308] =  {12'b110101111110, 12'b100001101000};
			assign coef[309] =  {12'b110101110010, 12'b100001101100};
			assign coef[310] =  {12'b110101100110, 12'b100001110000};
			assign coef[311] =  {12'b110101011010, 12'b100001110100};
			assign coef[312] =  {12'b110101001110, 12'b100001111001};
			assign coef[313] =  {12'b110101000011, 12'b100001111101};
			assign coef[314] =  {12'b110100110111, 12'b100010000001};
			assign coef[315] =  {12'b110100101011, 12'b100010000110};
			assign coef[316] =  {12'b110100011111, 12'b100010001010};
			assign coef[317] =  {12'b110100010100, 12'b100010001111};
			assign coef[318] =  {12'b110100001000, 12'b100010010011};
			assign coef[319] =  {12'b110011111100, 12'b100010011000};
			assign coef[320] =  {12'b110011110001, 12'b100010011101};
			assign coef[321] =  {12'b110011100101, 12'b100010100010};
			assign coef[322] =  {12'b110011011001, 12'b100010100111};
			assign coef[323] =  {12'b110011001110, 12'b100010101100};
			assign coef[324] =  {12'b110011000010, 12'b100010110001};
			assign coef[325] =  {12'b110010110111, 12'b100010110110};
			assign coef[326] =  {12'b110010101100, 12'b100010111011};
			assign coef[327] =  {12'b110010100000, 12'b100011000000};
			assign coef[328] =  {12'b110010010101, 12'b100011000101};
			assign coef[329] =  {12'b110010001001, 12'b100011001011};
			assign coef[330] =  {12'b110001111110, 12'b100011010000};
			assign coef[331] =  {12'b110001110011, 12'b100011010110};
			assign coef[332] =  {12'b110001101000, 12'b100011011100};
			assign coef[333] =  {12'b110001011100, 12'b100011100001};
			assign coef[334] =  {12'b110001010001, 12'b100011100111};
			assign coef[335] =  {12'b110001000110, 12'b100011101101};
			assign coef[336] =  {12'b110000111011, 12'b100011110011};
			assign coef[337] =  {12'b110000110000, 12'b100011111001};
			assign coef[338] =  {12'b110000100101, 12'b100011111111};
			assign coef[339] =  {12'b110000011010, 12'b100100000101};
			assign coef[340] =  {12'b110000001111, 12'b100100001011};
			assign coef[341] =  {12'b110000000100, 12'b100100010001};
			assign coef[342] =  {12'b101111111001, 12'b100100010111};
			assign coef[343] =  {12'b101111101110, 12'b100100011110};
			assign coef[344] =  {12'b101111100100, 12'b100100100100};
			assign coef[345] =  {12'b101111011001, 12'b100100101011};
			assign coef[346] =  {12'b101111001110, 12'b100100110001};
			assign coef[347] =  {12'b101111000011, 12'b100100111000};
			assign coef[348] =  {12'b101110111001, 12'b100100111111};
			assign coef[349] =  {12'b101110101110, 12'b100101000101};
			assign coef[350] =  {12'b101110100100, 12'b100101001100};
			assign coef[351] =  {12'b101110011001, 12'b100101010011};
			assign coef[352] =  {12'b101110001111, 12'b100101011010};
			assign coef[353] =  {12'b101110000100, 12'b100101100001};
			assign coef[354] =  {12'b101101111010, 12'b100101101000};
			assign coef[355] =  {12'b101101110000, 12'b100101101111};
			assign coef[356] =  {12'b101101100101, 12'b100101110110};
			assign coef[357] =  {12'b101101011011, 12'b100101111110};
			assign coef[358] =  {12'b101101010001, 12'b100110000101};
			assign coef[359] =  {12'b101101000111, 12'b100110001100};
			assign coef[360] =  {12'b101100111101, 12'b100110010100};
			assign coef[361] =  {12'b101100110010, 12'b100110011011};
			assign coef[362] =  {12'b101100101000, 12'b100110100011};
			assign coef[363] =  {12'b101100011110, 12'b100110101011};
			assign coef[364] =  {12'b101100010101, 12'b100110110010};
			assign coef[365] =  {12'b101100001011, 12'b100110111010};
			assign coef[366] =  {12'b101100000001, 12'b100111000010};
			assign coef[367] =  {12'b101011110111, 12'b100111001010};
			assign coef[368] =  {12'b101011101101, 12'b100111010010};
			assign coef[369] =  {12'b101011100100, 12'b100111011010};
			assign coef[370] =  {12'b101011011010, 12'b100111100010};
			assign coef[371] =  {12'b101011010000, 12'b100111101010};
			assign coef[372] =  {12'b101011000111, 12'b100111110010};
			assign coef[373] =  {12'b101010111101, 12'b100111111010};
			assign coef[374] =  {12'b101010110100, 12'b101000000010};
			assign coef[375] =  {12'b101010101011, 12'b101000001011};
			assign coef[376] =  {12'b101010100001, 12'b101000010011};
			assign coef[377] =  {12'b101010011000, 12'b101000011100};
			assign coef[378] =  {12'b101010001111, 12'b101000100100};
			assign coef[379] =  {12'b101010000110, 12'b101000101101};
			assign coef[380] =  {12'b101001111100, 12'b101000110101};
			assign coef[381] =  {12'b101001110011, 12'b101000111110};
			assign coef[382] =  {12'b101001101010, 12'b101001000111};
			assign coef[383] =  {12'b101001100001, 12'b101001010000};
			assign coef[384] =  {12'b101001011001, 12'b101001011001};
			assign coef[385] =  {12'b101001010000, 12'b101001100001};
			assign coef[386] =  {12'b101001000111, 12'b101001101010};
			assign coef[387] =  {12'b101000111110, 12'b101001110011};
			assign coef[388] =  {12'b101000110101, 12'b101001111100};
			assign coef[389] =  {12'b101000101101, 12'b101010000110};
			assign coef[390] =  {12'b101000100100, 12'b101010001111};
			assign coef[391] =  {12'b101000011100, 12'b101010011000};
			assign coef[392] =  {12'b101000010011, 12'b101010100001};
			assign coef[393] =  {12'b101000001011, 12'b101010101011};
			assign coef[394] =  {12'b101000000010, 12'b101010110100};
			assign coef[395] =  {12'b100111111010, 12'b101010111101};
			assign coef[396] =  {12'b100111110010, 12'b101011000111};
			assign coef[397] =  {12'b100111101010, 12'b101011010000};
			assign coef[398] =  {12'b100111100010, 12'b101011011010};
			assign coef[399] =  {12'b100111011010, 12'b101011100100};
			assign coef[400] =  {12'b100111010010, 12'b101011101101};
			assign coef[401] =  {12'b100111001010, 12'b101011110111};
			assign coef[402] =  {12'b100111000010, 12'b101100000001};
			assign coef[403] =  {12'b100110111010, 12'b101100001011};
			assign coef[404] =  {12'b100110110010, 12'b101100010101};
			assign coef[405] =  {12'b100110101011, 12'b101100011110};
			assign coef[406] =  {12'b100110100011, 12'b101100101000};
			assign coef[407] =  {12'b100110011011, 12'b101100110010};
			assign coef[408] =  {12'b100110010100, 12'b101100111101};
			assign coef[409] =  {12'b100110001100, 12'b101101000111};
			assign coef[410] =  {12'b100110000101, 12'b101101010001};
			assign coef[411] =  {12'b100101111110, 12'b101101011011};
			assign coef[412] =  {12'b100101110110, 12'b101101100101};
			assign coef[413] =  {12'b100101101111, 12'b101101110000};
			assign coef[414] =  {12'b100101101000, 12'b101101111010};
			assign coef[415] =  {12'b100101100001, 12'b101110000100};
			assign coef[416] =  {12'b100101011010, 12'b101110001111};
			assign coef[417] =  {12'b100101010011, 12'b101110011001};
			assign coef[418] =  {12'b100101001100, 12'b101110100100};
			assign coef[419] =  {12'b100101000101, 12'b101110101110};
			assign coef[420] =  {12'b100100111111, 12'b101110111001};
			assign coef[421] =  {12'b100100111000, 12'b101111000011};
			assign coef[422] =  {12'b100100110001, 12'b101111001110};
			assign coef[423] =  {12'b100100101011, 12'b101111011001};
			assign coef[424] =  {12'b100100100100, 12'b101111100100};
			assign coef[425] =  {12'b100100011110, 12'b101111101110};
			assign coef[426] =  {12'b100100010111, 12'b101111111001};
			assign coef[427] =  {12'b100100010001, 12'b110000000100};
			assign coef[428] =  {12'b100100001011, 12'b110000001111};
			assign coef[429] =  {12'b100100000101, 12'b110000011010};
			assign coef[430] =  {12'b100011111111, 12'b110000100101};
			assign coef[431] =  {12'b100011111001, 12'b110000110000};
			assign coef[432] =  {12'b100011110011, 12'b110000111011};
			assign coef[433] =  {12'b100011101101, 12'b110001000110};
			assign coef[434] =  {12'b100011100111, 12'b110001010001};
			assign coef[435] =  {12'b100011100001, 12'b110001011100};
			assign coef[436] =  {12'b100011011100, 12'b110001101000};
			assign coef[437] =  {12'b100011010110, 12'b110001110011};
			assign coef[438] =  {12'b100011010000, 12'b110001111110};
			assign coef[439] =  {12'b100011001011, 12'b110010001001};
			assign coef[440] =  {12'b100011000101, 12'b110010010101};
			assign coef[441] =  {12'b100011000000, 12'b110010100000};
			assign coef[442] =  {12'b100010111011, 12'b110010101100};
			assign coef[443] =  {12'b100010110110, 12'b110010110111};
			assign coef[444] =  {12'b100010110001, 12'b110011000010};
			assign coef[445] =  {12'b100010101100, 12'b110011001110};
			assign coef[446] =  {12'b100010100111, 12'b110011011001};
			assign coef[447] =  {12'b100010100010, 12'b110011100101};
			assign coef[448] =  {12'b100010011101, 12'b110011110001};
			assign coef[449] =  {12'b100010011000, 12'b110011111100};
			assign coef[450] =  {12'b100010010011, 12'b110100001000};
			assign coef[451] =  {12'b100010001111, 12'b110100010100};
			assign coef[452] =  {12'b100010001010, 12'b110100011111};
			assign coef[453] =  {12'b100010000110, 12'b110100101011};
			assign coef[454] =  {12'b100010000001, 12'b110100110111};
			assign coef[455] =  {12'b100001111101, 12'b110101000011};
			assign coef[456] =  {12'b100001111001, 12'b110101001110};
			assign coef[457] =  {12'b100001110100, 12'b110101011010};
			assign coef[458] =  {12'b100001110000, 12'b110101100110};
			assign coef[459] =  {12'b100001101100, 12'b110101110010};
			assign coef[460] =  {12'b100001101000, 12'b110101111110};
			assign coef[461] =  {12'b100001100100, 12'b110110001010};
			assign coef[462] =  {12'b100001100001, 12'b110110010110};
			assign coef[463] =  {12'b100001011101, 12'b110110100010};
			assign coef[464] =  {12'b100001011001, 12'b110110101110};
			assign coef[465] =  {12'b100001010101, 12'b110110111010};
			assign coef[466] =  {12'b100001010010, 12'b110111000110};
			assign coef[467] =  {12'b100001001110, 12'b110111010010};
			assign coef[468] =  {12'b100001001011, 12'b110111011110};
			assign coef[469] =  {12'b100001001000, 12'b110111101010};
			assign coef[470] =  {12'b100001000101, 12'b110111110110};
			assign coef[471] =  {12'b100001000001, 12'b111000000010};
			assign coef[472] =  {12'b100000111110, 12'b111000001111};
			assign coef[473] =  {12'b100000111011, 12'b111000011011};
			assign coef[474] =  {12'b100000111000, 12'b111000100111};
			assign coef[475] =  {12'b100000110101, 12'b111000110011};
			assign coef[476] =  {12'b100000110011, 12'b111000111111};
			assign coef[477] =  {12'b100000110000, 12'b111001001100};
			assign coef[478] =  {12'b100000101101, 12'b111001011000};
			assign coef[479] =  {12'b100000101011, 12'b111001100100};
			assign coef[480] =  {12'b100000101000, 12'b111001110001};
			assign coef[481] =  {12'b100000100110, 12'b111001111101};
			assign coef[482] =  {12'b100000100100, 12'b111010001001};
			assign coef[483] =  {12'b100000100001, 12'b111010010110};
			assign coef[484] =  {12'b100000011111, 12'b111010100010};
			assign coef[485] =  {12'b100000011101, 12'b111010101110};
			assign coef[486] =  {12'b100000011011, 12'b111010111011};
			assign coef[487] =  {12'b100000011001, 12'b111011000111};
			assign coef[488] =  {12'b100000010111, 12'b111011010100};
			assign coef[489] =  {12'b100000010101, 12'b111011100000};
			assign coef[490] =  {12'b100000010100, 12'b111011101100};
			assign coef[491] =  {12'b100000010010, 12'b111011111001};
			assign coef[492] =  {12'b100000010000, 12'b111100000101};
			assign coef[493] =  {12'b100000001111, 12'b111100010010};
			assign coef[494] =  {12'b100000001101, 12'b111100011110};
			assign coef[495] =  {12'b100000001100, 12'b111100101011};
			assign coef[496] =  {12'b100000001011, 12'b111100110111};
			assign coef[497] =  {12'b100000001010, 12'b111101000100};
			assign coef[498] =  {12'b100000001000, 12'b111101010000};
			assign coef[499] =  {12'b100000000111, 12'b111101011101};
			assign coef[500] =  {12'b100000000110, 12'b111101101001};
			assign coef[501] =  {12'b100000000110, 12'b111101110110};
			assign coef[502] =  {12'b100000000101, 12'b111110000010};
			assign coef[503] =  {12'b100000000100, 12'b111110001111};
			assign coef[504] =  {12'b100000000011, 12'b111110011100};
			assign coef[505] =  {12'b100000000011, 12'b111110101000};
			assign coef[506] =  {12'b100000000010, 12'b111110110101};
			assign coef[507] =  {12'b100000000010, 12'b111111000001};
			assign coef[508] =  {12'b100000000010, 12'b111111001110};
			assign coef[509] =  {12'b100000000001, 12'b111111011010};
			assign coef[510] =  {12'b100000000001, 12'b111111100111};
			assign coef[511] =  {12'b100000000001, 12'b111111110011};

		//--- fifo stage
			localparam depth=`LOG2(size);
			fifo #(.depth(depth)) inst_fifo(.clk(clk), .rst(rst), .stall_in(stall), .stall_out(stall_out));

			assign comb_stall = stall_out & stall;

		//--- input stage
			always @(posedge clk or posedge rst) begin
				if (rst) begin
					a0_wr[0]       <= 0;                           
					a0_wr[1]       <= 0;                           
					a0_wr[2]       <= 0;                           
					a0_wr[3]       <= 0;                           
					a0_wr[4]       <= 0;                           
					a0_wr[5]       <= 0;                           
					a0_wr[6]       <= 0;                           
					a0_wr[7]       <= 0;                           
					a0_wr[8]       <= 0;                           
					a0_wr[9]       <= 0;                           
					a0_wr[10]      <= 0;                           
					a0_wr[11]      <= 0;                           
					a0_wr[12]      <= 0;                           
					a0_wr[13]      <= 0;                           
					a0_wr[14]      <= 0;                           
					a0_wr[15]      <= 0;                           
					a0_wr[16]      <= 0;                           
					a0_wr[17]      <= 0;                           
					a0_wr[18]      <= 0;                           
					a0_wr[19]      <= 0;                           
					a0_wr[20]      <= 0;                           
					a0_wr[21]      <= 0;                           
					a0_wr[22]      <= 0;                           
					a0_wr[23]      <= 0;                           
					a0_wr[24]      <= 0;                           
					a0_wr[25]      <= 0;                           
					a0_wr[26]      <= 0;                           
					a0_wr[27]      <= 0;                           
					a0_wr[28]      <= 0;                           
					a0_wr[29]      <= 0;                           
					a0_wr[30]      <= 0;                           
					a0_wr[31]      <= 0;                           
					a0_wr[32]      <= 0;                           
					a0_wr[33]      <= 0;                           
					a0_wr[34]      <= 0;                           
					a0_wr[35]      <= 0;                           
					a0_wr[36]      <= 0;                           
					a0_wr[37]      <= 0;                           
					a0_wr[38]      <= 0;                           
					a0_wr[39]      <= 0;                           
					a0_wr[40]      <= 0;                           
					a0_wr[41]      <= 0;                           
					a0_wr[42]      <= 0;                           
					a0_wr[43]      <= 0;                           
					a0_wr[44]      <= 0;                           
					a0_wr[45]      <= 0;                           
					a0_wr[46]      <= 0;                           
					a0_wr[47]      <= 0;                           
					a0_wr[48]      <= 0;                           
					a0_wr[49]      <= 0;                           
					a0_wr[50]      <= 0;                           
					a0_wr[51]      <= 0;                           
					a0_wr[52]      <= 0;                           
					a0_wr[53]      <= 0;                           
					a0_wr[54]      <= 0;                           
					a0_wr[55]      <= 0;                           
					a0_wr[56]      <= 0;                           
					a0_wr[57]      <= 0;                           
					a0_wr[58]      <= 0;                           
					a0_wr[59]      <= 0;                           
					a0_wr[60]      <= 0;                           
					a0_wr[61]      <= 0;                           
					a0_wr[62]      <= 0;                           
					a0_wr[63]      <= 0;                           
					a0_wr[64]      <= 0;                           
					a0_wr[65]      <= 0;                           
					a0_wr[66]      <= 0;                           
					a0_wr[67]      <= 0;                           
					a0_wr[68]      <= 0;                           
					a0_wr[69]      <= 0;                           
					a0_wr[70]      <= 0;                           
					a0_wr[71]      <= 0;                           
					a0_wr[72]      <= 0;                           
					a0_wr[73]      <= 0;                           
					a0_wr[74]      <= 0;                           
					a0_wr[75]      <= 0;                           
					a0_wr[76]      <= 0;                           
					a0_wr[77]      <= 0;                           
					a0_wr[78]      <= 0;                           
					a0_wr[79]      <= 0;                           
					a0_wr[80]      <= 0;                           
					a0_wr[81]      <= 0;                           
					a0_wr[82]      <= 0;                           
					a0_wr[83]      <= 0;                           
					a0_wr[84]      <= 0;                           
					a0_wr[85]      <= 0;                           
					a0_wr[86]      <= 0;                           
					a0_wr[87]      <= 0;                           
					a0_wr[88]      <= 0;                           
					a0_wr[89]      <= 0;                           
					a0_wr[90]      <= 0;                           
					a0_wr[91]      <= 0;                           
					a0_wr[92]      <= 0;                           
					a0_wr[93]      <= 0;                           
					a0_wr[94]      <= 0;                           
					a0_wr[95]      <= 0;                           
					a0_wr[96]      <= 0;                           
					a0_wr[97]      <= 0;                           
					a0_wr[98]      <= 0;                           
					a0_wr[99]      <= 0;                           
					a0_wr[100]     <= 0;                           
					a0_wr[101]     <= 0;                           
					a0_wr[102]     <= 0;                           
					a0_wr[103]     <= 0;                           
					a0_wr[104]     <= 0;                           
					a0_wr[105]     <= 0;                           
					a0_wr[106]     <= 0;                           
					a0_wr[107]     <= 0;                           
					a0_wr[108]     <= 0;                           
					a0_wr[109]     <= 0;                           
					a0_wr[110]     <= 0;                           
					a0_wr[111]     <= 0;                           
					a0_wr[112]     <= 0;                           
					a0_wr[113]     <= 0;                           
					a0_wr[114]     <= 0;                           
					a0_wr[115]     <= 0;                           
					a0_wr[116]     <= 0;                           
					a0_wr[117]     <= 0;                           
					a0_wr[118]     <= 0;                           
					a0_wr[119]     <= 0;                           
					a0_wr[120]     <= 0;                           
					a0_wr[121]     <= 0;                           
					a0_wr[122]     <= 0;                           
					a0_wr[123]     <= 0;                           
					a0_wr[124]     <= 0;                           
					a0_wr[125]     <= 0;                           
					a0_wr[126]     <= 0;                           
					a0_wr[127]     <= 0;                           
					a0_wr[128]     <= 0;                           
					a0_wr[129]     <= 0;                           
					a0_wr[130]     <= 0;                           
					a0_wr[131]     <= 0;                           
					a0_wr[132]     <= 0;                           
					a0_wr[133]     <= 0;                           
					a0_wr[134]     <= 0;                           
					a0_wr[135]     <= 0;                           
					a0_wr[136]     <= 0;                           
					a0_wr[137]     <= 0;                           
					a0_wr[138]     <= 0;                           
					a0_wr[139]     <= 0;                           
					a0_wr[140]     <= 0;                           
					a0_wr[141]     <= 0;                           
					a0_wr[142]     <= 0;                           
					a0_wr[143]     <= 0;                           
					a0_wr[144]     <= 0;                           
					a0_wr[145]     <= 0;                           
					a0_wr[146]     <= 0;                           
					a0_wr[147]     <= 0;                           
					a0_wr[148]     <= 0;                           
					a0_wr[149]     <= 0;                           
					a0_wr[150]     <= 0;                           
					a0_wr[151]     <= 0;                           
					a0_wr[152]     <= 0;                           
					a0_wr[153]     <= 0;                           
					a0_wr[154]     <= 0;                           
					a0_wr[155]     <= 0;                           
					a0_wr[156]     <= 0;                           
					a0_wr[157]     <= 0;                           
					a0_wr[158]     <= 0;                           
					a0_wr[159]     <= 0;                           
					a0_wr[160]     <= 0;                           
					a0_wr[161]     <= 0;                           
					a0_wr[162]     <= 0;                           
					a0_wr[163]     <= 0;                           
					a0_wr[164]     <= 0;                           
					a0_wr[165]     <= 0;                           
					a0_wr[166]     <= 0;                           
					a0_wr[167]     <= 0;                           
					a0_wr[168]     <= 0;                           
					a0_wr[169]     <= 0;                           
					a0_wr[170]     <= 0;                           
					a0_wr[171]     <= 0;                           
					a0_wr[172]     <= 0;                           
					a0_wr[173]     <= 0;                           
					a0_wr[174]     <= 0;                           
					a0_wr[175]     <= 0;                           
					a0_wr[176]     <= 0;                           
					a0_wr[177]     <= 0;                           
					a0_wr[178]     <= 0;                           
					a0_wr[179]     <= 0;                           
					a0_wr[180]     <= 0;                           
					a0_wr[181]     <= 0;                           
					a0_wr[182]     <= 0;                           
					a0_wr[183]     <= 0;                           
					a0_wr[184]     <= 0;                           
					a0_wr[185]     <= 0;                           
					a0_wr[186]     <= 0;                           
					a0_wr[187]     <= 0;                           
					a0_wr[188]     <= 0;                           
					a0_wr[189]     <= 0;                           
					a0_wr[190]     <= 0;                           
					a0_wr[191]     <= 0;                           
					a0_wr[192]     <= 0;                           
					a0_wr[193]     <= 0;                           
					a0_wr[194]     <= 0;                           
					a0_wr[195]     <= 0;                           
					a0_wr[196]     <= 0;                           
					a0_wr[197]     <= 0;                           
					a0_wr[198]     <= 0;                           
					a0_wr[199]     <= 0;                           
					a0_wr[200]     <= 0;                           
					a0_wr[201]     <= 0;                           
					a0_wr[202]     <= 0;                           
					a0_wr[203]     <= 0;                           
					a0_wr[204]     <= 0;                           
					a0_wr[205]     <= 0;                           
					a0_wr[206]     <= 0;                           
					a0_wr[207]     <= 0;                           
					a0_wr[208]     <= 0;                           
					a0_wr[209]     <= 0;                           
					a0_wr[210]     <= 0;                           
					a0_wr[211]     <= 0;                           
					a0_wr[212]     <= 0;                           
					a0_wr[213]     <= 0;                           
					a0_wr[214]     <= 0;                           
					a0_wr[215]     <= 0;                           
					a0_wr[216]     <= 0;                           
					a0_wr[217]     <= 0;                           
					a0_wr[218]     <= 0;                           
					a0_wr[219]     <= 0;                           
					a0_wr[220]     <= 0;                           
					a0_wr[221]     <= 0;                           
					a0_wr[222]     <= 0;                           
					a0_wr[223]     <= 0;                           
					a0_wr[224]     <= 0;                           
					a0_wr[225]     <= 0;                           
					a0_wr[226]     <= 0;                           
					a0_wr[227]     <= 0;                           
					a0_wr[228]     <= 0;                           
					a0_wr[229]     <= 0;                           
					a0_wr[230]     <= 0;                           
					a0_wr[231]     <= 0;                           
					a0_wr[232]     <= 0;                           
					a0_wr[233]     <= 0;                           
					a0_wr[234]     <= 0;                           
					a0_wr[235]     <= 0;                           
					a0_wr[236]     <= 0;                           
					a0_wr[237]     <= 0;                           
					a0_wr[238]     <= 0;                           
					a0_wr[239]     <= 0;                           
					a0_wr[240]     <= 0;                           
					a0_wr[241]     <= 0;                           
					a0_wr[242]     <= 0;                           
					a0_wr[243]     <= 0;                           
					a0_wr[244]     <= 0;                           
					a0_wr[245]     <= 0;                           
					a0_wr[246]     <= 0;                           
					a0_wr[247]     <= 0;                           
					a0_wr[248]     <= 0;                           
					a0_wr[249]     <= 0;                           
					a0_wr[250]     <= 0;                           
					a0_wr[251]     <= 0;                           
					a0_wr[252]     <= 0;                           
					a0_wr[253]     <= 0;                           
					a0_wr[254]     <= 0;                           
					a0_wr[255]     <= 0;                           
					a0_wr[256]     <= 0;                           
					a0_wr[257]     <= 0;                           
					a0_wr[258]     <= 0;                           
					a0_wr[259]     <= 0;                           
					a0_wr[260]     <= 0;                           
					a0_wr[261]     <= 0;                           
					a0_wr[262]     <= 0;                           
					a0_wr[263]     <= 0;                           
					a0_wr[264]     <= 0;                           
					a0_wr[265]     <= 0;                           
					a0_wr[266]     <= 0;                           
					a0_wr[267]     <= 0;                           
					a0_wr[268]     <= 0;                           
					a0_wr[269]     <= 0;                           
					a0_wr[270]     <= 0;                           
					a0_wr[271]     <= 0;                           
					a0_wr[272]     <= 0;                           
					a0_wr[273]     <= 0;                           
					a0_wr[274]     <= 0;                           
					a0_wr[275]     <= 0;                           
					a0_wr[276]     <= 0;                           
					a0_wr[277]     <= 0;                           
					a0_wr[278]     <= 0;                           
					a0_wr[279]     <= 0;                           
					a0_wr[280]     <= 0;                           
					a0_wr[281]     <= 0;                           
					a0_wr[282]     <= 0;                           
					a0_wr[283]     <= 0;                           
					a0_wr[284]     <= 0;                           
					a0_wr[285]     <= 0;                           
					a0_wr[286]     <= 0;                           
					a0_wr[287]     <= 0;                           
					a0_wr[288]     <= 0;                           
					a0_wr[289]     <= 0;                           
					a0_wr[290]     <= 0;                           
					a0_wr[291]     <= 0;                           
					a0_wr[292]     <= 0;                           
					a0_wr[293]     <= 0;                           
					a0_wr[294]     <= 0;                           
					a0_wr[295]     <= 0;                           
					a0_wr[296]     <= 0;                           
					a0_wr[297]     <= 0;                           
					a0_wr[298]     <= 0;                           
					a0_wr[299]     <= 0;                           
					a0_wr[300]     <= 0;                           
					a0_wr[301]     <= 0;                           
					a0_wr[302]     <= 0;                           
					a0_wr[303]     <= 0;                           
					a0_wr[304]     <= 0;                           
					a0_wr[305]     <= 0;                           
					a0_wr[306]     <= 0;                           
					a0_wr[307]     <= 0;                           
					a0_wr[308]     <= 0;                           
					a0_wr[309]     <= 0;                           
					a0_wr[310]     <= 0;                           
					a0_wr[311]     <= 0;                           
					a0_wr[312]     <= 0;                           
					a0_wr[313]     <= 0;                           
					a0_wr[314]     <= 0;                           
					a0_wr[315]     <= 0;                           
					a0_wr[316]     <= 0;                           
					a0_wr[317]     <= 0;                           
					a0_wr[318]     <= 0;                           
					a0_wr[319]     <= 0;                           
					a0_wr[320]     <= 0;                           
					a0_wr[321]     <= 0;                           
					a0_wr[322]     <= 0;                           
					a0_wr[323]     <= 0;                           
					a0_wr[324]     <= 0;                           
					a0_wr[325]     <= 0;                           
					a0_wr[326]     <= 0;                           
					a0_wr[327]     <= 0;                           
					a0_wr[328]     <= 0;                           
					a0_wr[329]     <= 0;                           
					a0_wr[330]     <= 0;                           
					a0_wr[331]     <= 0;                           
					a0_wr[332]     <= 0;                           
					a0_wr[333]     <= 0;                           
					a0_wr[334]     <= 0;                           
					a0_wr[335]     <= 0;                           
					a0_wr[336]     <= 0;                           
					a0_wr[337]     <= 0;                           
					a0_wr[338]     <= 0;                           
					a0_wr[339]     <= 0;                           
					a0_wr[340]     <= 0;                           
					a0_wr[341]     <= 0;                           
					a0_wr[342]     <= 0;                           
					a0_wr[343]     <= 0;                           
					a0_wr[344]     <= 0;                           
					a0_wr[345]     <= 0;                           
					a0_wr[346]     <= 0;                           
					a0_wr[347]     <= 0;                           
					a0_wr[348]     <= 0;                           
					a0_wr[349]     <= 0;                           
					a0_wr[350]     <= 0;                           
					a0_wr[351]     <= 0;                           
					a0_wr[352]     <= 0;                           
					a0_wr[353]     <= 0;                           
					a0_wr[354]     <= 0;                           
					a0_wr[355]     <= 0;                           
					a0_wr[356]     <= 0;                           
					a0_wr[357]     <= 0;                           
					a0_wr[358]     <= 0;                           
					a0_wr[359]     <= 0;                           
					a0_wr[360]     <= 0;                           
					a0_wr[361]     <= 0;                           
					a0_wr[362]     <= 0;                           
					a0_wr[363]     <= 0;                           
					a0_wr[364]     <= 0;                           
					a0_wr[365]     <= 0;                           
					a0_wr[366]     <= 0;                           
					a0_wr[367]     <= 0;                           
					a0_wr[368]     <= 0;                           
					a0_wr[369]     <= 0;                           
					a0_wr[370]     <= 0;                           
					a0_wr[371]     <= 0;                           
					a0_wr[372]     <= 0;                           
					a0_wr[373]     <= 0;                           
					a0_wr[374]     <= 0;                           
					a0_wr[375]     <= 0;                           
					a0_wr[376]     <= 0;                           
					a0_wr[377]     <= 0;                           
					a0_wr[378]     <= 0;                           
					a0_wr[379]     <= 0;                           
					a0_wr[380]     <= 0;                           
					a0_wr[381]     <= 0;                           
					a0_wr[382]     <= 0;                           
					a0_wr[383]     <= 0;                           
					a0_wr[384]     <= 0;                           
					a0_wr[385]     <= 0;                           
					a0_wr[386]     <= 0;                           
					a0_wr[387]     <= 0;                           
					a0_wr[388]     <= 0;                           
					a0_wr[389]     <= 0;                           
					a0_wr[390]     <= 0;                           
					a0_wr[391]     <= 0;                           
					a0_wr[392]     <= 0;                           
					a0_wr[393]     <= 0;                           
					a0_wr[394]     <= 0;                           
					a0_wr[395]     <= 0;                           
					a0_wr[396]     <= 0;                           
					a0_wr[397]     <= 0;                           
					a0_wr[398]     <= 0;                           
					a0_wr[399]     <= 0;                           
					a0_wr[400]     <= 0;                           
					a0_wr[401]     <= 0;                           
					a0_wr[402]     <= 0;                           
					a0_wr[403]     <= 0;                           
					a0_wr[404]     <= 0;                           
					a0_wr[405]     <= 0;                           
					a0_wr[406]     <= 0;                           
					a0_wr[407]     <= 0;                           
					a0_wr[408]     <= 0;                           
					a0_wr[409]     <= 0;                           
					a0_wr[410]     <= 0;                           
					a0_wr[411]     <= 0;                           
					a0_wr[412]     <= 0;                           
					a0_wr[413]     <= 0;                           
					a0_wr[414]     <= 0;                           
					a0_wr[415]     <= 0;                           
					a0_wr[416]     <= 0;                           
					a0_wr[417]     <= 0;                           
					a0_wr[418]     <= 0;                           
					a0_wr[419]     <= 0;                           
					a0_wr[420]     <= 0;                           
					a0_wr[421]     <= 0;                           
					a0_wr[422]     <= 0;                           
					a0_wr[423]     <= 0;                           
					a0_wr[424]     <= 0;                           
					a0_wr[425]     <= 0;                           
					a0_wr[426]     <= 0;                           
					a0_wr[427]     <= 0;                           
					a0_wr[428]     <= 0;                           
					a0_wr[429]     <= 0;                           
					a0_wr[430]     <= 0;                           
					a0_wr[431]     <= 0;                           
					a0_wr[432]     <= 0;                           
					a0_wr[433]     <= 0;                           
					a0_wr[434]     <= 0;                           
					a0_wr[435]     <= 0;                           
					a0_wr[436]     <= 0;                           
					a0_wr[437]     <= 0;                           
					a0_wr[438]     <= 0;                           
					a0_wr[439]     <= 0;                           
					a0_wr[440]     <= 0;                           
					a0_wr[441]     <= 0;                           
					a0_wr[442]     <= 0;                           
					a0_wr[443]     <= 0;                           
					a0_wr[444]     <= 0;                           
					a0_wr[445]     <= 0;                           
					a0_wr[446]     <= 0;                           
					a0_wr[447]     <= 0;                           
					a0_wr[448]     <= 0;                           
					a0_wr[449]     <= 0;                           
					a0_wr[450]     <= 0;                           
					a0_wr[451]     <= 0;                           
					a0_wr[452]     <= 0;                           
					a0_wr[453]     <= 0;                           
					a0_wr[454]     <= 0;                           
					a0_wr[455]     <= 0;                           
					a0_wr[456]     <= 0;                           
					a0_wr[457]     <= 0;                           
					a0_wr[458]     <= 0;                           
					a0_wr[459]     <= 0;                           
					a0_wr[460]     <= 0;                           
					a0_wr[461]     <= 0;                           
					a0_wr[462]     <= 0;                           
					a0_wr[463]     <= 0;                           
					a0_wr[464]     <= 0;                           
					a0_wr[465]     <= 0;                           
					a0_wr[466]     <= 0;                           
					a0_wr[467]     <= 0;                           
					a0_wr[468]     <= 0;                           
					a0_wr[469]     <= 0;                           
					a0_wr[470]     <= 0;                           
					a0_wr[471]     <= 0;                           
					a0_wr[472]     <= 0;                           
					a0_wr[473]     <= 0;                           
					a0_wr[474]     <= 0;                           
					a0_wr[475]     <= 0;                           
					a0_wr[476]     <= 0;                           
					a0_wr[477]     <= 0;                           
					a0_wr[478]     <= 0;                           
					a0_wr[479]     <= 0;                           
					a0_wr[480]     <= 0;                           
					a0_wr[481]     <= 0;                           
					a0_wr[482]     <= 0;                           
					a0_wr[483]     <= 0;                           
					a0_wr[484]     <= 0;                           
					a0_wr[485]     <= 0;                           
					a0_wr[486]     <= 0;                           
					a0_wr[487]     <= 0;                           
					a0_wr[488]     <= 0;                           
					a0_wr[489]     <= 0;                           
					a0_wr[490]     <= 0;                           
					a0_wr[491]     <= 0;                           
					a0_wr[492]     <= 0;                           
					a0_wr[493]     <= 0;                           
					a0_wr[494]     <= 0;                           
					a0_wr[495]     <= 0;                           
					a0_wr[496]     <= 0;                           
					a0_wr[497]     <= 0;                           
					a0_wr[498]     <= 0;                           
					a0_wr[499]     <= 0;                           
					a0_wr[500]     <= 0;                           
					a0_wr[501]     <= 0;                           
					a0_wr[502]     <= 0;                           
					a0_wr[503]     <= 0;                           
					a0_wr[504]     <= 0;                           
					a0_wr[505]     <= 0;                           
					a0_wr[506]     <= 0;                           
					a0_wr[507]     <= 0;                           
					a0_wr[508]     <= 0;                           
					a0_wr[509]     <= 0;                           
					a0_wr[510]     <= 0;                           
					a0_wr[511]     <= 0;                           
					a0_wr[512]     <= 0;                           
					a0_wr[513]     <= 0;                           
					a0_wr[514]     <= 0;                           
					a0_wr[515]     <= 0;                           
					a0_wr[516]     <= 0;                           
					a0_wr[517]     <= 0;                           
					a0_wr[518]     <= 0;                           
					a0_wr[519]     <= 0;                           
					a0_wr[520]     <= 0;                           
					a0_wr[521]     <= 0;                           
					a0_wr[522]     <= 0;                           
					a0_wr[523]     <= 0;                           
					a0_wr[524]     <= 0;                           
					a0_wr[525]     <= 0;                           
					a0_wr[526]     <= 0;                           
					a0_wr[527]     <= 0;                           
					a0_wr[528]     <= 0;                           
					a0_wr[529]     <= 0;                           
					a0_wr[530]     <= 0;                           
					a0_wr[531]     <= 0;                           
					a0_wr[532]     <= 0;                           
					a0_wr[533]     <= 0;                           
					a0_wr[534]     <= 0;                           
					a0_wr[535]     <= 0;                           
					a0_wr[536]     <= 0;                           
					a0_wr[537]     <= 0;                           
					a0_wr[538]     <= 0;                           
					a0_wr[539]     <= 0;                           
					a0_wr[540]     <= 0;                           
					a0_wr[541]     <= 0;                           
					a0_wr[542]     <= 0;                           
					a0_wr[543]     <= 0;                           
					a0_wr[544]     <= 0;                           
					a0_wr[545]     <= 0;                           
					a0_wr[546]     <= 0;                           
					a0_wr[547]     <= 0;                           
					a0_wr[548]     <= 0;                           
					a0_wr[549]     <= 0;                           
					a0_wr[550]     <= 0;                           
					a0_wr[551]     <= 0;                           
					a0_wr[552]     <= 0;                           
					a0_wr[553]     <= 0;                           
					a0_wr[554]     <= 0;                           
					a0_wr[555]     <= 0;                           
					a0_wr[556]     <= 0;                           
					a0_wr[557]     <= 0;                           
					a0_wr[558]     <= 0;                           
					a0_wr[559]     <= 0;                           
					a0_wr[560]     <= 0;                           
					a0_wr[561]     <= 0;                           
					a0_wr[562]     <= 0;                           
					a0_wr[563]     <= 0;                           
					a0_wr[564]     <= 0;                           
					a0_wr[565]     <= 0;                           
					a0_wr[566]     <= 0;                           
					a0_wr[567]     <= 0;                           
					a0_wr[568]     <= 0;                           
					a0_wr[569]     <= 0;                           
					a0_wr[570]     <= 0;                           
					a0_wr[571]     <= 0;                           
					a0_wr[572]     <= 0;                           
					a0_wr[573]     <= 0;                           
					a0_wr[574]     <= 0;                           
					a0_wr[575]     <= 0;                           
					a0_wr[576]     <= 0;                           
					a0_wr[577]     <= 0;                           
					a0_wr[578]     <= 0;                           
					a0_wr[579]     <= 0;                           
					a0_wr[580]     <= 0;                           
					a0_wr[581]     <= 0;                           
					a0_wr[582]     <= 0;                           
					a0_wr[583]     <= 0;                           
					a0_wr[584]     <= 0;                           
					a0_wr[585]     <= 0;                           
					a0_wr[586]     <= 0;                           
					a0_wr[587]     <= 0;                           
					a0_wr[588]     <= 0;                           
					a0_wr[589]     <= 0;                           
					a0_wr[590]     <= 0;                           
					a0_wr[591]     <= 0;                           
					a0_wr[592]     <= 0;                           
					a0_wr[593]     <= 0;                           
					a0_wr[594]     <= 0;                           
					a0_wr[595]     <= 0;                           
					a0_wr[596]     <= 0;                           
					a0_wr[597]     <= 0;                           
					a0_wr[598]     <= 0;                           
					a0_wr[599]     <= 0;                           
					a0_wr[600]     <= 0;                           
					a0_wr[601]     <= 0;                           
					a0_wr[602]     <= 0;                           
					a0_wr[603]     <= 0;                           
					a0_wr[604]     <= 0;                           
					a0_wr[605]     <= 0;                           
					a0_wr[606]     <= 0;                           
					a0_wr[607]     <= 0;                           
					a0_wr[608]     <= 0;                           
					a0_wr[609]     <= 0;                           
					a0_wr[610]     <= 0;                           
					a0_wr[611]     <= 0;                           
					a0_wr[612]     <= 0;                           
					a0_wr[613]     <= 0;                           
					a0_wr[614]     <= 0;                           
					a0_wr[615]     <= 0;                           
					a0_wr[616]     <= 0;                           
					a0_wr[617]     <= 0;                           
					a0_wr[618]     <= 0;                           
					a0_wr[619]     <= 0;                           
					a0_wr[620]     <= 0;                           
					a0_wr[621]     <= 0;                           
					a0_wr[622]     <= 0;                           
					a0_wr[623]     <= 0;                           
					a0_wr[624]     <= 0;                           
					a0_wr[625]     <= 0;                           
					a0_wr[626]     <= 0;                           
					a0_wr[627]     <= 0;                           
					a0_wr[628]     <= 0;                           
					a0_wr[629]     <= 0;                           
					a0_wr[630]     <= 0;                           
					a0_wr[631]     <= 0;                           
					a0_wr[632]     <= 0;                           
					a0_wr[633]     <= 0;                           
					a0_wr[634]     <= 0;                           
					a0_wr[635]     <= 0;                           
					a0_wr[636]     <= 0;                           
					a0_wr[637]     <= 0;                           
					a0_wr[638]     <= 0;                           
					a0_wr[639]     <= 0;                           
					a0_wr[640]     <= 0;                           
					a0_wr[641]     <= 0;                           
					a0_wr[642]     <= 0;                           
					a0_wr[643]     <= 0;                           
					a0_wr[644]     <= 0;                           
					a0_wr[645]     <= 0;                           
					a0_wr[646]     <= 0;                           
					a0_wr[647]     <= 0;                           
					a0_wr[648]     <= 0;                           
					a0_wr[649]     <= 0;                           
					a0_wr[650]     <= 0;                           
					a0_wr[651]     <= 0;                           
					a0_wr[652]     <= 0;                           
					a0_wr[653]     <= 0;                           
					a0_wr[654]     <= 0;                           
					a0_wr[655]     <= 0;                           
					a0_wr[656]     <= 0;                           
					a0_wr[657]     <= 0;                           
					a0_wr[658]     <= 0;                           
					a0_wr[659]     <= 0;                           
					a0_wr[660]     <= 0;                           
					a0_wr[661]     <= 0;                           
					a0_wr[662]     <= 0;                           
					a0_wr[663]     <= 0;                           
					a0_wr[664]     <= 0;                           
					a0_wr[665]     <= 0;                           
					a0_wr[666]     <= 0;                           
					a0_wr[667]     <= 0;                           
					a0_wr[668]     <= 0;                           
					a0_wr[669]     <= 0;                           
					a0_wr[670]     <= 0;                           
					a0_wr[671]     <= 0;                           
					a0_wr[672]     <= 0;                           
					a0_wr[673]     <= 0;                           
					a0_wr[674]     <= 0;                           
					a0_wr[675]     <= 0;                           
					a0_wr[676]     <= 0;                           
					a0_wr[677]     <= 0;                           
					a0_wr[678]     <= 0;                           
					a0_wr[679]     <= 0;                           
					a0_wr[680]     <= 0;                           
					a0_wr[681]     <= 0;                           
					a0_wr[682]     <= 0;                           
					a0_wr[683]     <= 0;                           
					a0_wr[684]     <= 0;                           
					a0_wr[685]     <= 0;                           
					a0_wr[686]     <= 0;                           
					a0_wr[687]     <= 0;                           
					a0_wr[688]     <= 0;                           
					a0_wr[689]     <= 0;                           
					a0_wr[690]     <= 0;                           
					a0_wr[691]     <= 0;                           
					a0_wr[692]     <= 0;                           
					a0_wr[693]     <= 0;                           
					a0_wr[694]     <= 0;                           
					a0_wr[695]     <= 0;                           
					a0_wr[696]     <= 0;                           
					a0_wr[697]     <= 0;                           
					a0_wr[698]     <= 0;                           
					a0_wr[699]     <= 0;                           
					a0_wr[700]     <= 0;                           
					a0_wr[701]     <= 0;                           
					a0_wr[702]     <= 0;                           
					a0_wr[703]     <= 0;                           
					a0_wr[704]     <= 0;                           
					a0_wr[705]     <= 0;                           
					a0_wr[706]     <= 0;                           
					a0_wr[707]     <= 0;                           
					a0_wr[708]     <= 0;                           
					a0_wr[709]     <= 0;                           
					a0_wr[710]     <= 0;                           
					a0_wr[711]     <= 0;                           
					a0_wr[712]     <= 0;                           
					a0_wr[713]     <= 0;                           
					a0_wr[714]     <= 0;                           
					a0_wr[715]     <= 0;                           
					a0_wr[716]     <= 0;                           
					a0_wr[717]     <= 0;                           
					a0_wr[718]     <= 0;                           
					a0_wr[719]     <= 0;                           
					a0_wr[720]     <= 0;                           
					a0_wr[721]     <= 0;                           
					a0_wr[722]     <= 0;                           
					a0_wr[723]     <= 0;                           
					a0_wr[724]     <= 0;                           
					a0_wr[725]     <= 0;                           
					a0_wr[726]     <= 0;                           
					a0_wr[727]     <= 0;                           
					a0_wr[728]     <= 0;                           
					a0_wr[729]     <= 0;                           
					a0_wr[730]     <= 0;                           
					a0_wr[731]     <= 0;                           
					a0_wr[732]     <= 0;                           
					a0_wr[733]     <= 0;                           
					a0_wr[734]     <= 0;                           
					a0_wr[735]     <= 0;                           
					a0_wr[736]     <= 0;                           
					a0_wr[737]     <= 0;                           
					a0_wr[738]     <= 0;                           
					a0_wr[739]     <= 0;                           
					a0_wr[740]     <= 0;                           
					a0_wr[741]     <= 0;                           
					a0_wr[742]     <= 0;                           
					a0_wr[743]     <= 0;                           
					a0_wr[744]     <= 0;                           
					a0_wr[745]     <= 0;                           
					a0_wr[746]     <= 0;                           
					a0_wr[747]     <= 0;                           
					a0_wr[748]     <= 0;                           
					a0_wr[749]     <= 0;                           
					a0_wr[750]     <= 0;                           
					a0_wr[751]     <= 0;                           
					a0_wr[752]     <= 0;                           
					a0_wr[753]     <= 0;                           
					a0_wr[754]     <= 0;                           
					a0_wr[755]     <= 0;                           
					a0_wr[756]     <= 0;                           
					a0_wr[757]     <= 0;                           
					a0_wr[758]     <= 0;                           
					a0_wr[759]     <= 0;                           
					a0_wr[760]     <= 0;                           
					a0_wr[761]     <= 0;                           
					a0_wr[762]     <= 0;                           
					a0_wr[763]     <= 0;                           
					a0_wr[764]     <= 0;                           
					a0_wr[765]     <= 0;                           
					a0_wr[766]     <= 0;                           
					a0_wr[767]     <= 0;                           
					a0_wr[768]     <= 0;                           
					a0_wr[769]     <= 0;                           
					a0_wr[770]     <= 0;                           
					a0_wr[771]     <= 0;                           
					a0_wr[772]     <= 0;                           
					a0_wr[773]     <= 0;                           
					a0_wr[774]     <= 0;                           
					a0_wr[775]     <= 0;                           
					a0_wr[776]     <= 0;                           
					a0_wr[777]     <= 0;                           
					a0_wr[778]     <= 0;                           
					a0_wr[779]     <= 0;                           
					a0_wr[780]     <= 0;                           
					a0_wr[781]     <= 0;                           
					a0_wr[782]     <= 0;                           
					a0_wr[783]     <= 0;                           
					a0_wr[784]     <= 0;                           
					a0_wr[785]     <= 0;                           
					a0_wr[786]     <= 0;                           
					a0_wr[787]     <= 0;                           
					a0_wr[788]     <= 0;                           
					a0_wr[789]     <= 0;                           
					a0_wr[790]     <= 0;                           
					a0_wr[791]     <= 0;                           
					a0_wr[792]     <= 0;                           
					a0_wr[793]     <= 0;                           
					a0_wr[794]     <= 0;                           
					a0_wr[795]     <= 0;                           
					a0_wr[796]     <= 0;                           
					a0_wr[797]     <= 0;                           
					a0_wr[798]     <= 0;                           
					a0_wr[799]     <= 0;                           
					a0_wr[800]     <= 0;                           
					a0_wr[801]     <= 0;                           
					a0_wr[802]     <= 0;                           
					a0_wr[803]     <= 0;                           
					a0_wr[804]     <= 0;                           
					a0_wr[805]     <= 0;                           
					a0_wr[806]     <= 0;                           
					a0_wr[807]     <= 0;                           
					a0_wr[808]     <= 0;                           
					a0_wr[809]     <= 0;                           
					a0_wr[810]     <= 0;                           
					a0_wr[811]     <= 0;                           
					a0_wr[812]     <= 0;                           
					a0_wr[813]     <= 0;                           
					a0_wr[814]     <= 0;                           
					a0_wr[815]     <= 0;                           
					a0_wr[816]     <= 0;                           
					a0_wr[817]     <= 0;                           
					a0_wr[818]     <= 0;                           
					a0_wr[819]     <= 0;                           
					a0_wr[820]     <= 0;                           
					a0_wr[821]     <= 0;                           
					a0_wr[822]     <= 0;                           
					a0_wr[823]     <= 0;                           
					a0_wr[824]     <= 0;                           
					a0_wr[825]     <= 0;                           
					a0_wr[826]     <= 0;                           
					a0_wr[827]     <= 0;                           
					a0_wr[828]     <= 0;                           
					a0_wr[829]     <= 0;                           
					a0_wr[830]     <= 0;                           
					a0_wr[831]     <= 0;                           
					a0_wr[832]     <= 0;                           
					a0_wr[833]     <= 0;                           
					a0_wr[834]     <= 0;                           
					a0_wr[835]     <= 0;                           
					a0_wr[836]     <= 0;                           
					a0_wr[837]     <= 0;                           
					a0_wr[838]     <= 0;                           
					a0_wr[839]     <= 0;                           
					a0_wr[840]     <= 0;                           
					a0_wr[841]     <= 0;                           
					a0_wr[842]     <= 0;                           
					a0_wr[843]     <= 0;                           
					a0_wr[844]     <= 0;                           
					a0_wr[845]     <= 0;                           
					a0_wr[846]     <= 0;                           
					a0_wr[847]     <= 0;                           
					a0_wr[848]     <= 0;                           
					a0_wr[849]     <= 0;                           
					a0_wr[850]     <= 0;                           
					a0_wr[851]     <= 0;                           
					a0_wr[852]     <= 0;                           
					a0_wr[853]     <= 0;                           
					a0_wr[854]     <= 0;                           
					a0_wr[855]     <= 0;                           
					a0_wr[856]     <= 0;                           
					a0_wr[857]     <= 0;                           
					a0_wr[858]     <= 0;                           
					a0_wr[859]     <= 0;                           
					a0_wr[860]     <= 0;                           
					a0_wr[861]     <= 0;                           
					a0_wr[862]     <= 0;                           
					a0_wr[863]     <= 0;                           
					a0_wr[864]     <= 0;                           
					a0_wr[865]     <= 0;                           
					a0_wr[866]     <= 0;                           
					a0_wr[867]     <= 0;                           
					a0_wr[868]     <= 0;                           
					a0_wr[869]     <= 0;                           
					a0_wr[870]     <= 0;                           
					a0_wr[871]     <= 0;                           
					a0_wr[872]     <= 0;                           
					a0_wr[873]     <= 0;                           
					a0_wr[874]     <= 0;                           
					a0_wr[875]     <= 0;                           
					a0_wr[876]     <= 0;                           
					a0_wr[877]     <= 0;                           
					a0_wr[878]     <= 0;                           
					a0_wr[879]     <= 0;                           
					a0_wr[880]     <= 0;                           
					a0_wr[881]     <= 0;                           
					a0_wr[882]     <= 0;                           
					a0_wr[883]     <= 0;                           
					a0_wr[884]     <= 0;                           
					a0_wr[885]     <= 0;                           
					a0_wr[886]     <= 0;                           
					a0_wr[887]     <= 0;                           
					a0_wr[888]     <= 0;                           
					a0_wr[889]     <= 0;                           
					a0_wr[890]     <= 0;                           
					a0_wr[891]     <= 0;                           
					a0_wr[892]     <= 0;                           
					a0_wr[893]     <= 0;                           
					a0_wr[894]     <= 0;                           
					a0_wr[895]     <= 0;                           
					a0_wr[896]     <= 0;                           
					a0_wr[897]     <= 0;                           
					a0_wr[898]     <= 0;                           
					a0_wr[899]     <= 0;                           
					a0_wr[900]     <= 0;                           
					a0_wr[901]     <= 0;                           
					a0_wr[902]     <= 0;                           
					a0_wr[903]     <= 0;                           
					a0_wr[904]     <= 0;                           
					a0_wr[905]     <= 0;                           
					a0_wr[906]     <= 0;                           
					a0_wr[907]     <= 0;                           
					a0_wr[908]     <= 0;                           
					a0_wr[909]     <= 0;                           
					a0_wr[910]     <= 0;                           
					a0_wr[911]     <= 0;                           
					a0_wr[912]     <= 0;                           
					a0_wr[913]     <= 0;                           
					a0_wr[914]     <= 0;                           
					a0_wr[915]     <= 0;                           
					a0_wr[916]     <= 0;                           
					a0_wr[917]     <= 0;                           
					a0_wr[918]     <= 0;                           
					a0_wr[919]     <= 0;                           
					a0_wr[920]     <= 0;                           
					a0_wr[921]     <= 0;                           
					a0_wr[922]     <= 0;                           
					a0_wr[923]     <= 0;                           
					a0_wr[924]     <= 0;                           
					a0_wr[925]     <= 0;                           
					a0_wr[926]     <= 0;                           
					a0_wr[927]     <= 0;                           
					a0_wr[928]     <= 0;                           
					a0_wr[929]     <= 0;                           
					a0_wr[930]     <= 0;                           
					a0_wr[931]     <= 0;                           
					a0_wr[932]     <= 0;                           
					a0_wr[933]     <= 0;                           
					a0_wr[934]     <= 0;                           
					a0_wr[935]     <= 0;                           
					a0_wr[936]     <= 0;                           
					a0_wr[937]     <= 0;                           
					a0_wr[938]     <= 0;                           
					a0_wr[939]     <= 0;                           
					a0_wr[940]     <= 0;                           
					a0_wr[941]     <= 0;                           
					a0_wr[942]     <= 0;                           
					a0_wr[943]     <= 0;                           
					a0_wr[944]     <= 0;                           
					a0_wr[945]     <= 0;                           
					a0_wr[946]     <= 0;                           
					a0_wr[947]     <= 0;                           
					a0_wr[948]     <= 0;                           
					a0_wr[949]     <= 0;                           
					a0_wr[950]     <= 0;                           
					a0_wr[951]     <= 0;                           
					a0_wr[952]     <= 0;                           
					a0_wr[953]     <= 0;                           
					a0_wr[954]     <= 0;                           
					a0_wr[955]     <= 0;                           
					a0_wr[956]     <= 0;                           
					a0_wr[957]     <= 0;                           
					a0_wr[958]     <= 0;                           
					a0_wr[959]     <= 0;                           
					a0_wr[960]     <= 0;                           
					a0_wr[961]     <= 0;                           
					a0_wr[962]     <= 0;                           
					a0_wr[963]     <= 0;                           
					a0_wr[964]     <= 0;                           
					a0_wr[965]     <= 0;                           
					a0_wr[966]     <= 0;                           
					a0_wr[967]     <= 0;                           
					a0_wr[968]     <= 0;                           
					a0_wr[969]     <= 0;                           
					a0_wr[970]     <= 0;                           
					a0_wr[971]     <= 0;                           
					a0_wr[972]     <= 0;                           
					a0_wr[973]     <= 0;                           
					a0_wr[974]     <= 0;                           
					a0_wr[975]     <= 0;                           
					a0_wr[976]     <= 0;                           
					a0_wr[977]     <= 0;                           
					a0_wr[978]     <= 0;                           
					a0_wr[979]     <= 0;                           
					a0_wr[980]     <= 0;                           
					a0_wr[981]     <= 0;                           
					a0_wr[982]     <= 0;                           
					a0_wr[983]     <= 0;                           
					a0_wr[984]     <= 0;                           
					a0_wr[985]     <= 0;                           
					a0_wr[986]     <= 0;                           
					a0_wr[987]     <= 0;                           
					a0_wr[988]     <= 0;                           
					a0_wr[989]     <= 0;                           
					a0_wr[990]     <= 0;                           
					a0_wr[991]     <= 0;                           
					a0_wr[992]     <= 0;                           
					a0_wr[993]     <= 0;                           
					a0_wr[994]     <= 0;                           
					a0_wr[995]     <= 0;                           
					a0_wr[996]     <= 0;                           
					a0_wr[997]     <= 0;                           
					a0_wr[998]     <= 0;                           
					a0_wr[999]     <= 0;                           
					a0_wr[1000]    <= 0;                           
					a0_wr[1001]    <= 0;                           
					a0_wr[1002]    <= 0;                           
					a0_wr[1003]    <= 0;                           
					a0_wr[1004]    <= 0;                           
					a0_wr[1005]    <= 0;                           
					a0_wr[1006]    <= 0;                           
					a0_wr[1007]    <= 0;                           
					a0_wr[1008]    <= 0;                           
					a0_wr[1009]    <= 0;                           
					a0_wr[1010]    <= 0;                           
					a0_wr[1011]    <= 0;                           
					a0_wr[1012]    <= 0;                           
					a0_wr[1013]    <= 0;                           
					a0_wr[1014]    <= 0;                           
					a0_wr[1015]    <= 0;                           
					a0_wr[1016]    <= 0;                           
					a0_wr[1017]    <= 0;                           
					a0_wr[1018]    <= 0;                           
					a0_wr[1019]    <= 0;                           
					a0_wr[1020]    <= 0;                           
					a0_wr[1021]    <= 0;                           
					a0_wr[1022]    <= 0;                           
					a0_wr[1023]    <= 0;                           
				end
				else begin
					if (!stall) begin
						a0_wr[0]      <= x0_in;                       
						a0_wr[1]      <= x1_in;                       
						a0_wr[2]      <= x2_in;                       
						a0_wr[3]      <= x3_in;                       
						a0_wr[4]      <= x4_in;                       
						a0_wr[5]      <= x5_in;                       
						a0_wr[6]      <= x6_in;                       
						a0_wr[7]      <= x7_in;                       
						a0_wr[8]      <= x8_in;                       
						a0_wr[9]      <= x9_in;                       
						a0_wr[10]     <= x10_in;                      
						a0_wr[11]     <= x11_in;                      
						a0_wr[12]     <= x12_in;                      
						a0_wr[13]     <= x13_in;                      
						a0_wr[14]     <= x14_in;                      
						a0_wr[15]     <= x15_in;                      
						a0_wr[16]     <= x16_in;                      
						a0_wr[17]     <= x17_in;                      
						a0_wr[18]     <= x18_in;                      
						a0_wr[19]     <= x19_in;                      
						a0_wr[20]     <= x20_in;                      
						a0_wr[21]     <= x21_in;                      
						a0_wr[22]     <= x22_in;                      
						a0_wr[23]     <= x23_in;                      
						a0_wr[24]     <= x24_in;                      
						a0_wr[25]     <= x25_in;                      
						a0_wr[26]     <= x26_in;                      
						a0_wr[27]     <= x27_in;                      
						a0_wr[28]     <= x28_in;                      
						a0_wr[29]     <= x29_in;                      
						a0_wr[30]     <= x30_in;                      
						a0_wr[31]     <= x31_in;                      
						a0_wr[32]     <= x32_in;                      
						a0_wr[33]     <= x33_in;                      
						a0_wr[34]     <= x34_in;                      
						a0_wr[35]     <= x35_in;                      
						a0_wr[36]     <= x36_in;                      
						a0_wr[37]     <= x37_in;                      
						a0_wr[38]     <= x38_in;                      
						a0_wr[39]     <= x39_in;                      
						a0_wr[40]     <= x40_in;                      
						a0_wr[41]     <= x41_in;                      
						a0_wr[42]     <= x42_in;                      
						a0_wr[43]     <= x43_in;                      
						a0_wr[44]     <= x44_in;                      
						a0_wr[45]     <= x45_in;                      
						a0_wr[46]     <= x46_in;                      
						a0_wr[47]     <= x47_in;                      
						a0_wr[48]     <= x48_in;                      
						a0_wr[49]     <= x49_in;                      
						a0_wr[50]     <= x50_in;                      
						a0_wr[51]     <= x51_in;                      
						a0_wr[52]     <= x52_in;                      
						a0_wr[53]     <= x53_in;                      
						a0_wr[54]     <= x54_in;                      
						a0_wr[55]     <= x55_in;                      
						a0_wr[56]     <= x56_in;                      
						a0_wr[57]     <= x57_in;                      
						a0_wr[58]     <= x58_in;                      
						a0_wr[59]     <= x59_in;                      
						a0_wr[60]     <= x60_in;                      
						a0_wr[61]     <= x61_in;                      
						a0_wr[62]     <= x62_in;                      
						a0_wr[63]     <= x63_in;                      
						a0_wr[64]     <= x64_in;                      
						a0_wr[65]     <= x65_in;                      
						a0_wr[66]     <= x66_in;                      
						a0_wr[67]     <= x67_in;                      
						a0_wr[68]     <= x68_in;                      
						a0_wr[69]     <= x69_in;                      
						a0_wr[70]     <= x70_in;                      
						a0_wr[71]     <= x71_in;                      
						a0_wr[72]     <= x72_in;                      
						a0_wr[73]     <= x73_in;                      
						a0_wr[74]     <= x74_in;                      
						a0_wr[75]     <= x75_in;                      
						a0_wr[76]     <= x76_in;                      
						a0_wr[77]     <= x77_in;                      
						a0_wr[78]     <= x78_in;                      
						a0_wr[79]     <= x79_in;                      
						a0_wr[80]     <= x80_in;                      
						a0_wr[81]     <= x81_in;                      
						a0_wr[82]     <= x82_in;                      
						a0_wr[83]     <= x83_in;                      
						a0_wr[84]     <= x84_in;                      
						a0_wr[85]     <= x85_in;                      
						a0_wr[86]     <= x86_in;                      
						a0_wr[87]     <= x87_in;                      
						a0_wr[88]     <= x88_in;                      
						a0_wr[89]     <= x89_in;                      
						a0_wr[90]     <= x90_in;                      
						a0_wr[91]     <= x91_in;                      
						a0_wr[92]     <= x92_in;                      
						a0_wr[93]     <= x93_in;                      
						a0_wr[94]     <= x94_in;                      
						a0_wr[95]     <= x95_in;                      
						a0_wr[96]     <= x96_in;                      
						a0_wr[97]     <= x97_in;                      
						a0_wr[98]     <= x98_in;                      
						a0_wr[99]     <= x99_in;                      
						a0_wr[100]    <= x100_in;                     
						a0_wr[101]    <= x101_in;                     
						a0_wr[102]    <= x102_in;                     
						a0_wr[103]    <= x103_in;                     
						a0_wr[104]    <= x104_in;                     
						a0_wr[105]    <= x105_in;                     
						a0_wr[106]    <= x106_in;                     
						a0_wr[107]    <= x107_in;                     
						a0_wr[108]    <= x108_in;                     
						a0_wr[109]    <= x109_in;                     
						a0_wr[110]    <= x110_in;                     
						a0_wr[111]    <= x111_in;                     
						a0_wr[112]    <= x112_in;                     
						a0_wr[113]    <= x113_in;                     
						a0_wr[114]    <= x114_in;                     
						a0_wr[115]    <= x115_in;                     
						a0_wr[116]    <= x116_in;                     
						a0_wr[117]    <= x117_in;                     
						a0_wr[118]    <= x118_in;                     
						a0_wr[119]    <= x119_in;                     
						a0_wr[120]    <= x120_in;                     
						a0_wr[121]    <= x121_in;                     
						a0_wr[122]    <= x122_in;                     
						a0_wr[123]    <= x123_in;                     
						a0_wr[124]    <= x124_in;                     
						a0_wr[125]    <= x125_in;                     
						a0_wr[126]    <= x126_in;                     
						a0_wr[127]    <= x127_in;                     
						a0_wr[128]    <= x128_in;                     
						a0_wr[129]    <= x129_in;                     
						a0_wr[130]    <= x130_in;                     
						a0_wr[131]    <= x131_in;                     
						a0_wr[132]    <= x132_in;                     
						a0_wr[133]    <= x133_in;                     
						a0_wr[134]    <= x134_in;                     
						a0_wr[135]    <= x135_in;                     
						a0_wr[136]    <= x136_in;                     
						a0_wr[137]    <= x137_in;                     
						a0_wr[138]    <= x138_in;                     
						a0_wr[139]    <= x139_in;                     
						a0_wr[140]    <= x140_in;                     
						a0_wr[141]    <= x141_in;                     
						a0_wr[142]    <= x142_in;                     
						a0_wr[143]    <= x143_in;                     
						a0_wr[144]    <= x144_in;                     
						a0_wr[145]    <= x145_in;                     
						a0_wr[146]    <= x146_in;                     
						a0_wr[147]    <= x147_in;                     
						a0_wr[148]    <= x148_in;                     
						a0_wr[149]    <= x149_in;                     
						a0_wr[150]    <= x150_in;                     
						a0_wr[151]    <= x151_in;                     
						a0_wr[152]    <= x152_in;                     
						a0_wr[153]    <= x153_in;                     
						a0_wr[154]    <= x154_in;                     
						a0_wr[155]    <= x155_in;                     
						a0_wr[156]    <= x156_in;                     
						a0_wr[157]    <= x157_in;                     
						a0_wr[158]    <= x158_in;                     
						a0_wr[159]    <= x159_in;                     
						a0_wr[160]    <= x160_in;                     
						a0_wr[161]    <= x161_in;                     
						a0_wr[162]    <= x162_in;                     
						a0_wr[163]    <= x163_in;                     
						a0_wr[164]    <= x164_in;                     
						a0_wr[165]    <= x165_in;                     
						a0_wr[166]    <= x166_in;                     
						a0_wr[167]    <= x167_in;                     
						a0_wr[168]    <= x168_in;                     
						a0_wr[169]    <= x169_in;                     
						a0_wr[170]    <= x170_in;                     
						a0_wr[171]    <= x171_in;                     
						a0_wr[172]    <= x172_in;                     
						a0_wr[173]    <= x173_in;                     
						a0_wr[174]    <= x174_in;                     
						a0_wr[175]    <= x175_in;                     
						a0_wr[176]    <= x176_in;                     
						a0_wr[177]    <= x177_in;                     
						a0_wr[178]    <= x178_in;                     
						a0_wr[179]    <= x179_in;                     
						a0_wr[180]    <= x180_in;                     
						a0_wr[181]    <= x181_in;                     
						a0_wr[182]    <= x182_in;                     
						a0_wr[183]    <= x183_in;                     
						a0_wr[184]    <= x184_in;                     
						a0_wr[185]    <= x185_in;                     
						a0_wr[186]    <= x186_in;                     
						a0_wr[187]    <= x187_in;                     
						a0_wr[188]    <= x188_in;                     
						a0_wr[189]    <= x189_in;                     
						a0_wr[190]    <= x190_in;                     
						a0_wr[191]    <= x191_in;                     
						a0_wr[192]    <= x192_in;                     
						a0_wr[193]    <= x193_in;                     
						a0_wr[194]    <= x194_in;                     
						a0_wr[195]    <= x195_in;                     
						a0_wr[196]    <= x196_in;                     
						a0_wr[197]    <= x197_in;                     
						a0_wr[198]    <= x198_in;                     
						a0_wr[199]    <= x199_in;                     
						a0_wr[200]    <= x200_in;                     
						a0_wr[201]    <= x201_in;                     
						a0_wr[202]    <= x202_in;                     
						a0_wr[203]    <= x203_in;                     
						a0_wr[204]    <= x204_in;                     
						a0_wr[205]    <= x205_in;                     
						a0_wr[206]    <= x206_in;                     
						a0_wr[207]    <= x207_in;                     
						a0_wr[208]    <= x208_in;                     
						a0_wr[209]    <= x209_in;                     
						a0_wr[210]    <= x210_in;                     
						a0_wr[211]    <= x211_in;                     
						a0_wr[212]    <= x212_in;                     
						a0_wr[213]    <= x213_in;                     
						a0_wr[214]    <= x214_in;                     
						a0_wr[215]    <= x215_in;                     
						a0_wr[216]    <= x216_in;                     
						a0_wr[217]    <= x217_in;                     
						a0_wr[218]    <= x218_in;                     
						a0_wr[219]    <= x219_in;                     
						a0_wr[220]    <= x220_in;                     
						a0_wr[221]    <= x221_in;                     
						a0_wr[222]    <= x222_in;                     
						a0_wr[223]    <= x223_in;                     
						a0_wr[224]    <= x224_in;                     
						a0_wr[225]    <= x225_in;                     
						a0_wr[226]    <= x226_in;                     
						a0_wr[227]    <= x227_in;                     
						a0_wr[228]    <= x228_in;                     
						a0_wr[229]    <= x229_in;                     
						a0_wr[230]    <= x230_in;                     
						a0_wr[231]    <= x231_in;                     
						a0_wr[232]    <= x232_in;                     
						a0_wr[233]    <= x233_in;                     
						a0_wr[234]    <= x234_in;                     
						a0_wr[235]    <= x235_in;                     
						a0_wr[236]    <= x236_in;                     
						a0_wr[237]    <= x237_in;                     
						a0_wr[238]    <= x238_in;                     
						a0_wr[239]    <= x239_in;                     
						a0_wr[240]    <= x240_in;                     
						a0_wr[241]    <= x241_in;                     
						a0_wr[242]    <= x242_in;                     
						a0_wr[243]    <= x243_in;                     
						a0_wr[244]    <= x244_in;                     
						a0_wr[245]    <= x245_in;                     
						a0_wr[246]    <= x246_in;                     
						a0_wr[247]    <= x247_in;                     
						a0_wr[248]    <= x248_in;                     
						a0_wr[249]    <= x249_in;                     
						a0_wr[250]    <= x250_in;                     
						a0_wr[251]    <= x251_in;                     
						a0_wr[252]    <= x252_in;                     
						a0_wr[253]    <= x253_in;                     
						a0_wr[254]    <= x254_in;                     
						a0_wr[255]    <= x255_in;                     
						a0_wr[256]    <= x256_in;                     
						a0_wr[257]    <= x257_in;                     
						a0_wr[258]    <= x258_in;                     
						a0_wr[259]    <= x259_in;                     
						a0_wr[260]    <= x260_in;                     
						a0_wr[261]    <= x261_in;                     
						a0_wr[262]    <= x262_in;                     
						a0_wr[263]    <= x263_in;                     
						a0_wr[264]    <= x264_in;                     
						a0_wr[265]    <= x265_in;                     
						a0_wr[266]    <= x266_in;                     
						a0_wr[267]    <= x267_in;                     
						a0_wr[268]    <= x268_in;                     
						a0_wr[269]    <= x269_in;                     
						a0_wr[270]    <= x270_in;                     
						a0_wr[271]    <= x271_in;                     
						a0_wr[272]    <= x272_in;                     
						a0_wr[273]    <= x273_in;                     
						a0_wr[274]    <= x274_in;                     
						a0_wr[275]    <= x275_in;                     
						a0_wr[276]    <= x276_in;                     
						a0_wr[277]    <= x277_in;                     
						a0_wr[278]    <= x278_in;                     
						a0_wr[279]    <= x279_in;                     
						a0_wr[280]    <= x280_in;                     
						a0_wr[281]    <= x281_in;                     
						a0_wr[282]    <= x282_in;                     
						a0_wr[283]    <= x283_in;                     
						a0_wr[284]    <= x284_in;                     
						a0_wr[285]    <= x285_in;                     
						a0_wr[286]    <= x286_in;                     
						a0_wr[287]    <= x287_in;                     
						a0_wr[288]    <= x288_in;                     
						a0_wr[289]    <= x289_in;                     
						a0_wr[290]    <= x290_in;                     
						a0_wr[291]    <= x291_in;                     
						a0_wr[292]    <= x292_in;                     
						a0_wr[293]    <= x293_in;                     
						a0_wr[294]    <= x294_in;                     
						a0_wr[295]    <= x295_in;                     
						a0_wr[296]    <= x296_in;                     
						a0_wr[297]    <= x297_in;                     
						a0_wr[298]    <= x298_in;                     
						a0_wr[299]    <= x299_in;                     
						a0_wr[300]    <= x300_in;                     
						a0_wr[301]    <= x301_in;                     
						a0_wr[302]    <= x302_in;                     
						a0_wr[303]    <= x303_in;                     
						a0_wr[304]    <= x304_in;                     
						a0_wr[305]    <= x305_in;                     
						a0_wr[306]    <= x306_in;                     
						a0_wr[307]    <= x307_in;                     
						a0_wr[308]    <= x308_in;                     
						a0_wr[309]    <= x309_in;                     
						a0_wr[310]    <= x310_in;                     
						a0_wr[311]    <= x311_in;                     
						a0_wr[312]    <= x312_in;                     
						a0_wr[313]    <= x313_in;                     
						a0_wr[314]    <= x314_in;                     
						a0_wr[315]    <= x315_in;                     
						a0_wr[316]    <= x316_in;                     
						a0_wr[317]    <= x317_in;                     
						a0_wr[318]    <= x318_in;                     
						a0_wr[319]    <= x319_in;                     
						a0_wr[320]    <= x320_in;                     
						a0_wr[321]    <= x321_in;                     
						a0_wr[322]    <= x322_in;                     
						a0_wr[323]    <= x323_in;                     
						a0_wr[324]    <= x324_in;                     
						a0_wr[325]    <= x325_in;                     
						a0_wr[326]    <= x326_in;                     
						a0_wr[327]    <= x327_in;                     
						a0_wr[328]    <= x328_in;                     
						a0_wr[329]    <= x329_in;                     
						a0_wr[330]    <= x330_in;                     
						a0_wr[331]    <= x331_in;                     
						a0_wr[332]    <= x332_in;                     
						a0_wr[333]    <= x333_in;                     
						a0_wr[334]    <= x334_in;                     
						a0_wr[335]    <= x335_in;                     
						a0_wr[336]    <= x336_in;                     
						a0_wr[337]    <= x337_in;                     
						a0_wr[338]    <= x338_in;                     
						a0_wr[339]    <= x339_in;                     
						a0_wr[340]    <= x340_in;                     
						a0_wr[341]    <= x341_in;                     
						a0_wr[342]    <= x342_in;                     
						a0_wr[343]    <= x343_in;                     
						a0_wr[344]    <= x344_in;                     
						a0_wr[345]    <= x345_in;                     
						a0_wr[346]    <= x346_in;                     
						a0_wr[347]    <= x347_in;                     
						a0_wr[348]    <= x348_in;                     
						a0_wr[349]    <= x349_in;                     
						a0_wr[350]    <= x350_in;                     
						a0_wr[351]    <= x351_in;                     
						a0_wr[352]    <= x352_in;                     
						a0_wr[353]    <= x353_in;                     
						a0_wr[354]    <= x354_in;                     
						a0_wr[355]    <= x355_in;                     
						a0_wr[356]    <= x356_in;                     
						a0_wr[357]    <= x357_in;                     
						a0_wr[358]    <= x358_in;                     
						a0_wr[359]    <= x359_in;                     
						a0_wr[360]    <= x360_in;                     
						a0_wr[361]    <= x361_in;                     
						a0_wr[362]    <= x362_in;                     
						a0_wr[363]    <= x363_in;                     
						a0_wr[364]    <= x364_in;                     
						a0_wr[365]    <= x365_in;                     
						a0_wr[366]    <= x366_in;                     
						a0_wr[367]    <= x367_in;                     
						a0_wr[368]    <= x368_in;                     
						a0_wr[369]    <= x369_in;                     
						a0_wr[370]    <= x370_in;                     
						a0_wr[371]    <= x371_in;                     
						a0_wr[372]    <= x372_in;                     
						a0_wr[373]    <= x373_in;                     
						a0_wr[374]    <= x374_in;                     
						a0_wr[375]    <= x375_in;                     
						a0_wr[376]    <= x376_in;                     
						a0_wr[377]    <= x377_in;                     
						a0_wr[378]    <= x378_in;                     
						a0_wr[379]    <= x379_in;                     
						a0_wr[380]    <= x380_in;                     
						a0_wr[381]    <= x381_in;                     
						a0_wr[382]    <= x382_in;                     
						a0_wr[383]    <= x383_in;                     
						a0_wr[384]    <= x384_in;                     
						a0_wr[385]    <= x385_in;                     
						a0_wr[386]    <= x386_in;                     
						a0_wr[387]    <= x387_in;                     
						a0_wr[388]    <= x388_in;                     
						a0_wr[389]    <= x389_in;                     
						a0_wr[390]    <= x390_in;                     
						a0_wr[391]    <= x391_in;                     
						a0_wr[392]    <= x392_in;                     
						a0_wr[393]    <= x393_in;                     
						a0_wr[394]    <= x394_in;                     
						a0_wr[395]    <= x395_in;                     
						a0_wr[396]    <= x396_in;                     
						a0_wr[397]    <= x397_in;                     
						a0_wr[398]    <= x398_in;                     
						a0_wr[399]    <= x399_in;                     
						a0_wr[400]    <= x400_in;                     
						a0_wr[401]    <= x401_in;                     
						a0_wr[402]    <= x402_in;                     
						a0_wr[403]    <= x403_in;                     
						a0_wr[404]    <= x404_in;                     
						a0_wr[405]    <= x405_in;                     
						a0_wr[406]    <= x406_in;                     
						a0_wr[407]    <= x407_in;                     
						a0_wr[408]    <= x408_in;                     
						a0_wr[409]    <= x409_in;                     
						a0_wr[410]    <= x410_in;                     
						a0_wr[411]    <= x411_in;                     
						a0_wr[412]    <= x412_in;                     
						a0_wr[413]    <= x413_in;                     
						a0_wr[414]    <= x414_in;                     
						a0_wr[415]    <= x415_in;                     
						a0_wr[416]    <= x416_in;                     
						a0_wr[417]    <= x417_in;                     
						a0_wr[418]    <= x418_in;                     
						a0_wr[419]    <= x419_in;                     
						a0_wr[420]    <= x420_in;                     
						a0_wr[421]    <= x421_in;                     
						a0_wr[422]    <= x422_in;                     
						a0_wr[423]    <= x423_in;                     
						a0_wr[424]    <= x424_in;                     
						a0_wr[425]    <= x425_in;                     
						a0_wr[426]    <= x426_in;                     
						a0_wr[427]    <= x427_in;                     
						a0_wr[428]    <= x428_in;                     
						a0_wr[429]    <= x429_in;                     
						a0_wr[430]    <= x430_in;                     
						a0_wr[431]    <= x431_in;                     
						a0_wr[432]    <= x432_in;                     
						a0_wr[433]    <= x433_in;                     
						a0_wr[434]    <= x434_in;                     
						a0_wr[435]    <= x435_in;                     
						a0_wr[436]    <= x436_in;                     
						a0_wr[437]    <= x437_in;                     
						a0_wr[438]    <= x438_in;                     
						a0_wr[439]    <= x439_in;                     
						a0_wr[440]    <= x440_in;                     
						a0_wr[441]    <= x441_in;                     
						a0_wr[442]    <= x442_in;                     
						a0_wr[443]    <= x443_in;                     
						a0_wr[444]    <= x444_in;                     
						a0_wr[445]    <= x445_in;                     
						a0_wr[446]    <= x446_in;                     
						a0_wr[447]    <= x447_in;                     
						a0_wr[448]    <= x448_in;                     
						a0_wr[449]    <= x449_in;                     
						a0_wr[450]    <= x450_in;                     
						a0_wr[451]    <= x451_in;                     
						a0_wr[452]    <= x452_in;                     
						a0_wr[453]    <= x453_in;                     
						a0_wr[454]    <= x454_in;                     
						a0_wr[455]    <= x455_in;                     
						a0_wr[456]    <= x456_in;                     
						a0_wr[457]    <= x457_in;                     
						a0_wr[458]    <= x458_in;                     
						a0_wr[459]    <= x459_in;                     
						a0_wr[460]    <= x460_in;                     
						a0_wr[461]    <= x461_in;                     
						a0_wr[462]    <= x462_in;                     
						a0_wr[463]    <= x463_in;                     
						a0_wr[464]    <= x464_in;                     
						a0_wr[465]    <= x465_in;                     
						a0_wr[466]    <= x466_in;                     
						a0_wr[467]    <= x467_in;                     
						a0_wr[468]    <= x468_in;                     
						a0_wr[469]    <= x469_in;                     
						a0_wr[470]    <= x470_in;                     
						a0_wr[471]    <= x471_in;                     
						a0_wr[472]    <= x472_in;                     
						a0_wr[473]    <= x473_in;                     
						a0_wr[474]    <= x474_in;                     
						a0_wr[475]    <= x475_in;                     
						a0_wr[476]    <= x476_in;                     
						a0_wr[477]    <= x477_in;                     
						a0_wr[478]    <= x478_in;                     
						a0_wr[479]    <= x479_in;                     
						a0_wr[480]    <= x480_in;                     
						a0_wr[481]    <= x481_in;                     
						a0_wr[482]    <= x482_in;                     
						a0_wr[483]    <= x483_in;                     
						a0_wr[484]    <= x484_in;                     
						a0_wr[485]    <= x485_in;                     
						a0_wr[486]    <= x486_in;                     
						a0_wr[487]    <= x487_in;                     
						a0_wr[488]    <= x488_in;                     
						a0_wr[489]    <= x489_in;                     
						a0_wr[490]    <= x490_in;                     
						a0_wr[491]    <= x491_in;                     
						a0_wr[492]    <= x492_in;                     
						a0_wr[493]    <= x493_in;                     
						a0_wr[494]    <= x494_in;                     
						a0_wr[495]    <= x495_in;                     
						a0_wr[496]    <= x496_in;                     
						a0_wr[497]    <= x497_in;                     
						a0_wr[498]    <= x498_in;                     
						a0_wr[499]    <= x499_in;                     
						a0_wr[500]    <= x500_in;                     
						a0_wr[501]    <= x501_in;                     
						a0_wr[502]    <= x502_in;                     
						a0_wr[503]    <= x503_in;                     
						a0_wr[504]    <= x504_in;                     
						a0_wr[505]    <= x505_in;                     
						a0_wr[506]    <= x506_in;                     
						a0_wr[507]    <= x507_in;                     
						a0_wr[508]    <= x508_in;                     
						a0_wr[509]    <= x509_in;                     
						a0_wr[510]    <= x510_in;                     
						a0_wr[511]    <= x511_in;                     
						a0_wr[512]    <= x512_in;                     
						a0_wr[513]    <= x513_in;                     
						a0_wr[514]    <= x514_in;                     
						a0_wr[515]    <= x515_in;                     
						a0_wr[516]    <= x516_in;                     
						a0_wr[517]    <= x517_in;                     
						a0_wr[518]    <= x518_in;                     
						a0_wr[519]    <= x519_in;                     
						a0_wr[520]    <= x520_in;                     
						a0_wr[521]    <= x521_in;                     
						a0_wr[522]    <= x522_in;                     
						a0_wr[523]    <= x523_in;                     
						a0_wr[524]    <= x524_in;                     
						a0_wr[525]    <= x525_in;                     
						a0_wr[526]    <= x526_in;                     
						a0_wr[527]    <= x527_in;                     
						a0_wr[528]    <= x528_in;                     
						a0_wr[529]    <= x529_in;                     
						a0_wr[530]    <= x530_in;                     
						a0_wr[531]    <= x531_in;                     
						a0_wr[532]    <= x532_in;                     
						a0_wr[533]    <= x533_in;                     
						a0_wr[534]    <= x534_in;                     
						a0_wr[535]    <= x535_in;                     
						a0_wr[536]    <= x536_in;                     
						a0_wr[537]    <= x537_in;                     
						a0_wr[538]    <= x538_in;                     
						a0_wr[539]    <= x539_in;                     
						a0_wr[540]    <= x540_in;                     
						a0_wr[541]    <= x541_in;                     
						a0_wr[542]    <= x542_in;                     
						a0_wr[543]    <= x543_in;                     
						a0_wr[544]    <= x544_in;                     
						a0_wr[545]    <= x545_in;                     
						a0_wr[546]    <= x546_in;                     
						a0_wr[547]    <= x547_in;                     
						a0_wr[548]    <= x548_in;                     
						a0_wr[549]    <= x549_in;                     
						a0_wr[550]    <= x550_in;                     
						a0_wr[551]    <= x551_in;                     
						a0_wr[552]    <= x552_in;                     
						a0_wr[553]    <= x553_in;                     
						a0_wr[554]    <= x554_in;                     
						a0_wr[555]    <= x555_in;                     
						a0_wr[556]    <= x556_in;                     
						a0_wr[557]    <= x557_in;                     
						a0_wr[558]    <= x558_in;                     
						a0_wr[559]    <= x559_in;                     
						a0_wr[560]    <= x560_in;                     
						a0_wr[561]    <= x561_in;                     
						a0_wr[562]    <= x562_in;                     
						a0_wr[563]    <= x563_in;                     
						a0_wr[564]    <= x564_in;                     
						a0_wr[565]    <= x565_in;                     
						a0_wr[566]    <= x566_in;                     
						a0_wr[567]    <= x567_in;                     
						a0_wr[568]    <= x568_in;                     
						a0_wr[569]    <= x569_in;                     
						a0_wr[570]    <= x570_in;                     
						a0_wr[571]    <= x571_in;                     
						a0_wr[572]    <= x572_in;                     
						a0_wr[573]    <= x573_in;                     
						a0_wr[574]    <= x574_in;                     
						a0_wr[575]    <= x575_in;                     
						a0_wr[576]    <= x576_in;                     
						a0_wr[577]    <= x577_in;                     
						a0_wr[578]    <= x578_in;                     
						a0_wr[579]    <= x579_in;                     
						a0_wr[580]    <= x580_in;                     
						a0_wr[581]    <= x581_in;                     
						a0_wr[582]    <= x582_in;                     
						a0_wr[583]    <= x583_in;                     
						a0_wr[584]    <= x584_in;                     
						a0_wr[585]    <= x585_in;                     
						a0_wr[586]    <= x586_in;                     
						a0_wr[587]    <= x587_in;                     
						a0_wr[588]    <= x588_in;                     
						a0_wr[589]    <= x589_in;                     
						a0_wr[590]    <= x590_in;                     
						a0_wr[591]    <= x591_in;                     
						a0_wr[592]    <= x592_in;                     
						a0_wr[593]    <= x593_in;                     
						a0_wr[594]    <= x594_in;                     
						a0_wr[595]    <= x595_in;                     
						a0_wr[596]    <= x596_in;                     
						a0_wr[597]    <= x597_in;                     
						a0_wr[598]    <= x598_in;                     
						a0_wr[599]    <= x599_in;                     
						a0_wr[600]    <= x600_in;                     
						a0_wr[601]    <= x601_in;                     
						a0_wr[602]    <= x602_in;                     
						a0_wr[603]    <= x603_in;                     
						a0_wr[604]    <= x604_in;                     
						a0_wr[605]    <= x605_in;                     
						a0_wr[606]    <= x606_in;                     
						a0_wr[607]    <= x607_in;                     
						a0_wr[608]    <= x608_in;                     
						a0_wr[609]    <= x609_in;                     
						a0_wr[610]    <= x610_in;                     
						a0_wr[611]    <= x611_in;                     
						a0_wr[612]    <= x612_in;                     
						a0_wr[613]    <= x613_in;                     
						a0_wr[614]    <= x614_in;                     
						a0_wr[615]    <= x615_in;                     
						a0_wr[616]    <= x616_in;                     
						a0_wr[617]    <= x617_in;                     
						a0_wr[618]    <= x618_in;                     
						a0_wr[619]    <= x619_in;                     
						a0_wr[620]    <= x620_in;                     
						a0_wr[621]    <= x621_in;                     
						a0_wr[622]    <= x622_in;                     
						a0_wr[623]    <= x623_in;                     
						a0_wr[624]    <= x624_in;                     
						a0_wr[625]    <= x625_in;                     
						a0_wr[626]    <= x626_in;                     
						a0_wr[627]    <= x627_in;                     
						a0_wr[628]    <= x628_in;                     
						a0_wr[629]    <= x629_in;                     
						a0_wr[630]    <= x630_in;                     
						a0_wr[631]    <= x631_in;                     
						a0_wr[632]    <= x632_in;                     
						a0_wr[633]    <= x633_in;                     
						a0_wr[634]    <= x634_in;                     
						a0_wr[635]    <= x635_in;                     
						a0_wr[636]    <= x636_in;                     
						a0_wr[637]    <= x637_in;                     
						a0_wr[638]    <= x638_in;                     
						a0_wr[639]    <= x639_in;                     
						a0_wr[640]    <= x640_in;                     
						a0_wr[641]    <= x641_in;                     
						a0_wr[642]    <= x642_in;                     
						a0_wr[643]    <= x643_in;                     
						a0_wr[644]    <= x644_in;                     
						a0_wr[645]    <= x645_in;                     
						a0_wr[646]    <= x646_in;                     
						a0_wr[647]    <= x647_in;                     
						a0_wr[648]    <= x648_in;                     
						a0_wr[649]    <= x649_in;                     
						a0_wr[650]    <= x650_in;                     
						a0_wr[651]    <= x651_in;                     
						a0_wr[652]    <= x652_in;                     
						a0_wr[653]    <= x653_in;                     
						a0_wr[654]    <= x654_in;                     
						a0_wr[655]    <= x655_in;                     
						a0_wr[656]    <= x656_in;                     
						a0_wr[657]    <= x657_in;                     
						a0_wr[658]    <= x658_in;                     
						a0_wr[659]    <= x659_in;                     
						a0_wr[660]    <= x660_in;                     
						a0_wr[661]    <= x661_in;                     
						a0_wr[662]    <= x662_in;                     
						a0_wr[663]    <= x663_in;                     
						a0_wr[664]    <= x664_in;                     
						a0_wr[665]    <= x665_in;                     
						a0_wr[666]    <= x666_in;                     
						a0_wr[667]    <= x667_in;                     
						a0_wr[668]    <= x668_in;                     
						a0_wr[669]    <= x669_in;                     
						a0_wr[670]    <= x670_in;                     
						a0_wr[671]    <= x671_in;                     
						a0_wr[672]    <= x672_in;                     
						a0_wr[673]    <= x673_in;                     
						a0_wr[674]    <= x674_in;                     
						a0_wr[675]    <= x675_in;                     
						a0_wr[676]    <= x676_in;                     
						a0_wr[677]    <= x677_in;                     
						a0_wr[678]    <= x678_in;                     
						a0_wr[679]    <= x679_in;                     
						a0_wr[680]    <= x680_in;                     
						a0_wr[681]    <= x681_in;                     
						a0_wr[682]    <= x682_in;                     
						a0_wr[683]    <= x683_in;                     
						a0_wr[684]    <= x684_in;                     
						a0_wr[685]    <= x685_in;                     
						a0_wr[686]    <= x686_in;                     
						a0_wr[687]    <= x687_in;                     
						a0_wr[688]    <= x688_in;                     
						a0_wr[689]    <= x689_in;                     
						a0_wr[690]    <= x690_in;                     
						a0_wr[691]    <= x691_in;                     
						a0_wr[692]    <= x692_in;                     
						a0_wr[693]    <= x693_in;                     
						a0_wr[694]    <= x694_in;                     
						a0_wr[695]    <= x695_in;                     
						a0_wr[696]    <= x696_in;                     
						a0_wr[697]    <= x697_in;                     
						a0_wr[698]    <= x698_in;                     
						a0_wr[699]    <= x699_in;                     
						a0_wr[700]    <= x700_in;                     
						a0_wr[701]    <= x701_in;                     
						a0_wr[702]    <= x702_in;                     
						a0_wr[703]    <= x703_in;                     
						a0_wr[704]    <= x704_in;                     
						a0_wr[705]    <= x705_in;                     
						a0_wr[706]    <= x706_in;                     
						a0_wr[707]    <= x707_in;                     
						a0_wr[708]    <= x708_in;                     
						a0_wr[709]    <= x709_in;                     
						a0_wr[710]    <= x710_in;                     
						a0_wr[711]    <= x711_in;                     
						a0_wr[712]    <= x712_in;                     
						a0_wr[713]    <= x713_in;                     
						a0_wr[714]    <= x714_in;                     
						a0_wr[715]    <= x715_in;                     
						a0_wr[716]    <= x716_in;                     
						a0_wr[717]    <= x717_in;                     
						a0_wr[718]    <= x718_in;                     
						a0_wr[719]    <= x719_in;                     
						a0_wr[720]    <= x720_in;                     
						a0_wr[721]    <= x721_in;                     
						a0_wr[722]    <= x722_in;                     
						a0_wr[723]    <= x723_in;                     
						a0_wr[724]    <= x724_in;                     
						a0_wr[725]    <= x725_in;                     
						a0_wr[726]    <= x726_in;                     
						a0_wr[727]    <= x727_in;                     
						a0_wr[728]    <= x728_in;                     
						a0_wr[729]    <= x729_in;                     
						a0_wr[730]    <= x730_in;                     
						a0_wr[731]    <= x731_in;                     
						a0_wr[732]    <= x732_in;                     
						a0_wr[733]    <= x733_in;                     
						a0_wr[734]    <= x734_in;                     
						a0_wr[735]    <= x735_in;                     
						a0_wr[736]    <= x736_in;                     
						a0_wr[737]    <= x737_in;                     
						a0_wr[738]    <= x738_in;                     
						a0_wr[739]    <= x739_in;                     
						a0_wr[740]    <= x740_in;                     
						a0_wr[741]    <= x741_in;                     
						a0_wr[742]    <= x742_in;                     
						a0_wr[743]    <= x743_in;                     
						a0_wr[744]    <= x744_in;                     
						a0_wr[745]    <= x745_in;                     
						a0_wr[746]    <= x746_in;                     
						a0_wr[747]    <= x747_in;                     
						a0_wr[748]    <= x748_in;                     
						a0_wr[749]    <= x749_in;                     
						a0_wr[750]    <= x750_in;                     
						a0_wr[751]    <= x751_in;                     
						a0_wr[752]    <= x752_in;                     
						a0_wr[753]    <= x753_in;                     
						a0_wr[754]    <= x754_in;                     
						a0_wr[755]    <= x755_in;                     
						a0_wr[756]    <= x756_in;                     
						a0_wr[757]    <= x757_in;                     
						a0_wr[758]    <= x758_in;                     
						a0_wr[759]    <= x759_in;                     
						a0_wr[760]    <= x760_in;                     
						a0_wr[761]    <= x761_in;                     
						a0_wr[762]    <= x762_in;                     
						a0_wr[763]    <= x763_in;                     
						a0_wr[764]    <= x764_in;                     
						a0_wr[765]    <= x765_in;                     
						a0_wr[766]    <= x766_in;                     
						a0_wr[767]    <= x767_in;                     
						a0_wr[768]    <= x768_in;                     
						a0_wr[769]    <= x769_in;                     
						a0_wr[770]    <= x770_in;                     
						a0_wr[771]    <= x771_in;                     
						a0_wr[772]    <= x772_in;                     
						a0_wr[773]    <= x773_in;                     
						a0_wr[774]    <= x774_in;                     
						a0_wr[775]    <= x775_in;                     
						a0_wr[776]    <= x776_in;                     
						a0_wr[777]    <= x777_in;                     
						a0_wr[778]    <= x778_in;                     
						a0_wr[779]    <= x779_in;                     
						a0_wr[780]    <= x780_in;                     
						a0_wr[781]    <= x781_in;                     
						a0_wr[782]    <= x782_in;                     
						a0_wr[783]    <= x783_in;                     
						a0_wr[784]    <= x784_in;                     
						a0_wr[785]    <= x785_in;                     
						a0_wr[786]    <= x786_in;                     
						a0_wr[787]    <= x787_in;                     
						a0_wr[788]    <= x788_in;                     
						a0_wr[789]    <= x789_in;                     
						a0_wr[790]    <= x790_in;                     
						a0_wr[791]    <= x791_in;                     
						a0_wr[792]    <= x792_in;                     
						a0_wr[793]    <= x793_in;                     
						a0_wr[794]    <= x794_in;                     
						a0_wr[795]    <= x795_in;                     
						a0_wr[796]    <= x796_in;                     
						a0_wr[797]    <= x797_in;                     
						a0_wr[798]    <= x798_in;                     
						a0_wr[799]    <= x799_in;                     
						a0_wr[800]    <= x800_in;                     
						a0_wr[801]    <= x801_in;                     
						a0_wr[802]    <= x802_in;                     
						a0_wr[803]    <= x803_in;                     
						a0_wr[804]    <= x804_in;                     
						a0_wr[805]    <= x805_in;                     
						a0_wr[806]    <= x806_in;                     
						a0_wr[807]    <= x807_in;                     
						a0_wr[808]    <= x808_in;                     
						a0_wr[809]    <= x809_in;                     
						a0_wr[810]    <= x810_in;                     
						a0_wr[811]    <= x811_in;                     
						a0_wr[812]    <= x812_in;                     
						a0_wr[813]    <= x813_in;                     
						a0_wr[814]    <= x814_in;                     
						a0_wr[815]    <= x815_in;                     
						a0_wr[816]    <= x816_in;                     
						a0_wr[817]    <= x817_in;                     
						a0_wr[818]    <= x818_in;                     
						a0_wr[819]    <= x819_in;                     
						a0_wr[820]    <= x820_in;                     
						a0_wr[821]    <= x821_in;                     
						a0_wr[822]    <= x822_in;                     
						a0_wr[823]    <= x823_in;                     
						a0_wr[824]    <= x824_in;                     
						a0_wr[825]    <= x825_in;                     
						a0_wr[826]    <= x826_in;                     
						a0_wr[827]    <= x827_in;                     
						a0_wr[828]    <= x828_in;                     
						a0_wr[829]    <= x829_in;                     
						a0_wr[830]    <= x830_in;                     
						a0_wr[831]    <= x831_in;                     
						a0_wr[832]    <= x832_in;                     
						a0_wr[833]    <= x833_in;                     
						a0_wr[834]    <= x834_in;                     
						a0_wr[835]    <= x835_in;                     
						a0_wr[836]    <= x836_in;                     
						a0_wr[837]    <= x837_in;                     
						a0_wr[838]    <= x838_in;                     
						a0_wr[839]    <= x839_in;                     
						a0_wr[840]    <= x840_in;                     
						a0_wr[841]    <= x841_in;                     
						a0_wr[842]    <= x842_in;                     
						a0_wr[843]    <= x843_in;                     
						a0_wr[844]    <= x844_in;                     
						a0_wr[845]    <= x845_in;                     
						a0_wr[846]    <= x846_in;                     
						a0_wr[847]    <= x847_in;                     
						a0_wr[848]    <= x848_in;                     
						a0_wr[849]    <= x849_in;                     
						a0_wr[850]    <= x850_in;                     
						a0_wr[851]    <= x851_in;                     
						a0_wr[852]    <= x852_in;                     
						a0_wr[853]    <= x853_in;                     
						a0_wr[854]    <= x854_in;                     
						a0_wr[855]    <= x855_in;                     
						a0_wr[856]    <= x856_in;                     
						a0_wr[857]    <= x857_in;                     
						a0_wr[858]    <= x858_in;                     
						a0_wr[859]    <= x859_in;                     
						a0_wr[860]    <= x860_in;                     
						a0_wr[861]    <= x861_in;                     
						a0_wr[862]    <= x862_in;                     
						a0_wr[863]    <= x863_in;                     
						a0_wr[864]    <= x864_in;                     
						a0_wr[865]    <= x865_in;                     
						a0_wr[866]    <= x866_in;                     
						a0_wr[867]    <= x867_in;                     
						a0_wr[868]    <= x868_in;                     
						a0_wr[869]    <= x869_in;                     
						a0_wr[870]    <= x870_in;                     
						a0_wr[871]    <= x871_in;                     
						a0_wr[872]    <= x872_in;                     
						a0_wr[873]    <= x873_in;                     
						a0_wr[874]    <= x874_in;                     
						a0_wr[875]    <= x875_in;                     
						a0_wr[876]    <= x876_in;                     
						a0_wr[877]    <= x877_in;                     
						a0_wr[878]    <= x878_in;                     
						a0_wr[879]    <= x879_in;                     
						a0_wr[880]    <= x880_in;                     
						a0_wr[881]    <= x881_in;                     
						a0_wr[882]    <= x882_in;                     
						a0_wr[883]    <= x883_in;                     
						a0_wr[884]    <= x884_in;                     
						a0_wr[885]    <= x885_in;                     
						a0_wr[886]    <= x886_in;                     
						a0_wr[887]    <= x887_in;                     
						a0_wr[888]    <= x888_in;                     
						a0_wr[889]    <= x889_in;                     
						a0_wr[890]    <= x890_in;                     
						a0_wr[891]    <= x891_in;                     
						a0_wr[892]    <= x892_in;                     
						a0_wr[893]    <= x893_in;                     
						a0_wr[894]    <= x894_in;                     
						a0_wr[895]    <= x895_in;                     
						a0_wr[896]    <= x896_in;                     
						a0_wr[897]    <= x897_in;                     
						a0_wr[898]    <= x898_in;                     
						a0_wr[899]    <= x899_in;                     
						a0_wr[900]    <= x900_in;                     
						a0_wr[901]    <= x901_in;                     
						a0_wr[902]    <= x902_in;                     
						a0_wr[903]    <= x903_in;                     
						a0_wr[904]    <= x904_in;                     
						a0_wr[905]    <= x905_in;                     
						a0_wr[906]    <= x906_in;                     
						a0_wr[907]    <= x907_in;                     
						a0_wr[908]    <= x908_in;                     
						a0_wr[909]    <= x909_in;                     
						a0_wr[910]    <= x910_in;                     
						a0_wr[911]    <= x911_in;                     
						a0_wr[912]    <= x912_in;                     
						a0_wr[913]    <= x913_in;                     
						a0_wr[914]    <= x914_in;                     
						a0_wr[915]    <= x915_in;                     
						a0_wr[916]    <= x916_in;                     
						a0_wr[917]    <= x917_in;                     
						a0_wr[918]    <= x918_in;                     
						a0_wr[919]    <= x919_in;                     
						a0_wr[920]    <= x920_in;                     
						a0_wr[921]    <= x921_in;                     
						a0_wr[922]    <= x922_in;                     
						a0_wr[923]    <= x923_in;                     
						a0_wr[924]    <= x924_in;                     
						a0_wr[925]    <= x925_in;                     
						a0_wr[926]    <= x926_in;                     
						a0_wr[927]    <= x927_in;                     
						a0_wr[928]    <= x928_in;                     
						a0_wr[929]    <= x929_in;                     
						a0_wr[930]    <= x930_in;                     
						a0_wr[931]    <= x931_in;                     
						a0_wr[932]    <= x932_in;                     
						a0_wr[933]    <= x933_in;                     
						a0_wr[934]    <= x934_in;                     
						a0_wr[935]    <= x935_in;                     
						a0_wr[936]    <= x936_in;                     
						a0_wr[937]    <= x937_in;                     
						a0_wr[938]    <= x938_in;                     
						a0_wr[939]    <= x939_in;                     
						a0_wr[940]    <= x940_in;                     
						a0_wr[941]    <= x941_in;                     
						a0_wr[942]    <= x942_in;                     
						a0_wr[943]    <= x943_in;                     
						a0_wr[944]    <= x944_in;                     
						a0_wr[945]    <= x945_in;                     
						a0_wr[946]    <= x946_in;                     
						a0_wr[947]    <= x947_in;                     
						a0_wr[948]    <= x948_in;                     
						a0_wr[949]    <= x949_in;                     
						a0_wr[950]    <= x950_in;                     
						a0_wr[951]    <= x951_in;                     
						a0_wr[952]    <= x952_in;                     
						a0_wr[953]    <= x953_in;                     
						a0_wr[954]    <= x954_in;                     
						a0_wr[955]    <= x955_in;                     
						a0_wr[956]    <= x956_in;                     
						a0_wr[957]    <= x957_in;                     
						a0_wr[958]    <= x958_in;                     
						a0_wr[959]    <= x959_in;                     
						a0_wr[960]    <= x960_in;                     
						a0_wr[961]    <= x961_in;                     
						a0_wr[962]    <= x962_in;                     
						a0_wr[963]    <= x963_in;                     
						a0_wr[964]    <= x964_in;                     
						a0_wr[965]    <= x965_in;                     
						a0_wr[966]    <= x966_in;                     
						a0_wr[967]    <= x967_in;                     
						a0_wr[968]    <= x968_in;                     
						a0_wr[969]    <= x969_in;                     
						a0_wr[970]    <= x970_in;                     
						a0_wr[971]    <= x971_in;                     
						a0_wr[972]    <= x972_in;                     
						a0_wr[973]    <= x973_in;                     
						a0_wr[974]    <= x974_in;                     
						a0_wr[975]    <= x975_in;                     
						a0_wr[976]    <= x976_in;                     
						a0_wr[977]    <= x977_in;                     
						a0_wr[978]    <= x978_in;                     
						a0_wr[979]    <= x979_in;                     
						a0_wr[980]    <= x980_in;                     
						a0_wr[981]    <= x981_in;                     
						a0_wr[982]    <= x982_in;                     
						a0_wr[983]    <= x983_in;                     
						a0_wr[984]    <= x984_in;                     
						a0_wr[985]    <= x985_in;                     
						a0_wr[986]    <= x986_in;                     
						a0_wr[987]    <= x987_in;                     
						a0_wr[988]    <= x988_in;                     
						a0_wr[989]    <= x989_in;                     
						a0_wr[990]    <= x990_in;                     
						a0_wr[991]    <= x991_in;                     
						a0_wr[992]    <= x992_in;                     
						a0_wr[993]    <= x993_in;                     
						a0_wr[994]    <= x994_in;                     
						a0_wr[995]    <= x995_in;                     
						a0_wr[996]    <= x996_in;                     
						a0_wr[997]    <= x997_in;                     
						a0_wr[998]    <= x998_in;                     
						a0_wr[999]    <= x999_in;                     
						a0_wr[1000]   <= x1000_in;                    
						a0_wr[1001]   <= x1001_in;                    
						a0_wr[1002]   <= x1002_in;                    
						a0_wr[1003]   <= x1003_in;                    
						a0_wr[1004]   <= x1004_in;                    
						a0_wr[1005]   <= x1005_in;                    
						a0_wr[1006]   <= x1006_in;                    
						a0_wr[1007]   <= x1007_in;                    
						a0_wr[1008]   <= x1008_in;                    
						a0_wr[1009]   <= x1009_in;                    
						a0_wr[1010]   <= x1010_in;                    
						a0_wr[1011]   <= x1011_in;                    
						a0_wr[1012]   <= x1012_in;                    
						a0_wr[1013]   <= x1013_in;                    
						a0_wr[1014]   <= x1014_in;                    
						a0_wr[1015]   <= x1015_in;                    
						a0_wr[1016]   <= x1016_in;                    
						a0_wr[1017]   <= x1017_in;                    
						a0_wr[1018]   <= x1018_in;                    
						a0_wr[1019]   <= x1019_in;                    
						a0_wr[1020]   <= x1020_in;                    
						a0_wr[1021]   <= x1021_in;                    
						a0_wr[1022]   <= x1022_in;                    
						a0_wr[1023]   <= x1023_in;                    
					end
				end
			end

		//--- radix stage 0
			radix2 #(.width(width)) rd_st0_0   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[0]), .rdlo_in(a0_wr[512]),  .coef_in(coef[0]), .rdup_out(a1_wr[0]), .rdlo_out(a1_wr[512]));
			radix2 #(.width(width)) rd_st0_1   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[1]), .rdlo_in(a0_wr[513]),  .coef_in(coef[1]), .rdup_out(a1_wr[1]), .rdlo_out(a1_wr[513]));
			radix2 #(.width(width)) rd_st0_2   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[2]), .rdlo_in(a0_wr[514]),  .coef_in(coef[2]), .rdup_out(a1_wr[2]), .rdlo_out(a1_wr[514]));
			radix2 #(.width(width)) rd_st0_3   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[3]), .rdlo_in(a0_wr[515]),  .coef_in(coef[3]), .rdup_out(a1_wr[3]), .rdlo_out(a1_wr[515]));
			radix2 #(.width(width)) rd_st0_4   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[4]), .rdlo_in(a0_wr[516]),  .coef_in(coef[4]), .rdup_out(a1_wr[4]), .rdlo_out(a1_wr[516]));
			radix2 #(.width(width)) rd_st0_5   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[5]), .rdlo_in(a0_wr[517]),  .coef_in(coef[5]), .rdup_out(a1_wr[5]), .rdlo_out(a1_wr[517]));
			radix2 #(.width(width)) rd_st0_6   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[6]), .rdlo_in(a0_wr[518]),  .coef_in(coef[6]), .rdup_out(a1_wr[6]), .rdlo_out(a1_wr[518]));
			radix2 #(.width(width)) rd_st0_7   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[7]), .rdlo_in(a0_wr[519]),  .coef_in(coef[7]), .rdup_out(a1_wr[7]), .rdlo_out(a1_wr[519]));
			radix2 #(.width(width)) rd_st0_8   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[8]), .rdlo_in(a0_wr[520]),  .coef_in(coef[8]), .rdup_out(a1_wr[8]), .rdlo_out(a1_wr[520]));
			radix2 #(.width(width)) rd_st0_9   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[9]), .rdlo_in(a0_wr[521]),  .coef_in(coef[9]), .rdup_out(a1_wr[9]), .rdlo_out(a1_wr[521]));
			radix2 #(.width(width)) rd_st0_10  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[10]), .rdlo_in(a0_wr[522]),  .coef_in(coef[10]), .rdup_out(a1_wr[10]), .rdlo_out(a1_wr[522]));
			radix2 #(.width(width)) rd_st0_11  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[11]), .rdlo_in(a0_wr[523]),  .coef_in(coef[11]), .rdup_out(a1_wr[11]), .rdlo_out(a1_wr[523]));
			radix2 #(.width(width)) rd_st0_12  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[12]), .rdlo_in(a0_wr[524]),  .coef_in(coef[12]), .rdup_out(a1_wr[12]), .rdlo_out(a1_wr[524]));
			radix2 #(.width(width)) rd_st0_13  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[13]), .rdlo_in(a0_wr[525]),  .coef_in(coef[13]), .rdup_out(a1_wr[13]), .rdlo_out(a1_wr[525]));
			radix2 #(.width(width)) rd_st0_14  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[14]), .rdlo_in(a0_wr[526]),  .coef_in(coef[14]), .rdup_out(a1_wr[14]), .rdlo_out(a1_wr[526]));
			radix2 #(.width(width)) rd_st0_15  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[15]), .rdlo_in(a0_wr[527]),  .coef_in(coef[15]), .rdup_out(a1_wr[15]), .rdlo_out(a1_wr[527]));
			radix2 #(.width(width)) rd_st0_16  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[16]), .rdlo_in(a0_wr[528]),  .coef_in(coef[16]), .rdup_out(a1_wr[16]), .rdlo_out(a1_wr[528]));
			radix2 #(.width(width)) rd_st0_17  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[17]), .rdlo_in(a0_wr[529]),  .coef_in(coef[17]), .rdup_out(a1_wr[17]), .rdlo_out(a1_wr[529]));
			radix2 #(.width(width)) rd_st0_18  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[18]), .rdlo_in(a0_wr[530]),  .coef_in(coef[18]), .rdup_out(a1_wr[18]), .rdlo_out(a1_wr[530]));
			radix2 #(.width(width)) rd_st0_19  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[19]), .rdlo_in(a0_wr[531]),  .coef_in(coef[19]), .rdup_out(a1_wr[19]), .rdlo_out(a1_wr[531]));
			radix2 #(.width(width)) rd_st0_20  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[20]), .rdlo_in(a0_wr[532]),  .coef_in(coef[20]), .rdup_out(a1_wr[20]), .rdlo_out(a1_wr[532]));
			radix2 #(.width(width)) rd_st0_21  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[21]), .rdlo_in(a0_wr[533]),  .coef_in(coef[21]), .rdup_out(a1_wr[21]), .rdlo_out(a1_wr[533]));
			radix2 #(.width(width)) rd_st0_22  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[22]), .rdlo_in(a0_wr[534]),  .coef_in(coef[22]), .rdup_out(a1_wr[22]), .rdlo_out(a1_wr[534]));
			radix2 #(.width(width)) rd_st0_23  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[23]), .rdlo_in(a0_wr[535]),  .coef_in(coef[23]), .rdup_out(a1_wr[23]), .rdlo_out(a1_wr[535]));
			radix2 #(.width(width)) rd_st0_24  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[24]), .rdlo_in(a0_wr[536]),  .coef_in(coef[24]), .rdup_out(a1_wr[24]), .rdlo_out(a1_wr[536]));
			radix2 #(.width(width)) rd_st0_25  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[25]), .rdlo_in(a0_wr[537]),  .coef_in(coef[25]), .rdup_out(a1_wr[25]), .rdlo_out(a1_wr[537]));
			radix2 #(.width(width)) rd_st0_26  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[26]), .rdlo_in(a0_wr[538]),  .coef_in(coef[26]), .rdup_out(a1_wr[26]), .rdlo_out(a1_wr[538]));
			radix2 #(.width(width)) rd_st0_27  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[27]), .rdlo_in(a0_wr[539]),  .coef_in(coef[27]), .rdup_out(a1_wr[27]), .rdlo_out(a1_wr[539]));
			radix2 #(.width(width)) rd_st0_28  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[28]), .rdlo_in(a0_wr[540]),  .coef_in(coef[28]), .rdup_out(a1_wr[28]), .rdlo_out(a1_wr[540]));
			radix2 #(.width(width)) rd_st0_29  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[29]), .rdlo_in(a0_wr[541]),  .coef_in(coef[29]), .rdup_out(a1_wr[29]), .rdlo_out(a1_wr[541]));
			radix2 #(.width(width)) rd_st0_30  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[30]), .rdlo_in(a0_wr[542]),  .coef_in(coef[30]), .rdup_out(a1_wr[30]), .rdlo_out(a1_wr[542]));
			radix2 #(.width(width)) rd_st0_31  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[31]), .rdlo_in(a0_wr[543]),  .coef_in(coef[31]), .rdup_out(a1_wr[31]), .rdlo_out(a1_wr[543]));
			radix2 #(.width(width)) rd_st0_32  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[32]), .rdlo_in(a0_wr[544]),  .coef_in(coef[32]), .rdup_out(a1_wr[32]), .rdlo_out(a1_wr[544]));
			radix2 #(.width(width)) rd_st0_33  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[33]), .rdlo_in(a0_wr[545]),  .coef_in(coef[33]), .rdup_out(a1_wr[33]), .rdlo_out(a1_wr[545]));
			radix2 #(.width(width)) rd_st0_34  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[34]), .rdlo_in(a0_wr[546]),  .coef_in(coef[34]), .rdup_out(a1_wr[34]), .rdlo_out(a1_wr[546]));
			radix2 #(.width(width)) rd_st0_35  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[35]), .rdlo_in(a0_wr[547]),  .coef_in(coef[35]), .rdup_out(a1_wr[35]), .rdlo_out(a1_wr[547]));
			radix2 #(.width(width)) rd_st0_36  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[36]), .rdlo_in(a0_wr[548]),  .coef_in(coef[36]), .rdup_out(a1_wr[36]), .rdlo_out(a1_wr[548]));
			radix2 #(.width(width)) rd_st0_37  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[37]), .rdlo_in(a0_wr[549]),  .coef_in(coef[37]), .rdup_out(a1_wr[37]), .rdlo_out(a1_wr[549]));
			radix2 #(.width(width)) rd_st0_38  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[38]), .rdlo_in(a0_wr[550]),  .coef_in(coef[38]), .rdup_out(a1_wr[38]), .rdlo_out(a1_wr[550]));
			radix2 #(.width(width)) rd_st0_39  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[39]), .rdlo_in(a0_wr[551]),  .coef_in(coef[39]), .rdup_out(a1_wr[39]), .rdlo_out(a1_wr[551]));
			radix2 #(.width(width)) rd_st0_40  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[40]), .rdlo_in(a0_wr[552]),  .coef_in(coef[40]), .rdup_out(a1_wr[40]), .rdlo_out(a1_wr[552]));
			radix2 #(.width(width)) rd_st0_41  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[41]), .rdlo_in(a0_wr[553]),  .coef_in(coef[41]), .rdup_out(a1_wr[41]), .rdlo_out(a1_wr[553]));
			radix2 #(.width(width)) rd_st0_42  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[42]), .rdlo_in(a0_wr[554]),  .coef_in(coef[42]), .rdup_out(a1_wr[42]), .rdlo_out(a1_wr[554]));
			radix2 #(.width(width)) rd_st0_43  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[43]), .rdlo_in(a0_wr[555]),  .coef_in(coef[43]), .rdup_out(a1_wr[43]), .rdlo_out(a1_wr[555]));
			radix2 #(.width(width)) rd_st0_44  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[44]), .rdlo_in(a0_wr[556]),  .coef_in(coef[44]), .rdup_out(a1_wr[44]), .rdlo_out(a1_wr[556]));
			radix2 #(.width(width)) rd_st0_45  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[45]), .rdlo_in(a0_wr[557]),  .coef_in(coef[45]), .rdup_out(a1_wr[45]), .rdlo_out(a1_wr[557]));
			radix2 #(.width(width)) rd_st0_46  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[46]), .rdlo_in(a0_wr[558]),  .coef_in(coef[46]), .rdup_out(a1_wr[46]), .rdlo_out(a1_wr[558]));
			radix2 #(.width(width)) rd_st0_47  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[47]), .rdlo_in(a0_wr[559]),  .coef_in(coef[47]), .rdup_out(a1_wr[47]), .rdlo_out(a1_wr[559]));
			radix2 #(.width(width)) rd_st0_48  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[48]), .rdlo_in(a0_wr[560]),  .coef_in(coef[48]), .rdup_out(a1_wr[48]), .rdlo_out(a1_wr[560]));
			radix2 #(.width(width)) rd_st0_49  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[49]), .rdlo_in(a0_wr[561]),  .coef_in(coef[49]), .rdup_out(a1_wr[49]), .rdlo_out(a1_wr[561]));
			radix2 #(.width(width)) rd_st0_50  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[50]), .rdlo_in(a0_wr[562]),  .coef_in(coef[50]), .rdup_out(a1_wr[50]), .rdlo_out(a1_wr[562]));
			radix2 #(.width(width)) rd_st0_51  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[51]), .rdlo_in(a0_wr[563]),  .coef_in(coef[51]), .rdup_out(a1_wr[51]), .rdlo_out(a1_wr[563]));
			radix2 #(.width(width)) rd_st0_52  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[52]), .rdlo_in(a0_wr[564]),  .coef_in(coef[52]), .rdup_out(a1_wr[52]), .rdlo_out(a1_wr[564]));
			radix2 #(.width(width)) rd_st0_53  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[53]), .rdlo_in(a0_wr[565]),  .coef_in(coef[53]), .rdup_out(a1_wr[53]), .rdlo_out(a1_wr[565]));
			radix2 #(.width(width)) rd_st0_54  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[54]), .rdlo_in(a0_wr[566]),  .coef_in(coef[54]), .rdup_out(a1_wr[54]), .rdlo_out(a1_wr[566]));
			radix2 #(.width(width)) rd_st0_55  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[55]), .rdlo_in(a0_wr[567]),  .coef_in(coef[55]), .rdup_out(a1_wr[55]), .rdlo_out(a1_wr[567]));
			radix2 #(.width(width)) rd_st0_56  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[56]), .rdlo_in(a0_wr[568]),  .coef_in(coef[56]), .rdup_out(a1_wr[56]), .rdlo_out(a1_wr[568]));
			radix2 #(.width(width)) rd_st0_57  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[57]), .rdlo_in(a0_wr[569]),  .coef_in(coef[57]), .rdup_out(a1_wr[57]), .rdlo_out(a1_wr[569]));
			radix2 #(.width(width)) rd_st0_58  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[58]), .rdlo_in(a0_wr[570]),  .coef_in(coef[58]), .rdup_out(a1_wr[58]), .rdlo_out(a1_wr[570]));
			radix2 #(.width(width)) rd_st0_59  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[59]), .rdlo_in(a0_wr[571]),  .coef_in(coef[59]), .rdup_out(a1_wr[59]), .rdlo_out(a1_wr[571]));
			radix2 #(.width(width)) rd_st0_60  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[60]), .rdlo_in(a0_wr[572]),  .coef_in(coef[60]), .rdup_out(a1_wr[60]), .rdlo_out(a1_wr[572]));
			radix2 #(.width(width)) rd_st0_61  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[61]), .rdlo_in(a0_wr[573]),  .coef_in(coef[61]), .rdup_out(a1_wr[61]), .rdlo_out(a1_wr[573]));
			radix2 #(.width(width)) rd_st0_62  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[62]), .rdlo_in(a0_wr[574]),  .coef_in(coef[62]), .rdup_out(a1_wr[62]), .rdlo_out(a1_wr[574]));
			radix2 #(.width(width)) rd_st0_63  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[63]), .rdlo_in(a0_wr[575]),  .coef_in(coef[63]), .rdup_out(a1_wr[63]), .rdlo_out(a1_wr[575]));
			radix2 #(.width(width)) rd_st0_64  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[64]), .rdlo_in(a0_wr[576]),  .coef_in(coef[64]), .rdup_out(a1_wr[64]), .rdlo_out(a1_wr[576]));
			radix2 #(.width(width)) rd_st0_65  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[65]), .rdlo_in(a0_wr[577]),  .coef_in(coef[65]), .rdup_out(a1_wr[65]), .rdlo_out(a1_wr[577]));
			radix2 #(.width(width)) rd_st0_66  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[66]), .rdlo_in(a0_wr[578]),  .coef_in(coef[66]), .rdup_out(a1_wr[66]), .rdlo_out(a1_wr[578]));
			radix2 #(.width(width)) rd_st0_67  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[67]), .rdlo_in(a0_wr[579]),  .coef_in(coef[67]), .rdup_out(a1_wr[67]), .rdlo_out(a1_wr[579]));
			radix2 #(.width(width)) rd_st0_68  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[68]), .rdlo_in(a0_wr[580]),  .coef_in(coef[68]), .rdup_out(a1_wr[68]), .rdlo_out(a1_wr[580]));
			radix2 #(.width(width)) rd_st0_69  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[69]), .rdlo_in(a0_wr[581]),  .coef_in(coef[69]), .rdup_out(a1_wr[69]), .rdlo_out(a1_wr[581]));
			radix2 #(.width(width)) rd_st0_70  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[70]), .rdlo_in(a0_wr[582]),  .coef_in(coef[70]), .rdup_out(a1_wr[70]), .rdlo_out(a1_wr[582]));
			radix2 #(.width(width)) rd_st0_71  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[71]), .rdlo_in(a0_wr[583]),  .coef_in(coef[71]), .rdup_out(a1_wr[71]), .rdlo_out(a1_wr[583]));
			radix2 #(.width(width)) rd_st0_72  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[72]), .rdlo_in(a0_wr[584]),  .coef_in(coef[72]), .rdup_out(a1_wr[72]), .rdlo_out(a1_wr[584]));
			radix2 #(.width(width)) rd_st0_73  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[73]), .rdlo_in(a0_wr[585]),  .coef_in(coef[73]), .rdup_out(a1_wr[73]), .rdlo_out(a1_wr[585]));
			radix2 #(.width(width)) rd_st0_74  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[74]), .rdlo_in(a0_wr[586]),  .coef_in(coef[74]), .rdup_out(a1_wr[74]), .rdlo_out(a1_wr[586]));
			radix2 #(.width(width)) rd_st0_75  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[75]), .rdlo_in(a0_wr[587]),  .coef_in(coef[75]), .rdup_out(a1_wr[75]), .rdlo_out(a1_wr[587]));
			radix2 #(.width(width)) rd_st0_76  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[76]), .rdlo_in(a0_wr[588]),  .coef_in(coef[76]), .rdup_out(a1_wr[76]), .rdlo_out(a1_wr[588]));
			radix2 #(.width(width)) rd_st0_77  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[77]), .rdlo_in(a0_wr[589]),  .coef_in(coef[77]), .rdup_out(a1_wr[77]), .rdlo_out(a1_wr[589]));
			radix2 #(.width(width)) rd_st0_78  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[78]), .rdlo_in(a0_wr[590]),  .coef_in(coef[78]), .rdup_out(a1_wr[78]), .rdlo_out(a1_wr[590]));
			radix2 #(.width(width)) rd_st0_79  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[79]), .rdlo_in(a0_wr[591]),  .coef_in(coef[79]), .rdup_out(a1_wr[79]), .rdlo_out(a1_wr[591]));
			radix2 #(.width(width)) rd_st0_80  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[80]), .rdlo_in(a0_wr[592]),  .coef_in(coef[80]), .rdup_out(a1_wr[80]), .rdlo_out(a1_wr[592]));
			radix2 #(.width(width)) rd_st0_81  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[81]), .rdlo_in(a0_wr[593]),  .coef_in(coef[81]), .rdup_out(a1_wr[81]), .rdlo_out(a1_wr[593]));
			radix2 #(.width(width)) rd_st0_82  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[82]), .rdlo_in(a0_wr[594]),  .coef_in(coef[82]), .rdup_out(a1_wr[82]), .rdlo_out(a1_wr[594]));
			radix2 #(.width(width)) rd_st0_83  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[83]), .rdlo_in(a0_wr[595]),  .coef_in(coef[83]), .rdup_out(a1_wr[83]), .rdlo_out(a1_wr[595]));
			radix2 #(.width(width)) rd_st0_84  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[84]), .rdlo_in(a0_wr[596]),  .coef_in(coef[84]), .rdup_out(a1_wr[84]), .rdlo_out(a1_wr[596]));
			radix2 #(.width(width)) rd_st0_85  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[85]), .rdlo_in(a0_wr[597]),  .coef_in(coef[85]), .rdup_out(a1_wr[85]), .rdlo_out(a1_wr[597]));
			radix2 #(.width(width)) rd_st0_86  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[86]), .rdlo_in(a0_wr[598]),  .coef_in(coef[86]), .rdup_out(a1_wr[86]), .rdlo_out(a1_wr[598]));
			radix2 #(.width(width)) rd_st0_87  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[87]), .rdlo_in(a0_wr[599]),  .coef_in(coef[87]), .rdup_out(a1_wr[87]), .rdlo_out(a1_wr[599]));
			radix2 #(.width(width)) rd_st0_88  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[88]), .rdlo_in(a0_wr[600]),  .coef_in(coef[88]), .rdup_out(a1_wr[88]), .rdlo_out(a1_wr[600]));
			radix2 #(.width(width)) rd_st0_89  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[89]), .rdlo_in(a0_wr[601]),  .coef_in(coef[89]), .rdup_out(a1_wr[89]), .rdlo_out(a1_wr[601]));
			radix2 #(.width(width)) rd_st0_90  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[90]), .rdlo_in(a0_wr[602]),  .coef_in(coef[90]), .rdup_out(a1_wr[90]), .rdlo_out(a1_wr[602]));
			radix2 #(.width(width)) rd_st0_91  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[91]), .rdlo_in(a0_wr[603]),  .coef_in(coef[91]), .rdup_out(a1_wr[91]), .rdlo_out(a1_wr[603]));
			radix2 #(.width(width)) rd_st0_92  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[92]), .rdlo_in(a0_wr[604]),  .coef_in(coef[92]), .rdup_out(a1_wr[92]), .rdlo_out(a1_wr[604]));
			radix2 #(.width(width)) rd_st0_93  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[93]), .rdlo_in(a0_wr[605]),  .coef_in(coef[93]), .rdup_out(a1_wr[93]), .rdlo_out(a1_wr[605]));
			radix2 #(.width(width)) rd_st0_94  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[94]), .rdlo_in(a0_wr[606]),  .coef_in(coef[94]), .rdup_out(a1_wr[94]), .rdlo_out(a1_wr[606]));
			radix2 #(.width(width)) rd_st0_95  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[95]), .rdlo_in(a0_wr[607]),  .coef_in(coef[95]), .rdup_out(a1_wr[95]), .rdlo_out(a1_wr[607]));
			radix2 #(.width(width)) rd_st0_96  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[96]), .rdlo_in(a0_wr[608]),  .coef_in(coef[96]), .rdup_out(a1_wr[96]), .rdlo_out(a1_wr[608]));
			radix2 #(.width(width)) rd_st0_97  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[97]), .rdlo_in(a0_wr[609]),  .coef_in(coef[97]), .rdup_out(a1_wr[97]), .rdlo_out(a1_wr[609]));
			radix2 #(.width(width)) rd_st0_98  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[98]), .rdlo_in(a0_wr[610]),  .coef_in(coef[98]), .rdup_out(a1_wr[98]), .rdlo_out(a1_wr[610]));
			radix2 #(.width(width)) rd_st0_99  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[99]), .rdlo_in(a0_wr[611]),  .coef_in(coef[99]), .rdup_out(a1_wr[99]), .rdlo_out(a1_wr[611]));
			radix2 #(.width(width)) rd_st0_100  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[100]), .rdlo_in(a0_wr[612]),  .coef_in(coef[100]), .rdup_out(a1_wr[100]), .rdlo_out(a1_wr[612]));
			radix2 #(.width(width)) rd_st0_101  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[101]), .rdlo_in(a0_wr[613]),  .coef_in(coef[101]), .rdup_out(a1_wr[101]), .rdlo_out(a1_wr[613]));
			radix2 #(.width(width)) rd_st0_102  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[102]), .rdlo_in(a0_wr[614]),  .coef_in(coef[102]), .rdup_out(a1_wr[102]), .rdlo_out(a1_wr[614]));
			radix2 #(.width(width)) rd_st0_103  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[103]), .rdlo_in(a0_wr[615]),  .coef_in(coef[103]), .rdup_out(a1_wr[103]), .rdlo_out(a1_wr[615]));
			radix2 #(.width(width)) rd_st0_104  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[104]), .rdlo_in(a0_wr[616]),  .coef_in(coef[104]), .rdup_out(a1_wr[104]), .rdlo_out(a1_wr[616]));
			radix2 #(.width(width)) rd_st0_105  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[105]), .rdlo_in(a0_wr[617]),  .coef_in(coef[105]), .rdup_out(a1_wr[105]), .rdlo_out(a1_wr[617]));
			radix2 #(.width(width)) rd_st0_106  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[106]), .rdlo_in(a0_wr[618]),  .coef_in(coef[106]), .rdup_out(a1_wr[106]), .rdlo_out(a1_wr[618]));
			radix2 #(.width(width)) rd_st0_107  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[107]), .rdlo_in(a0_wr[619]),  .coef_in(coef[107]), .rdup_out(a1_wr[107]), .rdlo_out(a1_wr[619]));
			radix2 #(.width(width)) rd_st0_108  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[108]), .rdlo_in(a0_wr[620]),  .coef_in(coef[108]), .rdup_out(a1_wr[108]), .rdlo_out(a1_wr[620]));
			radix2 #(.width(width)) rd_st0_109  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[109]), .rdlo_in(a0_wr[621]),  .coef_in(coef[109]), .rdup_out(a1_wr[109]), .rdlo_out(a1_wr[621]));
			radix2 #(.width(width)) rd_st0_110  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[110]), .rdlo_in(a0_wr[622]),  .coef_in(coef[110]), .rdup_out(a1_wr[110]), .rdlo_out(a1_wr[622]));
			radix2 #(.width(width)) rd_st0_111  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[111]), .rdlo_in(a0_wr[623]),  .coef_in(coef[111]), .rdup_out(a1_wr[111]), .rdlo_out(a1_wr[623]));
			radix2 #(.width(width)) rd_st0_112  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[112]), .rdlo_in(a0_wr[624]),  .coef_in(coef[112]), .rdup_out(a1_wr[112]), .rdlo_out(a1_wr[624]));
			radix2 #(.width(width)) rd_st0_113  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[113]), .rdlo_in(a0_wr[625]),  .coef_in(coef[113]), .rdup_out(a1_wr[113]), .rdlo_out(a1_wr[625]));
			radix2 #(.width(width)) rd_st0_114  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[114]), .rdlo_in(a0_wr[626]),  .coef_in(coef[114]), .rdup_out(a1_wr[114]), .rdlo_out(a1_wr[626]));
			radix2 #(.width(width)) rd_st0_115  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[115]), .rdlo_in(a0_wr[627]),  .coef_in(coef[115]), .rdup_out(a1_wr[115]), .rdlo_out(a1_wr[627]));
			radix2 #(.width(width)) rd_st0_116  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[116]), .rdlo_in(a0_wr[628]),  .coef_in(coef[116]), .rdup_out(a1_wr[116]), .rdlo_out(a1_wr[628]));
			radix2 #(.width(width)) rd_st0_117  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[117]), .rdlo_in(a0_wr[629]),  .coef_in(coef[117]), .rdup_out(a1_wr[117]), .rdlo_out(a1_wr[629]));
			radix2 #(.width(width)) rd_st0_118  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[118]), .rdlo_in(a0_wr[630]),  .coef_in(coef[118]), .rdup_out(a1_wr[118]), .rdlo_out(a1_wr[630]));
			radix2 #(.width(width)) rd_st0_119  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[119]), .rdlo_in(a0_wr[631]),  .coef_in(coef[119]), .rdup_out(a1_wr[119]), .rdlo_out(a1_wr[631]));
			radix2 #(.width(width)) rd_st0_120  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[120]), .rdlo_in(a0_wr[632]),  .coef_in(coef[120]), .rdup_out(a1_wr[120]), .rdlo_out(a1_wr[632]));
			radix2 #(.width(width)) rd_st0_121  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[121]), .rdlo_in(a0_wr[633]),  .coef_in(coef[121]), .rdup_out(a1_wr[121]), .rdlo_out(a1_wr[633]));
			radix2 #(.width(width)) rd_st0_122  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[122]), .rdlo_in(a0_wr[634]),  .coef_in(coef[122]), .rdup_out(a1_wr[122]), .rdlo_out(a1_wr[634]));
			radix2 #(.width(width)) rd_st0_123  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[123]), .rdlo_in(a0_wr[635]),  .coef_in(coef[123]), .rdup_out(a1_wr[123]), .rdlo_out(a1_wr[635]));
			radix2 #(.width(width)) rd_st0_124  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[124]), .rdlo_in(a0_wr[636]),  .coef_in(coef[124]), .rdup_out(a1_wr[124]), .rdlo_out(a1_wr[636]));
			radix2 #(.width(width)) rd_st0_125  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[125]), .rdlo_in(a0_wr[637]),  .coef_in(coef[125]), .rdup_out(a1_wr[125]), .rdlo_out(a1_wr[637]));
			radix2 #(.width(width)) rd_st0_126  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[126]), .rdlo_in(a0_wr[638]),  .coef_in(coef[126]), .rdup_out(a1_wr[126]), .rdlo_out(a1_wr[638]));
			radix2 #(.width(width)) rd_st0_127  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[127]), .rdlo_in(a0_wr[639]),  .coef_in(coef[127]), .rdup_out(a1_wr[127]), .rdlo_out(a1_wr[639]));
			radix2 #(.width(width)) rd_st0_128  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[128]), .rdlo_in(a0_wr[640]),  .coef_in(coef[128]), .rdup_out(a1_wr[128]), .rdlo_out(a1_wr[640]));
			radix2 #(.width(width)) rd_st0_129  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[129]), .rdlo_in(a0_wr[641]),  .coef_in(coef[129]), .rdup_out(a1_wr[129]), .rdlo_out(a1_wr[641]));
			radix2 #(.width(width)) rd_st0_130  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[130]), .rdlo_in(a0_wr[642]),  .coef_in(coef[130]), .rdup_out(a1_wr[130]), .rdlo_out(a1_wr[642]));
			radix2 #(.width(width)) rd_st0_131  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[131]), .rdlo_in(a0_wr[643]),  .coef_in(coef[131]), .rdup_out(a1_wr[131]), .rdlo_out(a1_wr[643]));
			radix2 #(.width(width)) rd_st0_132  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[132]), .rdlo_in(a0_wr[644]),  .coef_in(coef[132]), .rdup_out(a1_wr[132]), .rdlo_out(a1_wr[644]));
			radix2 #(.width(width)) rd_st0_133  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[133]), .rdlo_in(a0_wr[645]),  .coef_in(coef[133]), .rdup_out(a1_wr[133]), .rdlo_out(a1_wr[645]));
			radix2 #(.width(width)) rd_st0_134  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[134]), .rdlo_in(a0_wr[646]),  .coef_in(coef[134]), .rdup_out(a1_wr[134]), .rdlo_out(a1_wr[646]));
			radix2 #(.width(width)) rd_st0_135  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[135]), .rdlo_in(a0_wr[647]),  .coef_in(coef[135]), .rdup_out(a1_wr[135]), .rdlo_out(a1_wr[647]));
			radix2 #(.width(width)) rd_st0_136  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[136]), .rdlo_in(a0_wr[648]),  .coef_in(coef[136]), .rdup_out(a1_wr[136]), .rdlo_out(a1_wr[648]));
			radix2 #(.width(width)) rd_st0_137  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[137]), .rdlo_in(a0_wr[649]),  .coef_in(coef[137]), .rdup_out(a1_wr[137]), .rdlo_out(a1_wr[649]));
			radix2 #(.width(width)) rd_st0_138  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[138]), .rdlo_in(a0_wr[650]),  .coef_in(coef[138]), .rdup_out(a1_wr[138]), .rdlo_out(a1_wr[650]));
			radix2 #(.width(width)) rd_st0_139  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[139]), .rdlo_in(a0_wr[651]),  .coef_in(coef[139]), .rdup_out(a1_wr[139]), .rdlo_out(a1_wr[651]));
			radix2 #(.width(width)) rd_st0_140  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[140]), .rdlo_in(a0_wr[652]),  .coef_in(coef[140]), .rdup_out(a1_wr[140]), .rdlo_out(a1_wr[652]));
			radix2 #(.width(width)) rd_st0_141  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[141]), .rdlo_in(a0_wr[653]),  .coef_in(coef[141]), .rdup_out(a1_wr[141]), .rdlo_out(a1_wr[653]));
			radix2 #(.width(width)) rd_st0_142  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[142]), .rdlo_in(a0_wr[654]),  .coef_in(coef[142]), .rdup_out(a1_wr[142]), .rdlo_out(a1_wr[654]));
			radix2 #(.width(width)) rd_st0_143  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[143]), .rdlo_in(a0_wr[655]),  .coef_in(coef[143]), .rdup_out(a1_wr[143]), .rdlo_out(a1_wr[655]));
			radix2 #(.width(width)) rd_st0_144  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[144]), .rdlo_in(a0_wr[656]),  .coef_in(coef[144]), .rdup_out(a1_wr[144]), .rdlo_out(a1_wr[656]));
			radix2 #(.width(width)) rd_st0_145  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[145]), .rdlo_in(a0_wr[657]),  .coef_in(coef[145]), .rdup_out(a1_wr[145]), .rdlo_out(a1_wr[657]));
			radix2 #(.width(width)) rd_st0_146  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[146]), .rdlo_in(a0_wr[658]),  .coef_in(coef[146]), .rdup_out(a1_wr[146]), .rdlo_out(a1_wr[658]));
			radix2 #(.width(width)) rd_st0_147  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[147]), .rdlo_in(a0_wr[659]),  .coef_in(coef[147]), .rdup_out(a1_wr[147]), .rdlo_out(a1_wr[659]));
			radix2 #(.width(width)) rd_st0_148  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[148]), .rdlo_in(a0_wr[660]),  .coef_in(coef[148]), .rdup_out(a1_wr[148]), .rdlo_out(a1_wr[660]));
			radix2 #(.width(width)) rd_st0_149  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[149]), .rdlo_in(a0_wr[661]),  .coef_in(coef[149]), .rdup_out(a1_wr[149]), .rdlo_out(a1_wr[661]));
			radix2 #(.width(width)) rd_st0_150  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[150]), .rdlo_in(a0_wr[662]),  .coef_in(coef[150]), .rdup_out(a1_wr[150]), .rdlo_out(a1_wr[662]));
			radix2 #(.width(width)) rd_st0_151  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[151]), .rdlo_in(a0_wr[663]),  .coef_in(coef[151]), .rdup_out(a1_wr[151]), .rdlo_out(a1_wr[663]));
			radix2 #(.width(width)) rd_st0_152  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[152]), .rdlo_in(a0_wr[664]),  .coef_in(coef[152]), .rdup_out(a1_wr[152]), .rdlo_out(a1_wr[664]));
			radix2 #(.width(width)) rd_st0_153  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[153]), .rdlo_in(a0_wr[665]),  .coef_in(coef[153]), .rdup_out(a1_wr[153]), .rdlo_out(a1_wr[665]));
			radix2 #(.width(width)) rd_st0_154  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[154]), .rdlo_in(a0_wr[666]),  .coef_in(coef[154]), .rdup_out(a1_wr[154]), .rdlo_out(a1_wr[666]));
			radix2 #(.width(width)) rd_st0_155  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[155]), .rdlo_in(a0_wr[667]),  .coef_in(coef[155]), .rdup_out(a1_wr[155]), .rdlo_out(a1_wr[667]));
			radix2 #(.width(width)) rd_st0_156  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[156]), .rdlo_in(a0_wr[668]),  .coef_in(coef[156]), .rdup_out(a1_wr[156]), .rdlo_out(a1_wr[668]));
			radix2 #(.width(width)) rd_st0_157  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[157]), .rdlo_in(a0_wr[669]),  .coef_in(coef[157]), .rdup_out(a1_wr[157]), .rdlo_out(a1_wr[669]));
			radix2 #(.width(width)) rd_st0_158  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[158]), .rdlo_in(a0_wr[670]),  .coef_in(coef[158]), .rdup_out(a1_wr[158]), .rdlo_out(a1_wr[670]));
			radix2 #(.width(width)) rd_st0_159  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[159]), .rdlo_in(a0_wr[671]),  .coef_in(coef[159]), .rdup_out(a1_wr[159]), .rdlo_out(a1_wr[671]));
			radix2 #(.width(width)) rd_st0_160  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[160]), .rdlo_in(a0_wr[672]),  .coef_in(coef[160]), .rdup_out(a1_wr[160]), .rdlo_out(a1_wr[672]));
			radix2 #(.width(width)) rd_st0_161  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[161]), .rdlo_in(a0_wr[673]),  .coef_in(coef[161]), .rdup_out(a1_wr[161]), .rdlo_out(a1_wr[673]));
			radix2 #(.width(width)) rd_st0_162  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[162]), .rdlo_in(a0_wr[674]),  .coef_in(coef[162]), .rdup_out(a1_wr[162]), .rdlo_out(a1_wr[674]));
			radix2 #(.width(width)) rd_st0_163  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[163]), .rdlo_in(a0_wr[675]),  .coef_in(coef[163]), .rdup_out(a1_wr[163]), .rdlo_out(a1_wr[675]));
			radix2 #(.width(width)) rd_st0_164  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[164]), .rdlo_in(a0_wr[676]),  .coef_in(coef[164]), .rdup_out(a1_wr[164]), .rdlo_out(a1_wr[676]));
			radix2 #(.width(width)) rd_st0_165  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[165]), .rdlo_in(a0_wr[677]),  .coef_in(coef[165]), .rdup_out(a1_wr[165]), .rdlo_out(a1_wr[677]));
			radix2 #(.width(width)) rd_st0_166  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[166]), .rdlo_in(a0_wr[678]),  .coef_in(coef[166]), .rdup_out(a1_wr[166]), .rdlo_out(a1_wr[678]));
			radix2 #(.width(width)) rd_st0_167  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[167]), .rdlo_in(a0_wr[679]),  .coef_in(coef[167]), .rdup_out(a1_wr[167]), .rdlo_out(a1_wr[679]));
			radix2 #(.width(width)) rd_st0_168  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[168]), .rdlo_in(a0_wr[680]),  .coef_in(coef[168]), .rdup_out(a1_wr[168]), .rdlo_out(a1_wr[680]));
			radix2 #(.width(width)) rd_st0_169  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[169]), .rdlo_in(a0_wr[681]),  .coef_in(coef[169]), .rdup_out(a1_wr[169]), .rdlo_out(a1_wr[681]));
			radix2 #(.width(width)) rd_st0_170  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[170]), .rdlo_in(a0_wr[682]),  .coef_in(coef[170]), .rdup_out(a1_wr[170]), .rdlo_out(a1_wr[682]));
			radix2 #(.width(width)) rd_st0_171  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[171]), .rdlo_in(a0_wr[683]),  .coef_in(coef[171]), .rdup_out(a1_wr[171]), .rdlo_out(a1_wr[683]));
			radix2 #(.width(width)) rd_st0_172  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[172]), .rdlo_in(a0_wr[684]),  .coef_in(coef[172]), .rdup_out(a1_wr[172]), .rdlo_out(a1_wr[684]));
			radix2 #(.width(width)) rd_st0_173  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[173]), .rdlo_in(a0_wr[685]),  .coef_in(coef[173]), .rdup_out(a1_wr[173]), .rdlo_out(a1_wr[685]));
			radix2 #(.width(width)) rd_st0_174  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[174]), .rdlo_in(a0_wr[686]),  .coef_in(coef[174]), .rdup_out(a1_wr[174]), .rdlo_out(a1_wr[686]));
			radix2 #(.width(width)) rd_st0_175  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[175]), .rdlo_in(a0_wr[687]),  .coef_in(coef[175]), .rdup_out(a1_wr[175]), .rdlo_out(a1_wr[687]));
			radix2 #(.width(width)) rd_st0_176  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[176]), .rdlo_in(a0_wr[688]),  .coef_in(coef[176]), .rdup_out(a1_wr[176]), .rdlo_out(a1_wr[688]));
			radix2 #(.width(width)) rd_st0_177  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[177]), .rdlo_in(a0_wr[689]),  .coef_in(coef[177]), .rdup_out(a1_wr[177]), .rdlo_out(a1_wr[689]));
			radix2 #(.width(width)) rd_st0_178  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[178]), .rdlo_in(a0_wr[690]),  .coef_in(coef[178]), .rdup_out(a1_wr[178]), .rdlo_out(a1_wr[690]));
			radix2 #(.width(width)) rd_st0_179  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[179]), .rdlo_in(a0_wr[691]),  .coef_in(coef[179]), .rdup_out(a1_wr[179]), .rdlo_out(a1_wr[691]));
			radix2 #(.width(width)) rd_st0_180  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[180]), .rdlo_in(a0_wr[692]),  .coef_in(coef[180]), .rdup_out(a1_wr[180]), .rdlo_out(a1_wr[692]));
			radix2 #(.width(width)) rd_st0_181  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[181]), .rdlo_in(a0_wr[693]),  .coef_in(coef[181]), .rdup_out(a1_wr[181]), .rdlo_out(a1_wr[693]));
			radix2 #(.width(width)) rd_st0_182  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[182]), .rdlo_in(a0_wr[694]),  .coef_in(coef[182]), .rdup_out(a1_wr[182]), .rdlo_out(a1_wr[694]));
			radix2 #(.width(width)) rd_st0_183  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[183]), .rdlo_in(a0_wr[695]),  .coef_in(coef[183]), .rdup_out(a1_wr[183]), .rdlo_out(a1_wr[695]));
			radix2 #(.width(width)) rd_st0_184  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[184]), .rdlo_in(a0_wr[696]),  .coef_in(coef[184]), .rdup_out(a1_wr[184]), .rdlo_out(a1_wr[696]));
			radix2 #(.width(width)) rd_st0_185  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[185]), .rdlo_in(a0_wr[697]),  .coef_in(coef[185]), .rdup_out(a1_wr[185]), .rdlo_out(a1_wr[697]));
			radix2 #(.width(width)) rd_st0_186  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[186]), .rdlo_in(a0_wr[698]),  .coef_in(coef[186]), .rdup_out(a1_wr[186]), .rdlo_out(a1_wr[698]));
			radix2 #(.width(width)) rd_st0_187  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[187]), .rdlo_in(a0_wr[699]),  .coef_in(coef[187]), .rdup_out(a1_wr[187]), .rdlo_out(a1_wr[699]));
			radix2 #(.width(width)) rd_st0_188  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[188]), .rdlo_in(a0_wr[700]),  .coef_in(coef[188]), .rdup_out(a1_wr[188]), .rdlo_out(a1_wr[700]));
			radix2 #(.width(width)) rd_st0_189  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[189]), .rdlo_in(a0_wr[701]),  .coef_in(coef[189]), .rdup_out(a1_wr[189]), .rdlo_out(a1_wr[701]));
			radix2 #(.width(width)) rd_st0_190  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[190]), .rdlo_in(a0_wr[702]),  .coef_in(coef[190]), .rdup_out(a1_wr[190]), .rdlo_out(a1_wr[702]));
			radix2 #(.width(width)) rd_st0_191  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[191]), .rdlo_in(a0_wr[703]),  .coef_in(coef[191]), .rdup_out(a1_wr[191]), .rdlo_out(a1_wr[703]));
			radix2 #(.width(width)) rd_st0_192  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[192]), .rdlo_in(a0_wr[704]),  .coef_in(coef[192]), .rdup_out(a1_wr[192]), .rdlo_out(a1_wr[704]));
			radix2 #(.width(width)) rd_st0_193  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[193]), .rdlo_in(a0_wr[705]),  .coef_in(coef[193]), .rdup_out(a1_wr[193]), .rdlo_out(a1_wr[705]));
			radix2 #(.width(width)) rd_st0_194  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[194]), .rdlo_in(a0_wr[706]),  .coef_in(coef[194]), .rdup_out(a1_wr[194]), .rdlo_out(a1_wr[706]));
			radix2 #(.width(width)) rd_st0_195  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[195]), .rdlo_in(a0_wr[707]),  .coef_in(coef[195]), .rdup_out(a1_wr[195]), .rdlo_out(a1_wr[707]));
			radix2 #(.width(width)) rd_st0_196  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[196]), .rdlo_in(a0_wr[708]),  .coef_in(coef[196]), .rdup_out(a1_wr[196]), .rdlo_out(a1_wr[708]));
			radix2 #(.width(width)) rd_st0_197  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[197]), .rdlo_in(a0_wr[709]),  .coef_in(coef[197]), .rdup_out(a1_wr[197]), .rdlo_out(a1_wr[709]));
			radix2 #(.width(width)) rd_st0_198  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[198]), .rdlo_in(a0_wr[710]),  .coef_in(coef[198]), .rdup_out(a1_wr[198]), .rdlo_out(a1_wr[710]));
			radix2 #(.width(width)) rd_st0_199  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[199]), .rdlo_in(a0_wr[711]),  .coef_in(coef[199]), .rdup_out(a1_wr[199]), .rdlo_out(a1_wr[711]));
			radix2 #(.width(width)) rd_st0_200  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[200]), .rdlo_in(a0_wr[712]),  .coef_in(coef[200]), .rdup_out(a1_wr[200]), .rdlo_out(a1_wr[712]));
			radix2 #(.width(width)) rd_st0_201  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[201]), .rdlo_in(a0_wr[713]),  .coef_in(coef[201]), .rdup_out(a1_wr[201]), .rdlo_out(a1_wr[713]));
			radix2 #(.width(width)) rd_st0_202  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[202]), .rdlo_in(a0_wr[714]),  .coef_in(coef[202]), .rdup_out(a1_wr[202]), .rdlo_out(a1_wr[714]));
			radix2 #(.width(width)) rd_st0_203  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[203]), .rdlo_in(a0_wr[715]),  .coef_in(coef[203]), .rdup_out(a1_wr[203]), .rdlo_out(a1_wr[715]));
			radix2 #(.width(width)) rd_st0_204  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[204]), .rdlo_in(a0_wr[716]),  .coef_in(coef[204]), .rdup_out(a1_wr[204]), .rdlo_out(a1_wr[716]));
			radix2 #(.width(width)) rd_st0_205  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[205]), .rdlo_in(a0_wr[717]),  .coef_in(coef[205]), .rdup_out(a1_wr[205]), .rdlo_out(a1_wr[717]));
			radix2 #(.width(width)) rd_st0_206  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[206]), .rdlo_in(a0_wr[718]),  .coef_in(coef[206]), .rdup_out(a1_wr[206]), .rdlo_out(a1_wr[718]));
			radix2 #(.width(width)) rd_st0_207  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[207]), .rdlo_in(a0_wr[719]),  .coef_in(coef[207]), .rdup_out(a1_wr[207]), .rdlo_out(a1_wr[719]));
			radix2 #(.width(width)) rd_st0_208  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[208]), .rdlo_in(a0_wr[720]),  .coef_in(coef[208]), .rdup_out(a1_wr[208]), .rdlo_out(a1_wr[720]));
			radix2 #(.width(width)) rd_st0_209  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[209]), .rdlo_in(a0_wr[721]),  .coef_in(coef[209]), .rdup_out(a1_wr[209]), .rdlo_out(a1_wr[721]));
			radix2 #(.width(width)) rd_st0_210  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[210]), .rdlo_in(a0_wr[722]),  .coef_in(coef[210]), .rdup_out(a1_wr[210]), .rdlo_out(a1_wr[722]));
			radix2 #(.width(width)) rd_st0_211  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[211]), .rdlo_in(a0_wr[723]),  .coef_in(coef[211]), .rdup_out(a1_wr[211]), .rdlo_out(a1_wr[723]));
			radix2 #(.width(width)) rd_st0_212  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[212]), .rdlo_in(a0_wr[724]),  .coef_in(coef[212]), .rdup_out(a1_wr[212]), .rdlo_out(a1_wr[724]));
			radix2 #(.width(width)) rd_st0_213  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[213]), .rdlo_in(a0_wr[725]),  .coef_in(coef[213]), .rdup_out(a1_wr[213]), .rdlo_out(a1_wr[725]));
			radix2 #(.width(width)) rd_st0_214  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[214]), .rdlo_in(a0_wr[726]),  .coef_in(coef[214]), .rdup_out(a1_wr[214]), .rdlo_out(a1_wr[726]));
			radix2 #(.width(width)) rd_st0_215  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[215]), .rdlo_in(a0_wr[727]),  .coef_in(coef[215]), .rdup_out(a1_wr[215]), .rdlo_out(a1_wr[727]));
			radix2 #(.width(width)) rd_st0_216  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[216]), .rdlo_in(a0_wr[728]),  .coef_in(coef[216]), .rdup_out(a1_wr[216]), .rdlo_out(a1_wr[728]));
			radix2 #(.width(width)) rd_st0_217  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[217]), .rdlo_in(a0_wr[729]),  .coef_in(coef[217]), .rdup_out(a1_wr[217]), .rdlo_out(a1_wr[729]));
			radix2 #(.width(width)) rd_st0_218  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[218]), .rdlo_in(a0_wr[730]),  .coef_in(coef[218]), .rdup_out(a1_wr[218]), .rdlo_out(a1_wr[730]));
			radix2 #(.width(width)) rd_st0_219  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[219]), .rdlo_in(a0_wr[731]),  .coef_in(coef[219]), .rdup_out(a1_wr[219]), .rdlo_out(a1_wr[731]));
			radix2 #(.width(width)) rd_st0_220  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[220]), .rdlo_in(a0_wr[732]),  .coef_in(coef[220]), .rdup_out(a1_wr[220]), .rdlo_out(a1_wr[732]));
			radix2 #(.width(width)) rd_st0_221  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[221]), .rdlo_in(a0_wr[733]),  .coef_in(coef[221]), .rdup_out(a1_wr[221]), .rdlo_out(a1_wr[733]));
			radix2 #(.width(width)) rd_st0_222  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[222]), .rdlo_in(a0_wr[734]),  .coef_in(coef[222]), .rdup_out(a1_wr[222]), .rdlo_out(a1_wr[734]));
			radix2 #(.width(width)) rd_st0_223  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[223]), .rdlo_in(a0_wr[735]),  .coef_in(coef[223]), .rdup_out(a1_wr[223]), .rdlo_out(a1_wr[735]));
			radix2 #(.width(width)) rd_st0_224  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[224]), .rdlo_in(a0_wr[736]),  .coef_in(coef[224]), .rdup_out(a1_wr[224]), .rdlo_out(a1_wr[736]));
			radix2 #(.width(width)) rd_st0_225  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[225]), .rdlo_in(a0_wr[737]),  .coef_in(coef[225]), .rdup_out(a1_wr[225]), .rdlo_out(a1_wr[737]));
			radix2 #(.width(width)) rd_st0_226  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[226]), .rdlo_in(a0_wr[738]),  .coef_in(coef[226]), .rdup_out(a1_wr[226]), .rdlo_out(a1_wr[738]));
			radix2 #(.width(width)) rd_st0_227  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[227]), .rdlo_in(a0_wr[739]),  .coef_in(coef[227]), .rdup_out(a1_wr[227]), .rdlo_out(a1_wr[739]));
			radix2 #(.width(width)) rd_st0_228  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[228]), .rdlo_in(a0_wr[740]),  .coef_in(coef[228]), .rdup_out(a1_wr[228]), .rdlo_out(a1_wr[740]));
			radix2 #(.width(width)) rd_st0_229  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[229]), .rdlo_in(a0_wr[741]),  .coef_in(coef[229]), .rdup_out(a1_wr[229]), .rdlo_out(a1_wr[741]));
			radix2 #(.width(width)) rd_st0_230  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[230]), .rdlo_in(a0_wr[742]),  .coef_in(coef[230]), .rdup_out(a1_wr[230]), .rdlo_out(a1_wr[742]));
			radix2 #(.width(width)) rd_st0_231  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[231]), .rdlo_in(a0_wr[743]),  .coef_in(coef[231]), .rdup_out(a1_wr[231]), .rdlo_out(a1_wr[743]));
			radix2 #(.width(width)) rd_st0_232  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[232]), .rdlo_in(a0_wr[744]),  .coef_in(coef[232]), .rdup_out(a1_wr[232]), .rdlo_out(a1_wr[744]));
			radix2 #(.width(width)) rd_st0_233  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[233]), .rdlo_in(a0_wr[745]),  .coef_in(coef[233]), .rdup_out(a1_wr[233]), .rdlo_out(a1_wr[745]));
			radix2 #(.width(width)) rd_st0_234  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[234]), .rdlo_in(a0_wr[746]),  .coef_in(coef[234]), .rdup_out(a1_wr[234]), .rdlo_out(a1_wr[746]));
			radix2 #(.width(width)) rd_st0_235  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[235]), .rdlo_in(a0_wr[747]),  .coef_in(coef[235]), .rdup_out(a1_wr[235]), .rdlo_out(a1_wr[747]));
			radix2 #(.width(width)) rd_st0_236  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[236]), .rdlo_in(a0_wr[748]),  .coef_in(coef[236]), .rdup_out(a1_wr[236]), .rdlo_out(a1_wr[748]));
			radix2 #(.width(width)) rd_st0_237  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[237]), .rdlo_in(a0_wr[749]),  .coef_in(coef[237]), .rdup_out(a1_wr[237]), .rdlo_out(a1_wr[749]));
			radix2 #(.width(width)) rd_st0_238  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[238]), .rdlo_in(a0_wr[750]),  .coef_in(coef[238]), .rdup_out(a1_wr[238]), .rdlo_out(a1_wr[750]));
			radix2 #(.width(width)) rd_st0_239  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[239]), .rdlo_in(a0_wr[751]),  .coef_in(coef[239]), .rdup_out(a1_wr[239]), .rdlo_out(a1_wr[751]));
			radix2 #(.width(width)) rd_st0_240  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[240]), .rdlo_in(a0_wr[752]),  .coef_in(coef[240]), .rdup_out(a1_wr[240]), .rdlo_out(a1_wr[752]));
			radix2 #(.width(width)) rd_st0_241  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[241]), .rdlo_in(a0_wr[753]),  .coef_in(coef[241]), .rdup_out(a1_wr[241]), .rdlo_out(a1_wr[753]));
			radix2 #(.width(width)) rd_st0_242  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[242]), .rdlo_in(a0_wr[754]),  .coef_in(coef[242]), .rdup_out(a1_wr[242]), .rdlo_out(a1_wr[754]));
			radix2 #(.width(width)) rd_st0_243  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[243]), .rdlo_in(a0_wr[755]),  .coef_in(coef[243]), .rdup_out(a1_wr[243]), .rdlo_out(a1_wr[755]));
			radix2 #(.width(width)) rd_st0_244  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[244]), .rdlo_in(a0_wr[756]),  .coef_in(coef[244]), .rdup_out(a1_wr[244]), .rdlo_out(a1_wr[756]));
			radix2 #(.width(width)) rd_st0_245  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[245]), .rdlo_in(a0_wr[757]),  .coef_in(coef[245]), .rdup_out(a1_wr[245]), .rdlo_out(a1_wr[757]));
			radix2 #(.width(width)) rd_st0_246  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[246]), .rdlo_in(a0_wr[758]),  .coef_in(coef[246]), .rdup_out(a1_wr[246]), .rdlo_out(a1_wr[758]));
			radix2 #(.width(width)) rd_st0_247  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[247]), .rdlo_in(a0_wr[759]),  .coef_in(coef[247]), .rdup_out(a1_wr[247]), .rdlo_out(a1_wr[759]));
			radix2 #(.width(width)) rd_st0_248  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[248]), .rdlo_in(a0_wr[760]),  .coef_in(coef[248]), .rdup_out(a1_wr[248]), .rdlo_out(a1_wr[760]));
			radix2 #(.width(width)) rd_st0_249  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[249]), .rdlo_in(a0_wr[761]),  .coef_in(coef[249]), .rdup_out(a1_wr[249]), .rdlo_out(a1_wr[761]));
			radix2 #(.width(width)) rd_st0_250  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[250]), .rdlo_in(a0_wr[762]),  .coef_in(coef[250]), .rdup_out(a1_wr[250]), .rdlo_out(a1_wr[762]));
			radix2 #(.width(width)) rd_st0_251  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[251]), .rdlo_in(a0_wr[763]),  .coef_in(coef[251]), .rdup_out(a1_wr[251]), .rdlo_out(a1_wr[763]));
			radix2 #(.width(width)) rd_st0_252  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[252]), .rdlo_in(a0_wr[764]),  .coef_in(coef[252]), .rdup_out(a1_wr[252]), .rdlo_out(a1_wr[764]));
			radix2 #(.width(width)) rd_st0_253  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[253]), .rdlo_in(a0_wr[765]),  .coef_in(coef[253]), .rdup_out(a1_wr[253]), .rdlo_out(a1_wr[765]));
			radix2 #(.width(width)) rd_st0_254  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[254]), .rdlo_in(a0_wr[766]),  .coef_in(coef[254]), .rdup_out(a1_wr[254]), .rdlo_out(a1_wr[766]));
			radix2 #(.width(width)) rd_st0_255  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[255]), .rdlo_in(a0_wr[767]),  .coef_in(coef[255]), .rdup_out(a1_wr[255]), .rdlo_out(a1_wr[767]));
			radix2 #(.width(width)) rd_st0_256  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[256]), .rdlo_in(a0_wr[768]),  .coef_in(coef[256]), .rdup_out(a1_wr[256]), .rdlo_out(a1_wr[768]));
			radix2 #(.width(width)) rd_st0_257  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[257]), .rdlo_in(a0_wr[769]),  .coef_in(coef[257]), .rdup_out(a1_wr[257]), .rdlo_out(a1_wr[769]));
			radix2 #(.width(width)) rd_st0_258  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[258]), .rdlo_in(a0_wr[770]),  .coef_in(coef[258]), .rdup_out(a1_wr[258]), .rdlo_out(a1_wr[770]));
			radix2 #(.width(width)) rd_st0_259  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[259]), .rdlo_in(a0_wr[771]),  .coef_in(coef[259]), .rdup_out(a1_wr[259]), .rdlo_out(a1_wr[771]));
			radix2 #(.width(width)) rd_st0_260  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[260]), .rdlo_in(a0_wr[772]),  .coef_in(coef[260]), .rdup_out(a1_wr[260]), .rdlo_out(a1_wr[772]));
			radix2 #(.width(width)) rd_st0_261  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[261]), .rdlo_in(a0_wr[773]),  .coef_in(coef[261]), .rdup_out(a1_wr[261]), .rdlo_out(a1_wr[773]));
			radix2 #(.width(width)) rd_st0_262  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[262]), .rdlo_in(a0_wr[774]),  .coef_in(coef[262]), .rdup_out(a1_wr[262]), .rdlo_out(a1_wr[774]));
			radix2 #(.width(width)) rd_st0_263  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[263]), .rdlo_in(a0_wr[775]),  .coef_in(coef[263]), .rdup_out(a1_wr[263]), .rdlo_out(a1_wr[775]));
			radix2 #(.width(width)) rd_st0_264  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[264]), .rdlo_in(a0_wr[776]),  .coef_in(coef[264]), .rdup_out(a1_wr[264]), .rdlo_out(a1_wr[776]));
			radix2 #(.width(width)) rd_st0_265  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[265]), .rdlo_in(a0_wr[777]),  .coef_in(coef[265]), .rdup_out(a1_wr[265]), .rdlo_out(a1_wr[777]));
			radix2 #(.width(width)) rd_st0_266  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[266]), .rdlo_in(a0_wr[778]),  .coef_in(coef[266]), .rdup_out(a1_wr[266]), .rdlo_out(a1_wr[778]));
			radix2 #(.width(width)) rd_st0_267  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[267]), .rdlo_in(a0_wr[779]),  .coef_in(coef[267]), .rdup_out(a1_wr[267]), .rdlo_out(a1_wr[779]));
			radix2 #(.width(width)) rd_st0_268  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[268]), .rdlo_in(a0_wr[780]),  .coef_in(coef[268]), .rdup_out(a1_wr[268]), .rdlo_out(a1_wr[780]));
			radix2 #(.width(width)) rd_st0_269  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[269]), .rdlo_in(a0_wr[781]),  .coef_in(coef[269]), .rdup_out(a1_wr[269]), .rdlo_out(a1_wr[781]));
			radix2 #(.width(width)) rd_st0_270  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[270]), .rdlo_in(a0_wr[782]),  .coef_in(coef[270]), .rdup_out(a1_wr[270]), .rdlo_out(a1_wr[782]));
			radix2 #(.width(width)) rd_st0_271  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[271]), .rdlo_in(a0_wr[783]),  .coef_in(coef[271]), .rdup_out(a1_wr[271]), .rdlo_out(a1_wr[783]));
			radix2 #(.width(width)) rd_st0_272  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[272]), .rdlo_in(a0_wr[784]),  .coef_in(coef[272]), .rdup_out(a1_wr[272]), .rdlo_out(a1_wr[784]));
			radix2 #(.width(width)) rd_st0_273  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[273]), .rdlo_in(a0_wr[785]),  .coef_in(coef[273]), .rdup_out(a1_wr[273]), .rdlo_out(a1_wr[785]));
			radix2 #(.width(width)) rd_st0_274  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[274]), .rdlo_in(a0_wr[786]),  .coef_in(coef[274]), .rdup_out(a1_wr[274]), .rdlo_out(a1_wr[786]));
			radix2 #(.width(width)) rd_st0_275  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[275]), .rdlo_in(a0_wr[787]),  .coef_in(coef[275]), .rdup_out(a1_wr[275]), .rdlo_out(a1_wr[787]));
			radix2 #(.width(width)) rd_st0_276  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[276]), .rdlo_in(a0_wr[788]),  .coef_in(coef[276]), .rdup_out(a1_wr[276]), .rdlo_out(a1_wr[788]));
			radix2 #(.width(width)) rd_st0_277  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[277]), .rdlo_in(a0_wr[789]),  .coef_in(coef[277]), .rdup_out(a1_wr[277]), .rdlo_out(a1_wr[789]));
			radix2 #(.width(width)) rd_st0_278  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[278]), .rdlo_in(a0_wr[790]),  .coef_in(coef[278]), .rdup_out(a1_wr[278]), .rdlo_out(a1_wr[790]));
			radix2 #(.width(width)) rd_st0_279  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[279]), .rdlo_in(a0_wr[791]),  .coef_in(coef[279]), .rdup_out(a1_wr[279]), .rdlo_out(a1_wr[791]));
			radix2 #(.width(width)) rd_st0_280  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[280]), .rdlo_in(a0_wr[792]),  .coef_in(coef[280]), .rdup_out(a1_wr[280]), .rdlo_out(a1_wr[792]));
			radix2 #(.width(width)) rd_st0_281  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[281]), .rdlo_in(a0_wr[793]),  .coef_in(coef[281]), .rdup_out(a1_wr[281]), .rdlo_out(a1_wr[793]));
			radix2 #(.width(width)) rd_st0_282  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[282]), .rdlo_in(a0_wr[794]),  .coef_in(coef[282]), .rdup_out(a1_wr[282]), .rdlo_out(a1_wr[794]));
			radix2 #(.width(width)) rd_st0_283  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[283]), .rdlo_in(a0_wr[795]),  .coef_in(coef[283]), .rdup_out(a1_wr[283]), .rdlo_out(a1_wr[795]));
			radix2 #(.width(width)) rd_st0_284  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[284]), .rdlo_in(a0_wr[796]),  .coef_in(coef[284]), .rdup_out(a1_wr[284]), .rdlo_out(a1_wr[796]));
			radix2 #(.width(width)) rd_st0_285  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[285]), .rdlo_in(a0_wr[797]),  .coef_in(coef[285]), .rdup_out(a1_wr[285]), .rdlo_out(a1_wr[797]));
			radix2 #(.width(width)) rd_st0_286  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[286]), .rdlo_in(a0_wr[798]),  .coef_in(coef[286]), .rdup_out(a1_wr[286]), .rdlo_out(a1_wr[798]));
			radix2 #(.width(width)) rd_st0_287  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[287]), .rdlo_in(a0_wr[799]),  .coef_in(coef[287]), .rdup_out(a1_wr[287]), .rdlo_out(a1_wr[799]));
			radix2 #(.width(width)) rd_st0_288  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[288]), .rdlo_in(a0_wr[800]),  .coef_in(coef[288]), .rdup_out(a1_wr[288]), .rdlo_out(a1_wr[800]));
			radix2 #(.width(width)) rd_st0_289  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[289]), .rdlo_in(a0_wr[801]),  .coef_in(coef[289]), .rdup_out(a1_wr[289]), .rdlo_out(a1_wr[801]));
			radix2 #(.width(width)) rd_st0_290  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[290]), .rdlo_in(a0_wr[802]),  .coef_in(coef[290]), .rdup_out(a1_wr[290]), .rdlo_out(a1_wr[802]));
			radix2 #(.width(width)) rd_st0_291  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[291]), .rdlo_in(a0_wr[803]),  .coef_in(coef[291]), .rdup_out(a1_wr[291]), .rdlo_out(a1_wr[803]));
			radix2 #(.width(width)) rd_st0_292  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[292]), .rdlo_in(a0_wr[804]),  .coef_in(coef[292]), .rdup_out(a1_wr[292]), .rdlo_out(a1_wr[804]));
			radix2 #(.width(width)) rd_st0_293  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[293]), .rdlo_in(a0_wr[805]),  .coef_in(coef[293]), .rdup_out(a1_wr[293]), .rdlo_out(a1_wr[805]));
			radix2 #(.width(width)) rd_st0_294  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[294]), .rdlo_in(a0_wr[806]),  .coef_in(coef[294]), .rdup_out(a1_wr[294]), .rdlo_out(a1_wr[806]));
			radix2 #(.width(width)) rd_st0_295  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[295]), .rdlo_in(a0_wr[807]),  .coef_in(coef[295]), .rdup_out(a1_wr[295]), .rdlo_out(a1_wr[807]));
			radix2 #(.width(width)) rd_st0_296  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[296]), .rdlo_in(a0_wr[808]),  .coef_in(coef[296]), .rdup_out(a1_wr[296]), .rdlo_out(a1_wr[808]));
			radix2 #(.width(width)) rd_st0_297  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[297]), .rdlo_in(a0_wr[809]),  .coef_in(coef[297]), .rdup_out(a1_wr[297]), .rdlo_out(a1_wr[809]));
			radix2 #(.width(width)) rd_st0_298  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[298]), .rdlo_in(a0_wr[810]),  .coef_in(coef[298]), .rdup_out(a1_wr[298]), .rdlo_out(a1_wr[810]));
			radix2 #(.width(width)) rd_st0_299  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[299]), .rdlo_in(a0_wr[811]),  .coef_in(coef[299]), .rdup_out(a1_wr[299]), .rdlo_out(a1_wr[811]));
			radix2 #(.width(width)) rd_st0_300  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[300]), .rdlo_in(a0_wr[812]),  .coef_in(coef[300]), .rdup_out(a1_wr[300]), .rdlo_out(a1_wr[812]));
			radix2 #(.width(width)) rd_st0_301  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[301]), .rdlo_in(a0_wr[813]),  .coef_in(coef[301]), .rdup_out(a1_wr[301]), .rdlo_out(a1_wr[813]));
			radix2 #(.width(width)) rd_st0_302  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[302]), .rdlo_in(a0_wr[814]),  .coef_in(coef[302]), .rdup_out(a1_wr[302]), .rdlo_out(a1_wr[814]));
			radix2 #(.width(width)) rd_st0_303  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[303]), .rdlo_in(a0_wr[815]),  .coef_in(coef[303]), .rdup_out(a1_wr[303]), .rdlo_out(a1_wr[815]));
			radix2 #(.width(width)) rd_st0_304  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[304]), .rdlo_in(a0_wr[816]),  .coef_in(coef[304]), .rdup_out(a1_wr[304]), .rdlo_out(a1_wr[816]));
			radix2 #(.width(width)) rd_st0_305  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[305]), .rdlo_in(a0_wr[817]),  .coef_in(coef[305]), .rdup_out(a1_wr[305]), .rdlo_out(a1_wr[817]));
			radix2 #(.width(width)) rd_st0_306  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[306]), .rdlo_in(a0_wr[818]),  .coef_in(coef[306]), .rdup_out(a1_wr[306]), .rdlo_out(a1_wr[818]));
			radix2 #(.width(width)) rd_st0_307  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[307]), .rdlo_in(a0_wr[819]),  .coef_in(coef[307]), .rdup_out(a1_wr[307]), .rdlo_out(a1_wr[819]));
			radix2 #(.width(width)) rd_st0_308  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[308]), .rdlo_in(a0_wr[820]),  .coef_in(coef[308]), .rdup_out(a1_wr[308]), .rdlo_out(a1_wr[820]));
			radix2 #(.width(width)) rd_st0_309  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[309]), .rdlo_in(a0_wr[821]),  .coef_in(coef[309]), .rdup_out(a1_wr[309]), .rdlo_out(a1_wr[821]));
			radix2 #(.width(width)) rd_st0_310  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[310]), .rdlo_in(a0_wr[822]),  .coef_in(coef[310]), .rdup_out(a1_wr[310]), .rdlo_out(a1_wr[822]));
			radix2 #(.width(width)) rd_st0_311  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[311]), .rdlo_in(a0_wr[823]),  .coef_in(coef[311]), .rdup_out(a1_wr[311]), .rdlo_out(a1_wr[823]));
			radix2 #(.width(width)) rd_st0_312  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[312]), .rdlo_in(a0_wr[824]),  .coef_in(coef[312]), .rdup_out(a1_wr[312]), .rdlo_out(a1_wr[824]));
			radix2 #(.width(width)) rd_st0_313  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[313]), .rdlo_in(a0_wr[825]),  .coef_in(coef[313]), .rdup_out(a1_wr[313]), .rdlo_out(a1_wr[825]));
			radix2 #(.width(width)) rd_st0_314  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[314]), .rdlo_in(a0_wr[826]),  .coef_in(coef[314]), .rdup_out(a1_wr[314]), .rdlo_out(a1_wr[826]));
			radix2 #(.width(width)) rd_st0_315  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[315]), .rdlo_in(a0_wr[827]),  .coef_in(coef[315]), .rdup_out(a1_wr[315]), .rdlo_out(a1_wr[827]));
			radix2 #(.width(width)) rd_st0_316  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[316]), .rdlo_in(a0_wr[828]),  .coef_in(coef[316]), .rdup_out(a1_wr[316]), .rdlo_out(a1_wr[828]));
			radix2 #(.width(width)) rd_st0_317  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[317]), .rdlo_in(a0_wr[829]),  .coef_in(coef[317]), .rdup_out(a1_wr[317]), .rdlo_out(a1_wr[829]));
			radix2 #(.width(width)) rd_st0_318  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[318]), .rdlo_in(a0_wr[830]),  .coef_in(coef[318]), .rdup_out(a1_wr[318]), .rdlo_out(a1_wr[830]));
			radix2 #(.width(width)) rd_st0_319  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[319]), .rdlo_in(a0_wr[831]),  .coef_in(coef[319]), .rdup_out(a1_wr[319]), .rdlo_out(a1_wr[831]));
			radix2 #(.width(width)) rd_st0_320  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[320]), .rdlo_in(a0_wr[832]),  .coef_in(coef[320]), .rdup_out(a1_wr[320]), .rdlo_out(a1_wr[832]));
			radix2 #(.width(width)) rd_st0_321  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[321]), .rdlo_in(a0_wr[833]),  .coef_in(coef[321]), .rdup_out(a1_wr[321]), .rdlo_out(a1_wr[833]));
			radix2 #(.width(width)) rd_st0_322  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[322]), .rdlo_in(a0_wr[834]),  .coef_in(coef[322]), .rdup_out(a1_wr[322]), .rdlo_out(a1_wr[834]));
			radix2 #(.width(width)) rd_st0_323  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[323]), .rdlo_in(a0_wr[835]),  .coef_in(coef[323]), .rdup_out(a1_wr[323]), .rdlo_out(a1_wr[835]));
			radix2 #(.width(width)) rd_st0_324  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[324]), .rdlo_in(a0_wr[836]),  .coef_in(coef[324]), .rdup_out(a1_wr[324]), .rdlo_out(a1_wr[836]));
			radix2 #(.width(width)) rd_st0_325  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[325]), .rdlo_in(a0_wr[837]),  .coef_in(coef[325]), .rdup_out(a1_wr[325]), .rdlo_out(a1_wr[837]));
			radix2 #(.width(width)) rd_st0_326  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[326]), .rdlo_in(a0_wr[838]),  .coef_in(coef[326]), .rdup_out(a1_wr[326]), .rdlo_out(a1_wr[838]));
			radix2 #(.width(width)) rd_st0_327  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[327]), .rdlo_in(a0_wr[839]),  .coef_in(coef[327]), .rdup_out(a1_wr[327]), .rdlo_out(a1_wr[839]));
			radix2 #(.width(width)) rd_st0_328  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[328]), .rdlo_in(a0_wr[840]),  .coef_in(coef[328]), .rdup_out(a1_wr[328]), .rdlo_out(a1_wr[840]));
			radix2 #(.width(width)) rd_st0_329  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[329]), .rdlo_in(a0_wr[841]),  .coef_in(coef[329]), .rdup_out(a1_wr[329]), .rdlo_out(a1_wr[841]));
			radix2 #(.width(width)) rd_st0_330  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[330]), .rdlo_in(a0_wr[842]),  .coef_in(coef[330]), .rdup_out(a1_wr[330]), .rdlo_out(a1_wr[842]));
			radix2 #(.width(width)) rd_st0_331  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[331]), .rdlo_in(a0_wr[843]),  .coef_in(coef[331]), .rdup_out(a1_wr[331]), .rdlo_out(a1_wr[843]));
			radix2 #(.width(width)) rd_st0_332  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[332]), .rdlo_in(a0_wr[844]),  .coef_in(coef[332]), .rdup_out(a1_wr[332]), .rdlo_out(a1_wr[844]));
			radix2 #(.width(width)) rd_st0_333  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[333]), .rdlo_in(a0_wr[845]),  .coef_in(coef[333]), .rdup_out(a1_wr[333]), .rdlo_out(a1_wr[845]));
			radix2 #(.width(width)) rd_st0_334  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[334]), .rdlo_in(a0_wr[846]),  .coef_in(coef[334]), .rdup_out(a1_wr[334]), .rdlo_out(a1_wr[846]));
			radix2 #(.width(width)) rd_st0_335  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[335]), .rdlo_in(a0_wr[847]),  .coef_in(coef[335]), .rdup_out(a1_wr[335]), .rdlo_out(a1_wr[847]));
			radix2 #(.width(width)) rd_st0_336  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[336]), .rdlo_in(a0_wr[848]),  .coef_in(coef[336]), .rdup_out(a1_wr[336]), .rdlo_out(a1_wr[848]));
			radix2 #(.width(width)) rd_st0_337  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[337]), .rdlo_in(a0_wr[849]),  .coef_in(coef[337]), .rdup_out(a1_wr[337]), .rdlo_out(a1_wr[849]));
			radix2 #(.width(width)) rd_st0_338  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[338]), .rdlo_in(a0_wr[850]),  .coef_in(coef[338]), .rdup_out(a1_wr[338]), .rdlo_out(a1_wr[850]));
			radix2 #(.width(width)) rd_st0_339  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[339]), .rdlo_in(a0_wr[851]),  .coef_in(coef[339]), .rdup_out(a1_wr[339]), .rdlo_out(a1_wr[851]));
			radix2 #(.width(width)) rd_st0_340  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[340]), .rdlo_in(a0_wr[852]),  .coef_in(coef[340]), .rdup_out(a1_wr[340]), .rdlo_out(a1_wr[852]));
			radix2 #(.width(width)) rd_st0_341  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[341]), .rdlo_in(a0_wr[853]),  .coef_in(coef[341]), .rdup_out(a1_wr[341]), .rdlo_out(a1_wr[853]));
			radix2 #(.width(width)) rd_st0_342  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[342]), .rdlo_in(a0_wr[854]),  .coef_in(coef[342]), .rdup_out(a1_wr[342]), .rdlo_out(a1_wr[854]));
			radix2 #(.width(width)) rd_st0_343  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[343]), .rdlo_in(a0_wr[855]),  .coef_in(coef[343]), .rdup_out(a1_wr[343]), .rdlo_out(a1_wr[855]));
			radix2 #(.width(width)) rd_st0_344  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[344]), .rdlo_in(a0_wr[856]),  .coef_in(coef[344]), .rdup_out(a1_wr[344]), .rdlo_out(a1_wr[856]));
			radix2 #(.width(width)) rd_st0_345  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[345]), .rdlo_in(a0_wr[857]),  .coef_in(coef[345]), .rdup_out(a1_wr[345]), .rdlo_out(a1_wr[857]));
			radix2 #(.width(width)) rd_st0_346  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[346]), .rdlo_in(a0_wr[858]),  .coef_in(coef[346]), .rdup_out(a1_wr[346]), .rdlo_out(a1_wr[858]));
			radix2 #(.width(width)) rd_st0_347  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[347]), .rdlo_in(a0_wr[859]),  .coef_in(coef[347]), .rdup_out(a1_wr[347]), .rdlo_out(a1_wr[859]));
			radix2 #(.width(width)) rd_st0_348  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[348]), .rdlo_in(a0_wr[860]),  .coef_in(coef[348]), .rdup_out(a1_wr[348]), .rdlo_out(a1_wr[860]));
			radix2 #(.width(width)) rd_st0_349  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[349]), .rdlo_in(a0_wr[861]),  .coef_in(coef[349]), .rdup_out(a1_wr[349]), .rdlo_out(a1_wr[861]));
			radix2 #(.width(width)) rd_st0_350  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[350]), .rdlo_in(a0_wr[862]),  .coef_in(coef[350]), .rdup_out(a1_wr[350]), .rdlo_out(a1_wr[862]));
			radix2 #(.width(width)) rd_st0_351  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[351]), .rdlo_in(a0_wr[863]),  .coef_in(coef[351]), .rdup_out(a1_wr[351]), .rdlo_out(a1_wr[863]));
			radix2 #(.width(width)) rd_st0_352  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[352]), .rdlo_in(a0_wr[864]),  .coef_in(coef[352]), .rdup_out(a1_wr[352]), .rdlo_out(a1_wr[864]));
			radix2 #(.width(width)) rd_st0_353  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[353]), .rdlo_in(a0_wr[865]),  .coef_in(coef[353]), .rdup_out(a1_wr[353]), .rdlo_out(a1_wr[865]));
			radix2 #(.width(width)) rd_st0_354  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[354]), .rdlo_in(a0_wr[866]),  .coef_in(coef[354]), .rdup_out(a1_wr[354]), .rdlo_out(a1_wr[866]));
			radix2 #(.width(width)) rd_st0_355  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[355]), .rdlo_in(a0_wr[867]),  .coef_in(coef[355]), .rdup_out(a1_wr[355]), .rdlo_out(a1_wr[867]));
			radix2 #(.width(width)) rd_st0_356  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[356]), .rdlo_in(a0_wr[868]),  .coef_in(coef[356]), .rdup_out(a1_wr[356]), .rdlo_out(a1_wr[868]));
			radix2 #(.width(width)) rd_st0_357  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[357]), .rdlo_in(a0_wr[869]),  .coef_in(coef[357]), .rdup_out(a1_wr[357]), .rdlo_out(a1_wr[869]));
			radix2 #(.width(width)) rd_st0_358  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[358]), .rdlo_in(a0_wr[870]),  .coef_in(coef[358]), .rdup_out(a1_wr[358]), .rdlo_out(a1_wr[870]));
			radix2 #(.width(width)) rd_st0_359  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[359]), .rdlo_in(a0_wr[871]),  .coef_in(coef[359]), .rdup_out(a1_wr[359]), .rdlo_out(a1_wr[871]));
			radix2 #(.width(width)) rd_st0_360  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[360]), .rdlo_in(a0_wr[872]),  .coef_in(coef[360]), .rdup_out(a1_wr[360]), .rdlo_out(a1_wr[872]));
			radix2 #(.width(width)) rd_st0_361  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[361]), .rdlo_in(a0_wr[873]),  .coef_in(coef[361]), .rdup_out(a1_wr[361]), .rdlo_out(a1_wr[873]));
			radix2 #(.width(width)) rd_st0_362  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[362]), .rdlo_in(a0_wr[874]),  .coef_in(coef[362]), .rdup_out(a1_wr[362]), .rdlo_out(a1_wr[874]));
			radix2 #(.width(width)) rd_st0_363  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[363]), .rdlo_in(a0_wr[875]),  .coef_in(coef[363]), .rdup_out(a1_wr[363]), .rdlo_out(a1_wr[875]));
			radix2 #(.width(width)) rd_st0_364  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[364]), .rdlo_in(a0_wr[876]),  .coef_in(coef[364]), .rdup_out(a1_wr[364]), .rdlo_out(a1_wr[876]));
			radix2 #(.width(width)) rd_st0_365  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[365]), .rdlo_in(a0_wr[877]),  .coef_in(coef[365]), .rdup_out(a1_wr[365]), .rdlo_out(a1_wr[877]));
			radix2 #(.width(width)) rd_st0_366  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[366]), .rdlo_in(a0_wr[878]),  .coef_in(coef[366]), .rdup_out(a1_wr[366]), .rdlo_out(a1_wr[878]));
			radix2 #(.width(width)) rd_st0_367  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[367]), .rdlo_in(a0_wr[879]),  .coef_in(coef[367]), .rdup_out(a1_wr[367]), .rdlo_out(a1_wr[879]));
			radix2 #(.width(width)) rd_st0_368  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[368]), .rdlo_in(a0_wr[880]),  .coef_in(coef[368]), .rdup_out(a1_wr[368]), .rdlo_out(a1_wr[880]));
			radix2 #(.width(width)) rd_st0_369  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[369]), .rdlo_in(a0_wr[881]),  .coef_in(coef[369]), .rdup_out(a1_wr[369]), .rdlo_out(a1_wr[881]));
			radix2 #(.width(width)) rd_st0_370  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[370]), .rdlo_in(a0_wr[882]),  .coef_in(coef[370]), .rdup_out(a1_wr[370]), .rdlo_out(a1_wr[882]));
			radix2 #(.width(width)) rd_st0_371  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[371]), .rdlo_in(a0_wr[883]),  .coef_in(coef[371]), .rdup_out(a1_wr[371]), .rdlo_out(a1_wr[883]));
			radix2 #(.width(width)) rd_st0_372  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[372]), .rdlo_in(a0_wr[884]),  .coef_in(coef[372]), .rdup_out(a1_wr[372]), .rdlo_out(a1_wr[884]));
			radix2 #(.width(width)) rd_st0_373  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[373]), .rdlo_in(a0_wr[885]),  .coef_in(coef[373]), .rdup_out(a1_wr[373]), .rdlo_out(a1_wr[885]));
			radix2 #(.width(width)) rd_st0_374  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[374]), .rdlo_in(a0_wr[886]),  .coef_in(coef[374]), .rdup_out(a1_wr[374]), .rdlo_out(a1_wr[886]));
			radix2 #(.width(width)) rd_st0_375  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[375]), .rdlo_in(a0_wr[887]),  .coef_in(coef[375]), .rdup_out(a1_wr[375]), .rdlo_out(a1_wr[887]));
			radix2 #(.width(width)) rd_st0_376  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[376]), .rdlo_in(a0_wr[888]),  .coef_in(coef[376]), .rdup_out(a1_wr[376]), .rdlo_out(a1_wr[888]));
			radix2 #(.width(width)) rd_st0_377  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[377]), .rdlo_in(a0_wr[889]),  .coef_in(coef[377]), .rdup_out(a1_wr[377]), .rdlo_out(a1_wr[889]));
			radix2 #(.width(width)) rd_st0_378  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[378]), .rdlo_in(a0_wr[890]),  .coef_in(coef[378]), .rdup_out(a1_wr[378]), .rdlo_out(a1_wr[890]));
			radix2 #(.width(width)) rd_st0_379  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[379]), .rdlo_in(a0_wr[891]),  .coef_in(coef[379]), .rdup_out(a1_wr[379]), .rdlo_out(a1_wr[891]));
			radix2 #(.width(width)) rd_st0_380  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[380]), .rdlo_in(a0_wr[892]),  .coef_in(coef[380]), .rdup_out(a1_wr[380]), .rdlo_out(a1_wr[892]));
			radix2 #(.width(width)) rd_st0_381  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[381]), .rdlo_in(a0_wr[893]),  .coef_in(coef[381]), .rdup_out(a1_wr[381]), .rdlo_out(a1_wr[893]));
			radix2 #(.width(width)) rd_st0_382  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[382]), .rdlo_in(a0_wr[894]),  .coef_in(coef[382]), .rdup_out(a1_wr[382]), .rdlo_out(a1_wr[894]));
			radix2 #(.width(width)) rd_st0_383  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[383]), .rdlo_in(a0_wr[895]),  .coef_in(coef[383]), .rdup_out(a1_wr[383]), .rdlo_out(a1_wr[895]));
			radix2 #(.width(width)) rd_st0_384  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[384]), .rdlo_in(a0_wr[896]),  .coef_in(coef[384]), .rdup_out(a1_wr[384]), .rdlo_out(a1_wr[896]));
			radix2 #(.width(width)) rd_st0_385  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[385]), .rdlo_in(a0_wr[897]),  .coef_in(coef[385]), .rdup_out(a1_wr[385]), .rdlo_out(a1_wr[897]));
			radix2 #(.width(width)) rd_st0_386  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[386]), .rdlo_in(a0_wr[898]),  .coef_in(coef[386]), .rdup_out(a1_wr[386]), .rdlo_out(a1_wr[898]));
			radix2 #(.width(width)) rd_st0_387  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[387]), .rdlo_in(a0_wr[899]),  .coef_in(coef[387]), .rdup_out(a1_wr[387]), .rdlo_out(a1_wr[899]));
			radix2 #(.width(width)) rd_st0_388  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[388]), .rdlo_in(a0_wr[900]),  .coef_in(coef[388]), .rdup_out(a1_wr[388]), .rdlo_out(a1_wr[900]));
			radix2 #(.width(width)) rd_st0_389  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[389]), .rdlo_in(a0_wr[901]),  .coef_in(coef[389]), .rdup_out(a1_wr[389]), .rdlo_out(a1_wr[901]));
			radix2 #(.width(width)) rd_st0_390  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[390]), .rdlo_in(a0_wr[902]),  .coef_in(coef[390]), .rdup_out(a1_wr[390]), .rdlo_out(a1_wr[902]));
			radix2 #(.width(width)) rd_st0_391  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[391]), .rdlo_in(a0_wr[903]),  .coef_in(coef[391]), .rdup_out(a1_wr[391]), .rdlo_out(a1_wr[903]));
			radix2 #(.width(width)) rd_st0_392  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[392]), .rdlo_in(a0_wr[904]),  .coef_in(coef[392]), .rdup_out(a1_wr[392]), .rdlo_out(a1_wr[904]));
			radix2 #(.width(width)) rd_st0_393  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[393]), .rdlo_in(a0_wr[905]),  .coef_in(coef[393]), .rdup_out(a1_wr[393]), .rdlo_out(a1_wr[905]));
			radix2 #(.width(width)) rd_st0_394  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[394]), .rdlo_in(a0_wr[906]),  .coef_in(coef[394]), .rdup_out(a1_wr[394]), .rdlo_out(a1_wr[906]));
			radix2 #(.width(width)) rd_st0_395  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[395]), .rdlo_in(a0_wr[907]),  .coef_in(coef[395]), .rdup_out(a1_wr[395]), .rdlo_out(a1_wr[907]));
			radix2 #(.width(width)) rd_st0_396  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[396]), .rdlo_in(a0_wr[908]),  .coef_in(coef[396]), .rdup_out(a1_wr[396]), .rdlo_out(a1_wr[908]));
			radix2 #(.width(width)) rd_st0_397  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[397]), .rdlo_in(a0_wr[909]),  .coef_in(coef[397]), .rdup_out(a1_wr[397]), .rdlo_out(a1_wr[909]));
			radix2 #(.width(width)) rd_st0_398  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[398]), .rdlo_in(a0_wr[910]),  .coef_in(coef[398]), .rdup_out(a1_wr[398]), .rdlo_out(a1_wr[910]));
			radix2 #(.width(width)) rd_st0_399  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[399]), .rdlo_in(a0_wr[911]),  .coef_in(coef[399]), .rdup_out(a1_wr[399]), .rdlo_out(a1_wr[911]));
			radix2 #(.width(width)) rd_st0_400  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[400]), .rdlo_in(a0_wr[912]),  .coef_in(coef[400]), .rdup_out(a1_wr[400]), .rdlo_out(a1_wr[912]));
			radix2 #(.width(width)) rd_st0_401  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[401]), .rdlo_in(a0_wr[913]),  .coef_in(coef[401]), .rdup_out(a1_wr[401]), .rdlo_out(a1_wr[913]));
			radix2 #(.width(width)) rd_st0_402  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[402]), .rdlo_in(a0_wr[914]),  .coef_in(coef[402]), .rdup_out(a1_wr[402]), .rdlo_out(a1_wr[914]));
			radix2 #(.width(width)) rd_st0_403  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[403]), .rdlo_in(a0_wr[915]),  .coef_in(coef[403]), .rdup_out(a1_wr[403]), .rdlo_out(a1_wr[915]));
			radix2 #(.width(width)) rd_st0_404  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[404]), .rdlo_in(a0_wr[916]),  .coef_in(coef[404]), .rdup_out(a1_wr[404]), .rdlo_out(a1_wr[916]));
			radix2 #(.width(width)) rd_st0_405  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[405]), .rdlo_in(a0_wr[917]),  .coef_in(coef[405]), .rdup_out(a1_wr[405]), .rdlo_out(a1_wr[917]));
			radix2 #(.width(width)) rd_st0_406  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[406]), .rdlo_in(a0_wr[918]),  .coef_in(coef[406]), .rdup_out(a1_wr[406]), .rdlo_out(a1_wr[918]));
			radix2 #(.width(width)) rd_st0_407  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[407]), .rdlo_in(a0_wr[919]),  .coef_in(coef[407]), .rdup_out(a1_wr[407]), .rdlo_out(a1_wr[919]));
			radix2 #(.width(width)) rd_st0_408  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[408]), .rdlo_in(a0_wr[920]),  .coef_in(coef[408]), .rdup_out(a1_wr[408]), .rdlo_out(a1_wr[920]));
			radix2 #(.width(width)) rd_st0_409  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[409]), .rdlo_in(a0_wr[921]),  .coef_in(coef[409]), .rdup_out(a1_wr[409]), .rdlo_out(a1_wr[921]));
			radix2 #(.width(width)) rd_st0_410  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[410]), .rdlo_in(a0_wr[922]),  .coef_in(coef[410]), .rdup_out(a1_wr[410]), .rdlo_out(a1_wr[922]));
			radix2 #(.width(width)) rd_st0_411  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[411]), .rdlo_in(a0_wr[923]),  .coef_in(coef[411]), .rdup_out(a1_wr[411]), .rdlo_out(a1_wr[923]));
			radix2 #(.width(width)) rd_st0_412  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[412]), .rdlo_in(a0_wr[924]),  .coef_in(coef[412]), .rdup_out(a1_wr[412]), .rdlo_out(a1_wr[924]));
			radix2 #(.width(width)) rd_st0_413  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[413]), .rdlo_in(a0_wr[925]),  .coef_in(coef[413]), .rdup_out(a1_wr[413]), .rdlo_out(a1_wr[925]));
			radix2 #(.width(width)) rd_st0_414  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[414]), .rdlo_in(a0_wr[926]),  .coef_in(coef[414]), .rdup_out(a1_wr[414]), .rdlo_out(a1_wr[926]));
			radix2 #(.width(width)) rd_st0_415  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[415]), .rdlo_in(a0_wr[927]),  .coef_in(coef[415]), .rdup_out(a1_wr[415]), .rdlo_out(a1_wr[927]));
			radix2 #(.width(width)) rd_st0_416  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[416]), .rdlo_in(a0_wr[928]),  .coef_in(coef[416]), .rdup_out(a1_wr[416]), .rdlo_out(a1_wr[928]));
			radix2 #(.width(width)) rd_st0_417  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[417]), .rdlo_in(a0_wr[929]),  .coef_in(coef[417]), .rdup_out(a1_wr[417]), .rdlo_out(a1_wr[929]));
			radix2 #(.width(width)) rd_st0_418  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[418]), .rdlo_in(a0_wr[930]),  .coef_in(coef[418]), .rdup_out(a1_wr[418]), .rdlo_out(a1_wr[930]));
			radix2 #(.width(width)) rd_st0_419  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[419]), .rdlo_in(a0_wr[931]),  .coef_in(coef[419]), .rdup_out(a1_wr[419]), .rdlo_out(a1_wr[931]));
			radix2 #(.width(width)) rd_st0_420  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[420]), .rdlo_in(a0_wr[932]),  .coef_in(coef[420]), .rdup_out(a1_wr[420]), .rdlo_out(a1_wr[932]));
			radix2 #(.width(width)) rd_st0_421  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[421]), .rdlo_in(a0_wr[933]),  .coef_in(coef[421]), .rdup_out(a1_wr[421]), .rdlo_out(a1_wr[933]));
			radix2 #(.width(width)) rd_st0_422  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[422]), .rdlo_in(a0_wr[934]),  .coef_in(coef[422]), .rdup_out(a1_wr[422]), .rdlo_out(a1_wr[934]));
			radix2 #(.width(width)) rd_st0_423  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[423]), .rdlo_in(a0_wr[935]),  .coef_in(coef[423]), .rdup_out(a1_wr[423]), .rdlo_out(a1_wr[935]));
			radix2 #(.width(width)) rd_st0_424  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[424]), .rdlo_in(a0_wr[936]),  .coef_in(coef[424]), .rdup_out(a1_wr[424]), .rdlo_out(a1_wr[936]));
			radix2 #(.width(width)) rd_st0_425  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[425]), .rdlo_in(a0_wr[937]),  .coef_in(coef[425]), .rdup_out(a1_wr[425]), .rdlo_out(a1_wr[937]));
			radix2 #(.width(width)) rd_st0_426  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[426]), .rdlo_in(a0_wr[938]),  .coef_in(coef[426]), .rdup_out(a1_wr[426]), .rdlo_out(a1_wr[938]));
			radix2 #(.width(width)) rd_st0_427  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[427]), .rdlo_in(a0_wr[939]),  .coef_in(coef[427]), .rdup_out(a1_wr[427]), .rdlo_out(a1_wr[939]));
			radix2 #(.width(width)) rd_st0_428  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[428]), .rdlo_in(a0_wr[940]),  .coef_in(coef[428]), .rdup_out(a1_wr[428]), .rdlo_out(a1_wr[940]));
			radix2 #(.width(width)) rd_st0_429  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[429]), .rdlo_in(a0_wr[941]),  .coef_in(coef[429]), .rdup_out(a1_wr[429]), .rdlo_out(a1_wr[941]));
			radix2 #(.width(width)) rd_st0_430  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[430]), .rdlo_in(a0_wr[942]),  .coef_in(coef[430]), .rdup_out(a1_wr[430]), .rdlo_out(a1_wr[942]));
			radix2 #(.width(width)) rd_st0_431  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[431]), .rdlo_in(a0_wr[943]),  .coef_in(coef[431]), .rdup_out(a1_wr[431]), .rdlo_out(a1_wr[943]));
			radix2 #(.width(width)) rd_st0_432  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[432]), .rdlo_in(a0_wr[944]),  .coef_in(coef[432]), .rdup_out(a1_wr[432]), .rdlo_out(a1_wr[944]));
			radix2 #(.width(width)) rd_st0_433  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[433]), .rdlo_in(a0_wr[945]),  .coef_in(coef[433]), .rdup_out(a1_wr[433]), .rdlo_out(a1_wr[945]));
			radix2 #(.width(width)) rd_st0_434  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[434]), .rdlo_in(a0_wr[946]),  .coef_in(coef[434]), .rdup_out(a1_wr[434]), .rdlo_out(a1_wr[946]));
			radix2 #(.width(width)) rd_st0_435  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[435]), .rdlo_in(a0_wr[947]),  .coef_in(coef[435]), .rdup_out(a1_wr[435]), .rdlo_out(a1_wr[947]));
			radix2 #(.width(width)) rd_st0_436  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[436]), .rdlo_in(a0_wr[948]),  .coef_in(coef[436]), .rdup_out(a1_wr[436]), .rdlo_out(a1_wr[948]));
			radix2 #(.width(width)) rd_st0_437  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[437]), .rdlo_in(a0_wr[949]),  .coef_in(coef[437]), .rdup_out(a1_wr[437]), .rdlo_out(a1_wr[949]));
			radix2 #(.width(width)) rd_st0_438  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[438]), .rdlo_in(a0_wr[950]),  .coef_in(coef[438]), .rdup_out(a1_wr[438]), .rdlo_out(a1_wr[950]));
			radix2 #(.width(width)) rd_st0_439  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[439]), .rdlo_in(a0_wr[951]),  .coef_in(coef[439]), .rdup_out(a1_wr[439]), .rdlo_out(a1_wr[951]));
			radix2 #(.width(width)) rd_st0_440  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[440]), .rdlo_in(a0_wr[952]),  .coef_in(coef[440]), .rdup_out(a1_wr[440]), .rdlo_out(a1_wr[952]));
			radix2 #(.width(width)) rd_st0_441  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[441]), .rdlo_in(a0_wr[953]),  .coef_in(coef[441]), .rdup_out(a1_wr[441]), .rdlo_out(a1_wr[953]));
			radix2 #(.width(width)) rd_st0_442  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[442]), .rdlo_in(a0_wr[954]),  .coef_in(coef[442]), .rdup_out(a1_wr[442]), .rdlo_out(a1_wr[954]));
			radix2 #(.width(width)) rd_st0_443  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[443]), .rdlo_in(a0_wr[955]),  .coef_in(coef[443]), .rdup_out(a1_wr[443]), .rdlo_out(a1_wr[955]));
			radix2 #(.width(width)) rd_st0_444  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[444]), .rdlo_in(a0_wr[956]),  .coef_in(coef[444]), .rdup_out(a1_wr[444]), .rdlo_out(a1_wr[956]));
			radix2 #(.width(width)) rd_st0_445  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[445]), .rdlo_in(a0_wr[957]),  .coef_in(coef[445]), .rdup_out(a1_wr[445]), .rdlo_out(a1_wr[957]));
			radix2 #(.width(width)) rd_st0_446  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[446]), .rdlo_in(a0_wr[958]),  .coef_in(coef[446]), .rdup_out(a1_wr[446]), .rdlo_out(a1_wr[958]));
			radix2 #(.width(width)) rd_st0_447  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[447]), .rdlo_in(a0_wr[959]),  .coef_in(coef[447]), .rdup_out(a1_wr[447]), .rdlo_out(a1_wr[959]));
			radix2 #(.width(width)) rd_st0_448  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[448]), .rdlo_in(a0_wr[960]),  .coef_in(coef[448]), .rdup_out(a1_wr[448]), .rdlo_out(a1_wr[960]));
			radix2 #(.width(width)) rd_st0_449  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[449]), .rdlo_in(a0_wr[961]),  .coef_in(coef[449]), .rdup_out(a1_wr[449]), .rdlo_out(a1_wr[961]));
			radix2 #(.width(width)) rd_st0_450  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[450]), .rdlo_in(a0_wr[962]),  .coef_in(coef[450]), .rdup_out(a1_wr[450]), .rdlo_out(a1_wr[962]));
			radix2 #(.width(width)) rd_st0_451  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[451]), .rdlo_in(a0_wr[963]),  .coef_in(coef[451]), .rdup_out(a1_wr[451]), .rdlo_out(a1_wr[963]));
			radix2 #(.width(width)) rd_st0_452  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[452]), .rdlo_in(a0_wr[964]),  .coef_in(coef[452]), .rdup_out(a1_wr[452]), .rdlo_out(a1_wr[964]));
			radix2 #(.width(width)) rd_st0_453  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[453]), .rdlo_in(a0_wr[965]),  .coef_in(coef[453]), .rdup_out(a1_wr[453]), .rdlo_out(a1_wr[965]));
			radix2 #(.width(width)) rd_st0_454  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[454]), .rdlo_in(a0_wr[966]),  .coef_in(coef[454]), .rdup_out(a1_wr[454]), .rdlo_out(a1_wr[966]));
			radix2 #(.width(width)) rd_st0_455  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[455]), .rdlo_in(a0_wr[967]),  .coef_in(coef[455]), .rdup_out(a1_wr[455]), .rdlo_out(a1_wr[967]));
			radix2 #(.width(width)) rd_st0_456  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[456]), .rdlo_in(a0_wr[968]),  .coef_in(coef[456]), .rdup_out(a1_wr[456]), .rdlo_out(a1_wr[968]));
			radix2 #(.width(width)) rd_st0_457  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[457]), .rdlo_in(a0_wr[969]),  .coef_in(coef[457]), .rdup_out(a1_wr[457]), .rdlo_out(a1_wr[969]));
			radix2 #(.width(width)) rd_st0_458  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[458]), .rdlo_in(a0_wr[970]),  .coef_in(coef[458]), .rdup_out(a1_wr[458]), .rdlo_out(a1_wr[970]));
			radix2 #(.width(width)) rd_st0_459  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[459]), .rdlo_in(a0_wr[971]),  .coef_in(coef[459]), .rdup_out(a1_wr[459]), .rdlo_out(a1_wr[971]));
			radix2 #(.width(width)) rd_st0_460  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[460]), .rdlo_in(a0_wr[972]),  .coef_in(coef[460]), .rdup_out(a1_wr[460]), .rdlo_out(a1_wr[972]));
			radix2 #(.width(width)) rd_st0_461  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[461]), .rdlo_in(a0_wr[973]),  .coef_in(coef[461]), .rdup_out(a1_wr[461]), .rdlo_out(a1_wr[973]));
			radix2 #(.width(width)) rd_st0_462  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[462]), .rdlo_in(a0_wr[974]),  .coef_in(coef[462]), .rdup_out(a1_wr[462]), .rdlo_out(a1_wr[974]));
			radix2 #(.width(width)) rd_st0_463  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[463]), .rdlo_in(a0_wr[975]),  .coef_in(coef[463]), .rdup_out(a1_wr[463]), .rdlo_out(a1_wr[975]));
			radix2 #(.width(width)) rd_st0_464  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[464]), .rdlo_in(a0_wr[976]),  .coef_in(coef[464]), .rdup_out(a1_wr[464]), .rdlo_out(a1_wr[976]));
			radix2 #(.width(width)) rd_st0_465  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[465]), .rdlo_in(a0_wr[977]),  .coef_in(coef[465]), .rdup_out(a1_wr[465]), .rdlo_out(a1_wr[977]));
			radix2 #(.width(width)) rd_st0_466  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[466]), .rdlo_in(a0_wr[978]),  .coef_in(coef[466]), .rdup_out(a1_wr[466]), .rdlo_out(a1_wr[978]));
			radix2 #(.width(width)) rd_st0_467  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[467]), .rdlo_in(a0_wr[979]),  .coef_in(coef[467]), .rdup_out(a1_wr[467]), .rdlo_out(a1_wr[979]));
			radix2 #(.width(width)) rd_st0_468  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[468]), .rdlo_in(a0_wr[980]),  .coef_in(coef[468]), .rdup_out(a1_wr[468]), .rdlo_out(a1_wr[980]));
			radix2 #(.width(width)) rd_st0_469  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[469]), .rdlo_in(a0_wr[981]),  .coef_in(coef[469]), .rdup_out(a1_wr[469]), .rdlo_out(a1_wr[981]));
			radix2 #(.width(width)) rd_st0_470  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[470]), .rdlo_in(a0_wr[982]),  .coef_in(coef[470]), .rdup_out(a1_wr[470]), .rdlo_out(a1_wr[982]));
			radix2 #(.width(width)) rd_st0_471  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[471]), .rdlo_in(a0_wr[983]),  .coef_in(coef[471]), .rdup_out(a1_wr[471]), .rdlo_out(a1_wr[983]));
			radix2 #(.width(width)) rd_st0_472  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[472]), .rdlo_in(a0_wr[984]),  .coef_in(coef[472]), .rdup_out(a1_wr[472]), .rdlo_out(a1_wr[984]));
			radix2 #(.width(width)) rd_st0_473  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[473]), .rdlo_in(a0_wr[985]),  .coef_in(coef[473]), .rdup_out(a1_wr[473]), .rdlo_out(a1_wr[985]));
			radix2 #(.width(width)) rd_st0_474  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[474]), .rdlo_in(a0_wr[986]),  .coef_in(coef[474]), .rdup_out(a1_wr[474]), .rdlo_out(a1_wr[986]));
			radix2 #(.width(width)) rd_st0_475  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[475]), .rdlo_in(a0_wr[987]),  .coef_in(coef[475]), .rdup_out(a1_wr[475]), .rdlo_out(a1_wr[987]));
			radix2 #(.width(width)) rd_st0_476  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[476]), .rdlo_in(a0_wr[988]),  .coef_in(coef[476]), .rdup_out(a1_wr[476]), .rdlo_out(a1_wr[988]));
			radix2 #(.width(width)) rd_st0_477  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[477]), .rdlo_in(a0_wr[989]),  .coef_in(coef[477]), .rdup_out(a1_wr[477]), .rdlo_out(a1_wr[989]));
			radix2 #(.width(width)) rd_st0_478  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[478]), .rdlo_in(a0_wr[990]),  .coef_in(coef[478]), .rdup_out(a1_wr[478]), .rdlo_out(a1_wr[990]));
			radix2 #(.width(width)) rd_st0_479  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[479]), .rdlo_in(a0_wr[991]),  .coef_in(coef[479]), .rdup_out(a1_wr[479]), .rdlo_out(a1_wr[991]));
			radix2 #(.width(width)) rd_st0_480  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[480]), .rdlo_in(a0_wr[992]),  .coef_in(coef[480]), .rdup_out(a1_wr[480]), .rdlo_out(a1_wr[992]));
			radix2 #(.width(width)) rd_st0_481  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[481]), .rdlo_in(a0_wr[993]),  .coef_in(coef[481]), .rdup_out(a1_wr[481]), .rdlo_out(a1_wr[993]));
			radix2 #(.width(width)) rd_st0_482  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[482]), .rdlo_in(a0_wr[994]),  .coef_in(coef[482]), .rdup_out(a1_wr[482]), .rdlo_out(a1_wr[994]));
			radix2 #(.width(width)) rd_st0_483  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[483]), .rdlo_in(a0_wr[995]),  .coef_in(coef[483]), .rdup_out(a1_wr[483]), .rdlo_out(a1_wr[995]));
			radix2 #(.width(width)) rd_st0_484  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[484]), .rdlo_in(a0_wr[996]),  .coef_in(coef[484]), .rdup_out(a1_wr[484]), .rdlo_out(a1_wr[996]));
			radix2 #(.width(width)) rd_st0_485  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[485]), .rdlo_in(a0_wr[997]),  .coef_in(coef[485]), .rdup_out(a1_wr[485]), .rdlo_out(a1_wr[997]));
			radix2 #(.width(width)) rd_st0_486  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[486]), .rdlo_in(a0_wr[998]),  .coef_in(coef[486]), .rdup_out(a1_wr[486]), .rdlo_out(a1_wr[998]));
			radix2 #(.width(width)) rd_st0_487  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[487]), .rdlo_in(a0_wr[999]),  .coef_in(coef[487]), .rdup_out(a1_wr[487]), .rdlo_out(a1_wr[999]));
			radix2 #(.width(width)) rd_st0_488  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[488]), .rdlo_in(a0_wr[1000]),  .coef_in(coef[488]), .rdup_out(a1_wr[488]), .rdlo_out(a1_wr[1000]));
			radix2 #(.width(width)) rd_st0_489  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[489]), .rdlo_in(a0_wr[1001]),  .coef_in(coef[489]), .rdup_out(a1_wr[489]), .rdlo_out(a1_wr[1001]));
			radix2 #(.width(width)) rd_st0_490  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[490]), .rdlo_in(a0_wr[1002]),  .coef_in(coef[490]), .rdup_out(a1_wr[490]), .rdlo_out(a1_wr[1002]));
			radix2 #(.width(width)) rd_st0_491  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[491]), .rdlo_in(a0_wr[1003]),  .coef_in(coef[491]), .rdup_out(a1_wr[491]), .rdlo_out(a1_wr[1003]));
			radix2 #(.width(width)) rd_st0_492  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[492]), .rdlo_in(a0_wr[1004]),  .coef_in(coef[492]), .rdup_out(a1_wr[492]), .rdlo_out(a1_wr[1004]));
			radix2 #(.width(width)) rd_st0_493  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[493]), .rdlo_in(a0_wr[1005]),  .coef_in(coef[493]), .rdup_out(a1_wr[493]), .rdlo_out(a1_wr[1005]));
			radix2 #(.width(width)) rd_st0_494  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[494]), .rdlo_in(a0_wr[1006]),  .coef_in(coef[494]), .rdup_out(a1_wr[494]), .rdlo_out(a1_wr[1006]));
			radix2 #(.width(width)) rd_st0_495  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[495]), .rdlo_in(a0_wr[1007]),  .coef_in(coef[495]), .rdup_out(a1_wr[495]), .rdlo_out(a1_wr[1007]));
			radix2 #(.width(width)) rd_st0_496  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[496]), .rdlo_in(a0_wr[1008]),  .coef_in(coef[496]), .rdup_out(a1_wr[496]), .rdlo_out(a1_wr[1008]));
			radix2 #(.width(width)) rd_st0_497  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[497]), .rdlo_in(a0_wr[1009]),  .coef_in(coef[497]), .rdup_out(a1_wr[497]), .rdlo_out(a1_wr[1009]));
			radix2 #(.width(width)) rd_st0_498  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[498]), .rdlo_in(a0_wr[1010]),  .coef_in(coef[498]), .rdup_out(a1_wr[498]), .rdlo_out(a1_wr[1010]));
			radix2 #(.width(width)) rd_st0_499  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[499]), .rdlo_in(a0_wr[1011]),  .coef_in(coef[499]), .rdup_out(a1_wr[499]), .rdlo_out(a1_wr[1011]));
			radix2 #(.width(width)) rd_st0_500  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[500]), .rdlo_in(a0_wr[1012]),  .coef_in(coef[500]), .rdup_out(a1_wr[500]), .rdlo_out(a1_wr[1012]));
			radix2 #(.width(width)) rd_st0_501  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[501]), .rdlo_in(a0_wr[1013]),  .coef_in(coef[501]), .rdup_out(a1_wr[501]), .rdlo_out(a1_wr[1013]));
			radix2 #(.width(width)) rd_st0_502  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[502]), .rdlo_in(a0_wr[1014]),  .coef_in(coef[502]), .rdup_out(a1_wr[502]), .rdlo_out(a1_wr[1014]));
			radix2 #(.width(width)) rd_st0_503  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[503]), .rdlo_in(a0_wr[1015]),  .coef_in(coef[503]), .rdup_out(a1_wr[503]), .rdlo_out(a1_wr[1015]));
			radix2 #(.width(width)) rd_st0_504  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[504]), .rdlo_in(a0_wr[1016]),  .coef_in(coef[504]), .rdup_out(a1_wr[504]), .rdlo_out(a1_wr[1016]));
			radix2 #(.width(width)) rd_st0_505  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[505]), .rdlo_in(a0_wr[1017]),  .coef_in(coef[505]), .rdup_out(a1_wr[505]), .rdlo_out(a1_wr[1017]));
			radix2 #(.width(width)) rd_st0_506  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[506]), .rdlo_in(a0_wr[1018]),  .coef_in(coef[506]), .rdup_out(a1_wr[506]), .rdlo_out(a1_wr[1018]));
			radix2 #(.width(width)) rd_st0_507  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[507]), .rdlo_in(a0_wr[1019]),  .coef_in(coef[507]), .rdup_out(a1_wr[507]), .rdlo_out(a1_wr[1019]));
			radix2 #(.width(width)) rd_st0_508  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[508]), .rdlo_in(a0_wr[1020]),  .coef_in(coef[508]), .rdup_out(a1_wr[508]), .rdlo_out(a1_wr[1020]));
			radix2 #(.width(width)) rd_st0_509  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[509]), .rdlo_in(a0_wr[1021]),  .coef_in(coef[509]), .rdup_out(a1_wr[509]), .rdlo_out(a1_wr[1021]));
			radix2 #(.width(width)) rd_st0_510  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[510]), .rdlo_in(a0_wr[1022]),  .coef_in(coef[510]), .rdup_out(a1_wr[510]), .rdlo_out(a1_wr[1022]));
			radix2 #(.width(width)) rd_st0_511  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[511]), .rdlo_in(a0_wr[1023]),  .coef_in(coef[511]), .rdup_out(a1_wr[511]), .rdlo_out(a1_wr[1023]));

		//--- radix stage 1
			radix2 #(.width(width)) rd_st1_0   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[0]), .rdlo_in(a1_wr[256]),  .coef_in(coef[0]), .rdup_out(a2_wr[0]), .rdlo_out(a2_wr[256]));
			radix2 #(.width(width)) rd_st1_1   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1]), .rdlo_in(a1_wr[257]),  .coef_in(coef[2]), .rdup_out(a2_wr[1]), .rdlo_out(a2_wr[257]));
			radix2 #(.width(width)) rd_st1_2   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[2]), .rdlo_in(a1_wr[258]),  .coef_in(coef[4]), .rdup_out(a2_wr[2]), .rdlo_out(a2_wr[258]));
			radix2 #(.width(width)) rd_st1_3   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[3]), .rdlo_in(a1_wr[259]),  .coef_in(coef[6]), .rdup_out(a2_wr[3]), .rdlo_out(a2_wr[259]));
			radix2 #(.width(width)) rd_st1_4   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[4]), .rdlo_in(a1_wr[260]),  .coef_in(coef[8]), .rdup_out(a2_wr[4]), .rdlo_out(a2_wr[260]));
			radix2 #(.width(width)) rd_st1_5   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[5]), .rdlo_in(a1_wr[261]),  .coef_in(coef[10]), .rdup_out(a2_wr[5]), .rdlo_out(a2_wr[261]));
			radix2 #(.width(width)) rd_st1_6   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[6]), .rdlo_in(a1_wr[262]),  .coef_in(coef[12]), .rdup_out(a2_wr[6]), .rdlo_out(a2_wr[262]));
			radix2 #(.width(width)) rd_st1_7   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[7]), .rdlo_in(a1_wr[263]),  .coef_in(coef[14]), .rdup_out(a2_wr[7]), .rdlo_out(a2_wr[263]));
			radix2 #(.width(width)) rd_st1_8   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[8]), .rdlo_in(a1_wr[264]),  .coef_in(coef[16]), .rdup_out(a2_wr[8]), .rdlo_out(a2_wr[264]));
			radix2 #(.width(width)) rd_st1_9   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[9]), .rdlo_in(a1_wr[265]),  .coef_in(coef[18]), .rdup_out(a2_wr[9]), .rdlo_out(a2_wr[265]));
			radix2 #(.width(width)) rd_st1_10  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[10]), .rdlo_in(a1_wr[266]),  .coef_in(coef[20]), .rdup_out(a2_wr[10]), .rdlo_out(a2_wr[266]));
			radix2 #(.width(width)) rd_st1_11  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[11]), .rdlo_in(a1_wr[267]),  .coef_in(coef[22]), .rdup_out(a2_wr[11]), .rdlo_out(a2_wr[267]));
			radix2 #(.width(width)) rd_st1_12  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[12]), .rdlo_in(a1_wr[268]),  .coef_in(coef[24]), .rdup_out(a2_wr[12]), .rdlo_out(a2_wr[268]));
			radix2 #(.width(width)) rd_st1_13  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[13]), .rdlo_in(a1_wr[269]),  .coef_in(coef[26]), .rdup_out(a2_wr[13]), .rdlo_out(a2_wr[269]));
			radix2 #(.width(width)) rd_st1_14  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[14]), .rdlo_in(a1_wr[270]),  .coef_in(coef[28]), .rdup_out(a2_wr[14]), .rdlo_out(a2_wr[270]));
			radix2 #(.width(width)) rd_st1_15  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[15]), .rdlo_in(a1_wr[271]),  .coef_in(coef[30]), .rdup_out(a2_wr[15]), .rdlo_out(a2_wr[271]));
			radix2 #(.width(width)) rd_st1_16  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[16]), .rdlo_in(a1_wr[272]),  .coef_in(coef[32]), .rdup_out(a2_wr[16]), .rdlo_out(a2_wr[272]));
			radix2 #(.width(width)) rd_st1_17  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[17]), .rdlo_in(a1_wr[273]),  .coef_in(coef[34]), .rdup_out(a2_wr[17]), .rdlo_out(a2_wr[273]));
			radix2 #(.width(width)) rd_st1_18  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[18]), .rdlo_in(a1_wr[274]),  .coef_in(coef[36]), .rdup_out(a2_wr[18]), .rdlo_out(a2_wr[274]));
			radix2 #(.width(width)) rd_st1_19  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[19]), .rdlo_in(a1_wr[275]),  .coef_in(coef[38]), .rdup_out(a2_wr[19]), .rdlo_out(a2_wr[275]));
			radix2 #(.width(width)) rd_st1_20  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[20]), .rdlo_in(a1_wr[276]),  .coef_in(coef[40]), .rdup_out(a2_wr[20]), .rdlo_out(a2_wr[276]));
			radix2 #(.width(width)) rd_st1_21  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[21]), .rdlo_in(a1_wr[277]),  .coef_in(coef[42]), .rdup_out(a2_wr[21]), .rdlo_out(a2_wr[277]));
			radix2 #(.width(width)) rd_st1_22  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[22]), .rdlo_in(a1_wr[278]),  .coef_in(coef[44]), .rdup_out(a2_wr[22]), .rdlo_out(a2_wr[278]));
			radix2 #(.width(width)) rd_st1_23  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[23]), .rdlo_in(a1_wr[279]),  .coef_in(coef[46]), .rdup_out(a2_wr[23]), .rdlo_out(a2_wr[279]));
			radix2 #(.width(width)) rd_st1_24  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[24]), .rdlo_in(a1_wr[280]),  .coef_in(coef[48]), .rdup_out(a2_wr[24]), .rdlo_out(a2_wr[280]));
			radix2 #(.width(width)) rd_st1_25  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[25]), .rdlo_in(a1_wr[281]),  .coef_in(coef[50]), .rdup_out(a2_wr[25]), .rdlo_out(a2_wr[281]));
			radix2 #(.width(width)) rd_st1_26  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[26]), .rdlo_in(a1_wr[282]),  .coef_in(coef[52]), .rdup_out(a2_wr[26]), .rdlo_out(a2_wr[282]));
			radix2 #(.width(width)) rd_st1_27  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[27]), .rdlo_in(a1_wr[283]),  .coef_in(coef[54]), .rdup_out(a2_wr[27]), .rdlo_out(a2_wr[283]));
			radix2 #(.width(width)) rd_st1_28  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[28]), .rdlo_in(a1_wr[284]),  .coef_in(coef[56]), .rdup_out(a2_wr[28]), .rdlo_out(a2_wr[284]));
			radix2 #(.width(width)) rd_st1_29  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[29]), .rdlo_in(a1_wr[285]),  .coef_in(coef[58]), .rdup_out(a2_wr[29]), .rdlo_out(a2_wr[285]));
			radix2 #(.width(width)) rd_st1_30  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[30]), .rdlo_in(a1_wr[286]),  .coef_in(coef[60]), .rdup_out(a2_wr[30]), .rdlo_out(a2_wr[286]));
			radix2 #(.width(width)) rd_st1_31  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[31]), .rdlo_in(a1_wr[287]),  .coef_in(coef[62]), .rdup_out(a2_wr[31]), .rdlo_out(a2_wr[287]));
			radix2 #(.width(width)) rd_st1_32  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[32]), .rdlo_in(a1_wr[288]),  .coef_in(coef[64]), .rdup_out(a2_wr[32]), .rdlo_out(a2_wr[288]));
			radix2 #(.width(width)) rd_st1_33  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[33]), .rdlo_in(a1_wr[289]),  .coef_in(coef[66]), .rdup_out(a2_wr[33]), .rdlo_out(a2_wr[289]));
			radix2 #(.width(width)) rd_st1_34  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[34]), .rdlo_in(a1_wr[290]),  .coef_in(coef[68]), .rdup_out(a2_wr[34]), .rdlo_out(a2_wr[290]));
			radix2 #(.width(width)) rd_st1_35  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[35]), .rdlo_in(a1_wr[291]),  .coef_in(coef[70]), .rdup_out(a2_wr[35]), .rdlo_out(a2_wr[291]));
			radix2 #(.width(width)) rd_st1_36  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[36]), .rdlo_in(a1_wr[292]),  .coef_in(coef[72]), .rdup_out(a2_wr[36]), .rdlo_out(a2_wr[292]));
			radix2 #(.width(width)) rd_st1_37  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[37]), .rdlo_in(a1_wr[293]),  .coef_in(coef[74]), .rdup_out(a2_wr[37]), .rdlo_out(a2_wr[293]));
			radix2 #(.width(width)) rd_st1_38  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[38]), .rdlo_in(a1_wr[294]),  .coef_in(coef[76]), .rdup_out(a2_wr[38]), .rdlo_out(a2_wr[294]));
			radix2 #(.width(width)) rd_st1_39  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[39]), .rdlo_in(a1_wr[295]),  .coef_in(coef[78]), .rdup_out(a2_wr[39]), .rdlo_out(a2_wr[295]));
			radix2 #(.width(width)) rd_st1_40  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[40]), .rdlo_in(a1_wr[296]),  .coef_in(coef[80]), .rdup_out(a2_wr[40]), .rdlo_out(a2_wr[296]));
			radix2 #(.width(width)) rd_st1_41  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[41]), .rdlo_in(a1_wr[297]),  .coef_in(coef[82]), .rdup_out(a2_wr[41]), .rdlo_out(a2_wr[297]));
			radix2 #(.width(width)) rd_st1_42  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[42]), .rdlo_in(a1_wr[298]),  .coef_in(coef[84]), .rdup_out(a2_wr[42]), .rdlo_out(a2_wr[298]));
			radix2 #(.width(width)) rd_st1_43  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[43]), .rdlo_in(a1_wr[299]),  .coef_in(coef[86]), .rdup_out(a2_wr[43]), .rdlo_out(a2_wr[299]));
			radix2 #(.width(width)) rd_st1_44  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[44]), .rdlo_in(a1_wr[300]),  .coef_in(coef[88]), .rdup_out(a2_wr[44]), .rdlo_out(a2_wr[300]));
			radix2 #(.width(width)) rd_st1_45  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[45]), .rdlo_in(a1_wr[301]),  .coef_in(coef[90]), .rdup_out(a2_wr[45]), .rdlo_out(a2_wr[301]));
			radix2 #(.width(width)) rd_st1_46  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[46]), .rdlo_in(a1_wr[302]),  .coef_in(coef[92]), .rdup_out(a2_wr[46]), .rdlo_out(a2_wr[302]));
			radix2 #(.width(width)) rd_st1_47  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[47]), .rdlo_in(a1_wr[303]),  .coef_in(coef[94]), .rdup_out(a2_wr[47]), .rdlo_out(a2_wr[303]));
			radix2 #(.width(width)) rd_st1_48  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[48]), .rdlo_in(a1_wr[304]),  .coef_in(coef[96]), .rdup_out(a2_wr[48]), .rdlo_out(a2_wr[304]));
			radix2 #(.width(width)) rd_st1_49  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[49]), .rdlo_in(a1_wr[305]),  .coef_in(coef[98]), .rdup_out(a2_wr[49]), .rdlo_out(a2_wr[305]));
			radix2 #(.width(width)) rd_st1_50  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[50]), .rdlo_in(a1_wr[306]),  .coef_in(coef[100]), .rdup_out(a2_wr[50]), .rdlo_out(a2_wr[306]));
			radix2 #(.width(width)) rd_st1_51  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[51]), .rdlo_in(a1_wr[307]),  .coef_in(coef[102]), .rdup_out(a2_wr[51]), .rdlo_out(a2_wr[307]));
			radix2 #(.width(width)) rd_st1_52  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[52]), .rdlo_in(a1_wr[308]),  .coef_in(coef[104]), .rdup_out(a2_wr[52]), .rdlo_out(a2_wr[308]));
			radix2 #(.width(width)) rd_st1_53  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[53]), .rdlo_in(a1_wr[309]),  .coef_in(coef[106]), .rdup_out(a2_wr[53]), .rdlo_out(a2_wr[309]));
			radix2 #(.width(width)) rd_st1_54  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[54]), .rdlo_in(a1_wr[310]),  .coef_in(coef[108]), .rdup_out(a2_wr[54]), .rdlo_out(a2_wr[310]));
			radix2 #(.width(width)) rd_st1_55  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[55]), .rdlo_in(a1_wr[311]),  .coef_in(coef[110]), .rdup_out(a2_wr[55]), .rdlo_out(a2_wr[311]));
			radix2 #(.width(width)) rd_st1_56  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[56]), .rdlo_in(a1_wr[312]),  .coef_in(coef[112]), .rdup_out(a2_wr[56]), .rdlo_out(a2_wr[312]));
			radix2 #(.width(width)) rd_st1_57  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[57]), .rdlo_in(a1_wr[313]),  .coef_in(coef[114]), .rdup_out(a2_wr[57]), .rdlo_out(a2_wr[313]));
			radix2 #(.width(width)) rd_st1_58  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[58]), .rdlo_in(a1_wr[314]),  .coef_in(coef[116]), .rdup_out(a2_wr[58]), .rdlo_out(a2_wr[314]));
			radix2 #(.width(width)) rd_st1_59  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[59]), .rdlo_in(a1_wr[315]),  .coef_in(coef[118]), .rdup_out(a2_wr[59]), .rdlo_out(a2_wr[315]));
			radix2 #(.width(width)) rd_st1_60  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[60]), .rdlo_in(a1_wr[316]),  .coef_in(coef[120]), .rdup_out(a2_wr[60]), .rdlo_out(a2_wr[316]));
			radix2 #(.width(width)) rd_st1_61  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[61]), .rdlo_in(a1_wr[317]),  .coef_in(coef[122]), .rdup_out(a2_wr[61]), .rdlo_out(a2_wr[317]));
			radix2 #(.width(width)) rd_st1_62  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[62]), .rdlo_in(a1_wr[318]),  .coef_in(coef[124]), .rdup_out(a2_wr[62]), .rdlo_out(a2_wr[318]));
			radix2 #(.width(width)) rd_st1_63  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[63]), .rdlo_in(a1_wr[319]),  .coef_in(coef[126]), .rdup_out(a2_wr[63]), .rdlo_out(a2_wr[319]));
			radix2 #(.width(width)) rd_st1_64  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[64]), .rdlo_in(a1_wr[320]),  .coef_in(coef[128]), .rdup_out(a2_wr[64]), .rdlo_out(a2_wr[320]));
			radix2 #(.width(width)) rd_st1_65  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[65]), .rdlo_in(a1_wr[321]),  .coef_in(coef[130]), .rdup_out(a2_wr[65]), .rdlo_out(a2_wr[321]));
			radix2 #(.width(width)) rd_st1_66  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[66]), .rdlo_in(a1_wr[322]),  .coef_in(coef[132]), .rdup_out(a2_wr[66]), .rdlo_out(a2_wr[322]));
			radix2 #(.width(width)) rd_st1_67  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[67]), .rdlo_in(a1_wr[323]),  .coef_in(coef[134]), .rdup_out(a2_wr[67]), .rdlo_out(a2_wr[323]));
			radix2 #(.width(width)) rd_st1_68  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[68]), .rdlo_in(a1_wr[324]),  .coef_in(coef[136]), .rdup_out(a2_wr[68]), .rdlo_out(a2_wr[324]));
			radix2 #(.width(width)) rd_st1_69  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[69]), .rdlo_in(a1_wr[325]),  .coef_in(coef[138]), .rdup_out(a2_wr[69]), .rdlo_out(a2_wr[325]));
			radix2 #(.width(width)) rd_st1_70  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[70]), .rdlo_in(a1_wr[326]),  .coef_in(coef[140]), .rdup_out(a2_wr[70]), .rdlo_out(a2_wr[326]));
			radix2 #(.width(width)) rd_st1_71  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[71]), .rdlo_in(a1_wr[327]),  .coef_in(coef[142]), .rdup_out(a2_wr[71]), .rdlo_out(a2_wr[327]));
			radix2 #(.width(width)) rd_st1_72  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[72]), .rdlo_in(a1_wr[328]),  .coef_in(coef[144]), .rdup_out(a2_wr[72]), .rdlo_out(a2_wr[328]));
			radix2 #(.width(width)) rd_st1_73  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[73]), .rdlo_in(a1_wr[329]),  .coef_in(coef[146]), .rdup_out(a2_wr[73]), .rdlo_out(a2_wr[329]));
			radix2 #(.width(width)) rd_st1_74  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[74]), .rdlo_in(a1_wr[330]),  .coef_in(coef[148]), .rdup_out(a2_wr[74]), .rdlo_out(a2_wr[330]));
			radix2 #(.width(width)) rd_st1_75  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[75]), .rdlo_in(a1_wr[331]),  .coef_in(coef[150]), .rdup_out(a2_wr[75]), .rdlo_out(a2_wr[331]));
			radix2 #(.width(width)) rd_st1_76  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[76]), .rdlo_in(a1_wr[332]),  .coef_in(coef[152]), .rdup_out(a2_wr[76]), .rdlo_out(a2_wr[332]));
			radix2 #(.width(width)) rd_st1_77  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[77]), .rdlo_in(a1_wr[333]),  .coef_in(coef[154]), .rdup_out(a2_wr[77]), .rdlo_out(a2_wr[333]));
			radix2 #(.width(width)) rd_st1_78  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[78]), .rdlo_in(a1_wr[334]),  .coef_in(coef[156]), .rdup_out(a2_wr[78]), .rdlo_out(a2_wr[334]));
			radix2 #(.width(width)) rd_st1_79  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[79]), .rdlo_in(a1_wr[335]),  .coef_in(coef[158]), .rdup_out(a2_wr[79]), .rdlo_out(a2_wr[335]));
			radix2 #(.width(width)) rd_st1_80  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[80]), .rdlo_in(a1_wr[336]),  .coef_in(coef[160]), .rdup_out(a2_wr[80]), .rdlo_out(a2_wr[336]));
			radix2 #(.width(width)) rd_st1_81  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[81]), .rdlo_in(a1_wr[337]),  .coef_in(coef[162]), .rdup_out(a2_wr[81]), .rdlo_out(a2_wr[337]));
			radix2 #(.width(width)) rd_st1_82  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[82]), .rdlo_in(a1_wr[338]),  .coef_in(coef[164]), .rdup_out(a2_wr[82]), .rdlo_out(a2_wr[338]));
			radix2 #(.width(width)) rd_st1_83  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[83]), .rdlo_in(a1_wr[339]),  .coef_in(coef[166]), .rdup_out(a2_wr[83]), .rdlo_out(a2_wr[339]));
			radix2 #(.width(width)) rd_st1_84  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[84]), .rdlo_in(a1_wr[340]),  .coef_in(coef[168]), .rdup_out(a2_wr[84]), .rdlo_out(a2_wr[340]));
			radix2 #(.width(width)) rd_st1_85  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[85]), .rdlo_in(a1_wr[341]),  .coef_in(coef[170]), .rdup_out(a2_wr[85]), .rdlo_out(a2_wr[341]));
			radix2 #(.width(width)) rd_st1_86  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[86]), .rdlo_in(a1_wr[342]),  .coef_in(coef[172]), .rdup_out(a2_wr[86]), .rdlo_out(a2_wr[342]));
			radix2 #(.width(width)) rd_st1_87  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[87]), .rdlo_in(a1_wr[343]),  .coef_in(coef[174]), .rdup_out(a2_wr[87]), .rdlo_out(a2_wr[343]));
			radix2 #(.width(width)) rd_st1_88  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[88]), .rdlo_in(a1_wr[344]),  .coef_in(coef[176]), .rdup_out(a2_wr[88]), .rdlo_out(a2_wr[344]));
			radix2 #(.width(width)) rd_st1_89  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[89]), .rdlo_in(a1_wr[345]),  .coef_in(coef[178]), .rdup_out(a2_wr[89]), .rdlo_out(a2_wr[345]));
			radix2 #(.width(width)) rd_st1_90  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[90]), .rdlo_in(a1_wr[346]),  .coef_in(coef[180]), .rdup_out(a2_wr[90]), .rdlo_out(a2_wr[346]));
			radix2 #(.width(width)) rd_st1_91  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[91]), .rdlo_in(a1_wr[347]),  .coef_in(coef[182]), .rdup_out(a2_wr[91]), .rdlo_out(a2_wr[347]));
			radix2 #(.width(width)) rd_st1_92  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[92]), .rdlo_in(a1_wr[348]),  .coef_in(coef[184]), .rdup_out(a2_wr[92]), .rdlo_out(a2_wr[348]));
			radix2 #(.width(width)) rd_st1_93  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[93]), .rdlo_in(a1_wr[349]),  .coef_in(coef[186]), .rdup_out(a2_wr[93]), .rdlo_out(a2_wr[349]));
			radix2 #(.width(width)) rd_st1_94  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[94]), .rdlo_in(a1_wr[350]),  .coef_in(coef[188]), .rdup_out(a2_wr[94]), .rdlo_out(a2_wr[350]));
			radix2 #(.width(width)) rd_st1_95  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[95]), .rdlo_in(a1_wr[351]),  .coef_in(coef[190]), .rdup_out(a2_wr[95]), .rdlo_out(a2_wr[351]));
			radix2 #(.width(width)) rd_st1_96  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[96]), .rdlo_in(a1_wr[352]),  .coef_in(coef[192]), .rdup_out(a2_wr[96]), .rdlo_out(a2_wr[352]));
			radix2 #(.width(width)) rd_st1_97  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[97]), .rdlo_in(a1_wr[353]),  .coef_in(coef[194]), .rdup_out(a2_wr[97]), .rdlo_out(a2_wr[353]));
			radix2 #(.width(width)) rd_st1_98  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[98]), .rdlo_in(a1_wr[354]),  .coef_in(coef[196]), .rdup_out(a2_wr[98]), .rdlo_out(a2_wr[354]));
			radix2 #(.width(width)) rd_st1_99  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[99]), .rdlo_in(a1_wr[355]),  .coef_in(coef[198]), .rdup_out(a2_wr[99]), .rdlo_out(a2_wr[355]));
			radix2 #(.width(width)) rd_st1_100  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[100]), .rdlo_in(a1_wr[356]),  .coef_in(coef[200]), .rdup_out(a2_wr[100]), .rdlo_out(a2_wr[356]));
			radix2 #(.width(width)) rd_st1_101  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[101]), .rdlo_in(a1_wr[357]),  .coef_in(coef[202]), .rdup_out(a2_wr[101]), .rdlo_out(a2_wr[357]));
			radix2 #(.width(width)) rd_st1_102  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[102]), .rdlo_in(a1_wr[358]),  .coef_in(coef[204]), .rdup_out(a2_wr[102]), .rdlo_out(a2_wr[358]));
			radix2 #(.width(width)) rd_st1_103  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[103]), .rdlo_in(a1_wr[359]),  .coef_in(coef[206]), .rdup_out(a2_wr[103]), .rdlo_out(a2_wr[359]));
			radix2 #(.width(width)) rd_st1_104  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[104]), .rdlo_in(a1_wr[360]),  .coef_in(coef[208]), .rdup_out(a2_wr[104]), .rdlo_out(a2_wr[360]));
			radix2 #(.width(width)) rd_st1_105  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[105]), .rdlo_in(a1_wr[361]),  .coef_in(coef[210]), .rdup_out(a2_wr[105]), .rdlo_out(a2_wr[361]));
			radix2 #(.width(width)) rd_st1_106  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[106]), .rdlo_in(a1_wr[362]),  .coef_in(coef[212]), .rdup_out(a2_wr[106]), .rdlo_out(a2_wr[362]));
			radix2 #(.width(width)) rd_st1_107  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[107]), .rdlo_in(a1_wr[363]),  .coef_in(coef[214]), .rdup_out(a2_wr[107]), .rdlo_out(a2_wr[363]));
			radix2 #(.width(width)) rd_st1_108  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[108]), .rdlo_in(a1_wr[364]),  .coef_in(coef[216]), .rdup_out(a2_wr[108]), .rdlo_out(a2_wr[364]));
			radix2 #(.width(width)) rd_st1_109  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[109]), .rdlo_in(a1_wr[365]),  .coef_in(coef[218]), .rdup_out(a2_wr[109]), .rdlo_out(a2_wr[365]));
			radix2 #(.width(width)) rd_st1_110  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[110]), .rdlo_in(a1_wr[366]),  .coef_in(coef[220]), .rdup_out(a2_wr[110]), .rdlo_out(a2_wr[366]));
			radix2 #(.width(width)) rd_st1_111  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[111]), .rdlo_in(a1_wr[367]),  .coef_in(coef[222]), .rdup_out(a2_wr[111]), .rdlo_out(a2_wr[367]));
			radix2 #(.width(width)) rd_st1_112  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[112]), .rdlo_in(a1_wr[368]),  .coef_in(coef[224]), .rdup_out(a2_wr[112]), .rdlo_out(a2_wr[368]));
			radix2 #(.width(width)) rd_st1_113  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[113]), .rdlo_in(a1_wr[369]),  .coef_in(coef[226]), .rdup_out(a2_wr[113]), .rdlo_out(a2_wr[369]));
			radix2 #(.width(width)) rd_st1_114  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[114]), .rdlo_in(a1_wr[370]),  .coef_in(coef[228]), .rdup_out(a2_wr[114]), .rdlo_out(a2_wr[370]));
			radix2 #(.width(width)) rd_st1_115  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[115]), .rdlo_in(a1_wr[371]),  .coef_in(coef[230]), .rdup_out(a2_wr[115]), .rdlo_out(a2_wr[371]));
			radix2 #(.width(width)) rd_st1_116  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[116]), .rdlo_in(a1_wr[372]),  .coef_in(coef[232]), .rdup_out(a2_wr[116]), .rdlo_out(a2_wr[372]));
			radix2 #(.width(width)) rd_st1_117  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[117]), .rdlo_in(a1_wr[373]),  .coef_in(coef[234]), .rdup_out(a2_wr[117]), .rdlo_out(a2_wr[373]));
			radix2 #(.width(width)) rd_st1_118  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[118]), .rdlo_in(a1_wr[374]),  .coef_in(coef[236]), .rdup_out(a2_wr[118]), .rdlo_out(a2_wr[374]));
			radix2 #(.width(width)) rd_st1_119  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[119]), .rdlo_in(a1_wr[375]),  .coef_in(coef[238]), .rdup_out(a2_wr[119]), .rdlo_out(a2_wr[375]));
			radix2 #(.width(width)) rd_st1_120  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[120]), .rdlo_in(a1_wr[376]),  .coef_in(coef[240]), .rdup_out(a2_wr[120]), .rdlo_out(a2_wr[376]));
			radix2 #(.width(width)) rd_st1_121  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[121]), .rdlo_in(a1_wr[377]),  .coef_in(coef[242]), .rdup_out(a2_wr[121]), .rdlo_out(a2_wr[377]));
			radix2 #(.width(width)) rd_st1_122  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[122]), .rdlo_in(a1_wr[378]),  .coef_in(coef[244]), .rdup_out(a2_wr[122]), .rdlo_out(a2_wr[378]));
			radix2 #(.width(width)) rd_st1_123  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[123]), .rdlo_in(a1_wr[379]),  .coef_in(coef[246]), .rdup_out(a2_wr[123]), .rdlo_out(a2_wr[379]));
			radix2 #(.width(width)) rd_st1_124  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[124]), .rdlo_in(a1_wr[380]),  .coef_in(coef[248]), .rdup_out(a2_wr[124]), .rdlo_out(a2_wr[380]));
			radix2 #(.width(width)) rd_st1_125  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[125]), .rdlo_in(a1_wr[381]),  .coef_in(coef[250]), .rdup_out(a2_wr[125]), .rdlo_out(a2_wr[381]));
			radix2 #(.width(width)) rd_st1_126  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[126]), .rdlo_in(a1_wr[382]),  .coef_in(coef[252]), .rdup_out(a2_wr[126]), .rdlo_out(a2_wr[382]));
			radix2 #(.width(width)) rd_st1_127  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[127]), .rdlo_in(a1_wr[383]),  .coef_in(coef[254]), .rdup_out(a2_wr[127]), .rdlo_out(a2_wr[383]));
			radix2 #(.width(width)) rd_st1_128  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[128]), .rdlo_in(a1_wr[384]),  .coef_in(coef[256]), .rdup_out(a2_wr[128]), .rdlo_out(a2_wr[384]));
			radix2 #(.width(width)) rd_st1_129  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[129]), .rdlo_in(a1_wr[385]),  .coef_in(coef[258]), .rdup_out(a2_wr[129]), .rdlo_out(a2_wr[385]));
			radix2 #(.width(width)) rd_st1_130  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[130]), .rdlo_in(a1_wr[386]),  .coef_in(coef[260]), .rdup_out(a2_wr[130]), .rdlo_out(a2_wr[386]));
			radix2 #(.width(width)) rd_st1_131  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[131]), .rdlo_in(a1_wr[387]),  .coef_in(coef[262]), .rdup_out(a2_wr[131]), .rdlo_out(a2_wr[387]));
			radix2 #(.width(width)) rd_st1_132  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[132]), .rdlo_in(a1_wr[388]),  .coef_in(coef[264]), .rdup_out(a2_wr[132]), .rdlo_out(a2_wr[388]));
			radix2 #(.width(width)) rd_st1_133  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[133]), .rdlo_in(a1_wr[389]),  .coef_in(coef[266]), .rdup_out(a2_wr[133]), .rdlo_out(a2_wr[389]));
			radix2 #(.width(width)) rd_st1_134  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[134]), .rdlo_in(a1_wr[390]),  .coef_in(coef[268]), .rdup_out(a2_wr[134]), .rdlo_out(a2_wr[390]));
			radix2 #(.width(width)) rd_st1_135  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[135]), .rdlo_in(a1_wr[391]),  .coef_in(coef[270]), .rdup_out(a2_wr[135]), .rdlo_out(a2_wr[391]));
			radix2 #(.width(width)) rd_st1_136  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[136]), .rdlo_in(a1_wr[392]),  .coef_in(coef[272]), .rdup_out(a2_wr[136]), .rdlo_out(a2_wr[392]));
			radix2 #(.width(width)) rd_st1_137  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[137]), .rdlo_in(a1_wr[393]),  .coef_in(coef[274]), .rdup_out(a2_wr[137]), .rdlo_out(a2_wr[393]));
			radix2 #(.width(width)) rd_st1_138  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[138]), .rdlo_in(a1_wr[394]),  .coef_in(coef[276]), .rdup_out(a2_wr[138]), .rdlo_out(a2_wr[394]));
			radix2 #(.width(width)) rd_st1_139  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[139]), .rdlo_in(a1_wr[395]),  .coef_in(coef[278]), .rdup_out(a2_wr[139]), .rdlo_out(a2_wr[395]));
			radix2 #(.width(width)) rd_st1_140  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[140]), .rdlo_in(a1_wr[396]),  .coef_in(coef[280]), .rdup_out(a2_wr[140]), .rdlo_out(a2_wr[396]));
			radix2 #(.width(width)) rd_st1_141  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[141]), .rdlo_in(a1_wr[397]),  .coef_in(coef[282]), .rdup_out(a2_wr[141]), .rdlo_out(a2_wr[397]));
			radix2 #(.width(width)) rd_st1_142  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[142]), .rdlo_in(a1_wr[398]),  .coef_in(coef[284]), .rdup_out(a2_wr[142]), .rdlo_out(a2_wr[398]));
			radix2 #(.width(width)) rd_st1_143  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[143]), .rdlo_in(a1_wr[399]),  .coef_in(coef[286]), .rdup_out(a2_wr[143]), .rdlo_out(a2_wr[399]));
			radix2 #(.width(width)) rd_st1_144  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[144]), .rdlo_in(a1_wr[400]),  .coef_in(coef[288]), .rdup_out(a2_wr[144]), .rdlo_out(a2_wr[400]));
			radix2 #(.width(width)) rd_st1_145  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[145]), .rdlo_in(a1_wr[401]),  .coef_in(coef[290]), .rdup_out(a2_wr[145]), .rdlo_out(a2_wr[401]));
			radix2 #(.width(width)) rd_st1_146  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[146]), .rdlo_in(a1_wr[402]),  .coef_in(coef[292]), .rdup_out(a2_wr[146]), .rdlo_out(a2_wr[402]));
			radix2 #(.width(width)) rd_st1_147  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[147]), .rdlo_in(a1_wr[403]),  .coef_in(coef[294]), .rdup_out(a2_wr[147]), .rdlo_out(a2_wr[403]));
			radix2 #(.width(width)) rd_st1_148  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[148]), .rdlo_in(a1_wr[404]),  .coef_in(coef[296]), .rdup_out(a2_wr[148]), .rdlo_out(a2_wr[404]));
			radix2 #(.width(width)) rd_st1_149  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[149]), .rdlo_in(a1_wr[405]),  .coef_in(coef[298]), .rdup_out(a2_wr[149]), .rdlo_out(a2_wr[405]));
			radix2 #(.width(width)) rd_st1_150  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[150]), .rdlo_in(a1_wr[406]),  .coef_in(coef[300]), .rdup_out(a2_wr[150]), .rdlo_out(a2_wr[406]));
			radix2 #(.width(width)) rd_st1_151  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[151]), .rdlo_in(a1_wr[407]),  .coef_in(coef[302]), .rdup_out(a2_wr[151]), .rdlo_out(a2_wr[407]));
			radix2 #(.width(width)) rd_st1_152  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[152]), .rdlo_in(a1_wr[408]),  .coef_in(coef[304]), .rdup_out(a2_wr[152]), .rdlo_out(a2_wr[408]));
			radix2 #(.width(width)) rd_st1_153  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[153]), .rdlo_in(a1_wr[409]),  .coef_in(coef[306]), .rdup_out(a2_wr[153]), .rdlo_out(a2_wr[409]));
			radix2 #(.width(width)) rd_st1_154  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[154]), .rdlo_in(a1_wr[410]),  .coef_in(coef[308]), .rdup_out(a2_wr[154]), .rdlo_out(a2_wr[410]));
			radix2 #(.width(width)) rd_st1_155  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[155]), .rdlo_in(a1_wr[411]),  .coef_in(coef[310]), .rdup_out(a2_wr[155]), .rdlo_out(a2_wr[411]));
			radix2 #(.width(width)) rd_st1_156  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[156]), .rdlo_in(a1_wr[412]),  .coef_in(coef[312]), .rdup_out(a2_wr[156]), .rdlo_out(a2_wr[412]));
			radix2 #(.width(width)) rd_st1_157  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[157]), .rdlo_in(a1_wr[413]),  .coef_in(coef[314]), .rdup_out(a2_wr[157]), .rdlo_out(a2_wr[413]));
			radix2 #(.width(width)) rd_st1_158  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[158]), .rdlo_in(a1_wr[414]),  .coef_in(coef[316]), .rdup_out(a2_wr[158]), .rdlo_out(a2_wr[414]));
			radix2 #(.width(width)) rd_st1_159  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[159]), .rdlo_in(a1_wr[415]),  .coef_in(coef[318]), .rdup_out(a2_wr[159]), .rdlo_out(a2_wr[415]));
			radix2 #(.width(width)) rd_st1_160  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[160]), .rdlo_in(a1_wr[416]),  .coef_in(coef[320]), .rdup_out(a2_wr[160]), .rdlo_out(a2_wr[416]));
			radix2 #(.width(width)) rd_st1_161  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[161]), .rdlo_in(a1_wr[417]),  .coef_in(coef[322]), .rdup_out(a2_wr[161]), .rdlo_out(a2_wr[417]));
			radix2 #(.width(width)) rd_st1_162  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[162]), .rdlo_in(a1_wr[418]),  .coef_in(coef[324]), .rdup_out(a2_wr[162]), .rdlo_out(a2_wr[418]));
			radix2 #(.width(width)) rd_st1_163  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[163]), .rdlo_in(a1_wr[419]),  .coef_in(coef[326]), .rdup_out(a2_wr[163]), .rdlo_out(a2_wr[419]));
			radix2 #(.width(width)) rd_st1_164  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[164]), .rdlo_in(a1_wr[420]),  .coef_in(coef[328]), .rdup_out(a2_wr[164]), .rdlo_out(a2_wr[420]));
			radix2 #(.width(width)) rd_st1_165  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[165]), .rdlo_in(a1_wr[421]),  .coef_in(coef[330]), .rdup_out(a2_wr[165]), .rdlo_out(a2_wr[421]));
			radix2 #(.width(width)) rd_st1_166  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[166]), .rdlo_in(a1_wr[422]),  .coef_in(coef[332]), .rdup_out(a2_wr[166]), .rdlo_out(a2_wr[422]));
			radix2 #(.width(width)) rd_st1_167  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[167]), .rdlo_in(a1_wr[423]),  .coef_in(coef[334]), .rdup_out(a2_wr[167]), .rdlo_out(a2_wr[423]));
			radix2 #(.width(width)) rd_st1_168  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[168]), .rdlo_in(a1_wr[424]),  .coef_in(coef[336]), .rdup_out(a2_wr[168]), .rdlo_out(a2_wr[424]));
			radix2 #(.width(width)) rd_st1_169  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[169]), .rdlo_in(a1_wr[425]),  .coef_in(coef[338]), .rdup_out(a2_wr[169]), .rdlo_out(a2_wr[425]));
			radix2 #(.width(width)) rd_st1_170  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[170]), .rdlo_in(a1_wr[426]),  .coef_in(coef[340]), .rdup_out(a2_wr[170]), .rdlo_out(a2_wr[426]));
			radix2 #(.width(width)) rd_st1_171  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[171]), .rdlo_in(a1_wr[427]),  .coef_in(coef[342]), .rdup_out(a2_wr[171]), .rdlo_out(a2_wr[427]));
			radix2 #(.width(width)) rd_st1_172  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[172]), .rdlo_in(a1_wr[428]),  .coef_in(coef[344]), .rdup_out(a2_wr[172]), .rdlo_out(a2_wr[428]));
			radix2 #(.width(width)) rd_st1_173  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[173]), .rdlo_in(a1_wr[429]),  .coef_in(coef[346]), .rdup_out(a2_wr[173]), .rdlo_out(a2_wr[429]));
			radix2 #(.width(width)) rd_st1_174  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[174]), .rdlo_in(a1_wr[430]),  .coef_in(coef[348]), .rdup_out(a2_wr[174]), .rdlo_out(a2_wr[430]));
			radix2 #(.width(width)) rd_st1_175  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[175]), .rdlo_in(a1_wr[431]),  .coef_in(coef[350]), .rdup_out(a2_wr[175]), .rdlo_out(a2_wr[431]));
			radix2 #(.width(width)) rd_st1_176  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[176]), .rdlo_in(a1_wr[432]),  .coef_in(coef[352]), .rdup_out(a2_wr[176]), .rdlo_out(a2_wr[432]));
			radix2 #(.width(width)) rd_st1_177  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[177]), .rdlo_in(a1_wr[433]),  .coef_in(coef[354]), .rdup_out(a2_wr[177]), .rdlo_out(a2_wr[433]));
			radix2 #(.width(width)) rd_st1_178  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[178]), .rdlo_in(a1_wr[434]),  .coef_in(coef[356]), .rdup_out(a2_wr[178]), .rdlo_out(a2_wr[434]));
			radix2 #(.width(width)) rd_st1_179  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[179]), .rdlo_in(a1_wr[435]),  .coef_in(coef[358]), .rdup_out(a2_wr[179]), .rdlo_out(a2_wr[435]));
			radix2 #(.width(width)) rd_st1_180  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[180]), .rdlo_in(a1_wr[436]),  .coef_in(coef[360]), .rdup_out(a2_wr[180]), .rdlo_out(a2_wr[436]));
			radix2 #(.width(width)) rd_st1_181  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[181]), .rdlo_in(a1_wr[437]),  .coef_in(coef[362]), .rdup_out(a2_wr[181]), .rdlo_out(a2_wr[437]));
			radix2 #(.width(width)) rd_st1_182  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[182]), .rdlo_in(a1_wr[438]),  .coef_in(coef[364]), .rdup_out(a2_wr[182]), .rdlo_out(a2_wr[438]));
			radix2 #(.width(width)) rd_st1_183  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[183]), .rdlo_in(a1_wr[439]),  .coef_in(coef[366]), .rdup_out(a2_wr[183]), .rdlo_out(a2_wr[439]));
			radix2 #(.width(width)) rd_st1_184  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[184]), .rdlo_in(a1_wr[440]),  .coef_in(coef[368]), .rdup_out(a2_wr[184]), .rdlo_out(a2_wr[440]));
			radix2 #(.width(width)) rd_st1_185  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[185]), .rdlo_in(a1_wr[441]),  .coef_in(coef[370]), .rdup_out(a2_wr[185]), .rdlo_out(a2_wr[441]));
			radix2 #(.width(width)) rd_st1_186  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[186]), .rdlo_in(a1_wr[442]),  .coef_in(coef[372]), .rdup_out(a2_wr[186]), .rdlo_out(a2_wr[442]));
			radix2 #(.width(width)) rd_st1_187  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[187]), .rdlo_in(a1_wr[443]),  .coef_in(coef[374]), .rdup_out(a2_wr[187]), .rdlo_out(a2_wr[443]));
			radix2 #(.width(width)) rd_st1_188  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[188]), .rdlo_in(a1_wr[444]),  .coef_in(coef[376]), .rdup_out(a2_wr[188]), .rdlo_out(a2_wr[444]));
			radix2 #(.width(width)) rd_st1_189  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[189]), .rdlo_in(a1_wr[445]),  .coef_in(coef[378]), .rdup_out(a2_wr[189]), .rdlo_out(a2_wr[445]));
			radix2 #(.width(width)) rd_st1_190  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[190]), .rdlo_in(a1_wr[446]),  .coef_in(coef[380]), .rdup_out(a2_wr[190]), .rdlo_out(a2_wr[446]));
			radix2 #(.width(width)) rd_st1_191  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[191]), .rdlo_in(a1_wr[447]),  .coef_in(coef[382]), .rdup_out(a2_wr[191]), .rdlo_out(a2_wr[447]));
			radix2 #(.width(width)) rd_st1_192  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[192]), .rdlo_in(a1_wr[448]),  .coef_in(coef[384]), .rdup_out(a2_wr[192]), .rdlo_out(a2_wr[448]));
			radix2 #(.width(width)) rd_st1_193  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[193]), .rdlo_in(a1_wr[449]),  .coef_in(coef[386]), .rdup_out(a2_wr[193]), .rdlo_out(a2_wr[449]));
			radix2 #(.width(width)) rd_st1_194  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[194]), .rdlo_in(a1_wr[450]),  .coef_in(coef[388]), .rdup_out(a2_wr[194]), .rdlo_out(a2_wr[450]));
			radix2 #(.width(width)) rd_st1_195  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[195]), .rdlo_in(a1_wr[451]),  .coef_in(coef[390]), .rdup_out(a2_wr[195]), .rdlo_out(a2_wr[451]));
			radix2 #(.width(width)) rd_st1_196  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[196]), .rdlo_in(a1_wr[452]),  .coef_in(coef[392]), .rdup_out(a2_wr[196]), .rdlo_out(a2_wr[452]));
			radix2 #(.width(width)) rd_st1_197  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[197]), .rdlo_in(a1_wr[453]),  .coef_in(coef[394]), .rdup_out(a2_wr[197]), .rdlo_out(a2_wr[453]));
			radix2 #(.width(width)) rd_st1_198  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[198]), .rdlo_in(a1_wr[454]),  .coef_in(coef[396]), .rdup_out(a2_wr[198]), .rdlo_out(a2_wr[454]));
			radix2 #(.width(width)) rd_st1_199  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[199]), .rdlo_in(a1_wr[455]),  .coef_in(coef[398]), .rdup_out(a2_wr[199]), .rdlo_out(a2_wr[455]));
			radix2 #(.width(width)) rd_st1_200  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[200]), .rdlo_in(a1_wr[456]),  .coef_in(coef[400]), .rdup_out(a2_wr[200]), .rdlo_out(a2_wr[456]));
			radix2 #(.width(width)) rd_st1_201  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[201]), .rdlo_in(a1_wr[457]),  .coef_in(coef[402]), .rdup_out(a2_wr[201]), .rdlo_out(a2_wr[457]));
			radix2 #(.width(width)) rd_st1_202  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[202]), .rdlo_in(a1_wr[458]),  .coef_in(coef[404]), .rdup_out(a2_wr[202]), .rdlo_out(a2_wr[458]));
			radix2 #(.width(width)) rd_st1_203  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[203]), .rdlo_in(a1_wr[459]),  .coef_in(coef[406]), .rdup_out(a2_wr[203]), .rdlo_out(a2_wr[459]));
			radix2 #(.width(width)) rd_st1_204  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[204]), .rdlo_in(a1_wr[460]),  .coef_in(coef[408]), .rdup_out(a2_wr[204]), .rdlo_out(a2_wr[460]));
			radix2 #(.width(width)) rd_st1_205  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[205]), .rdlo_in(a1_wr[461]),  .coef_in(coef[410]), .rdup_out(a2_wr[205]), .rdlo_out(a2_wr[461]));
			radix2 #(.width(width)) rd_st1_206  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[206]), .rdlo_in(a1_wr[462]),  .coef_in(coef[412]), .rdup_out(a2_wr[206]), .rdlo_out(a2_wr[462]));
			radix2 #(.width(width)) rd_st1_207  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[207]), .rdlo_in(a1_wr[463]),  .coef_in(coef[414]), .rdup_out(a2_wr[207]), .rdlo_out(a2_wr[463]));
			radix2 #(.width(width)) rd_st1_208  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[208]), .rdlo_in(a1_wr[464]),  .coef_in(coef[416]), .rdup_out(a2_wr[208]), .rdlo_out(a2_wr[464]));
			radix2 #(.width(width)) rd_st1_209  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[209]), .rdlo_in(a1_wr[465]),  .coef_in(coef[418]), .rdup_out(a2_wr[209]), .rdlo_out(a2_wr[465]));
			radix2 #(.width(width)) rd_st1_210  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[210]), .rdlo_in(a1_wr[466]),  .coef_in(coef[420]), .rdup_out(a2_wr[210]), .rdlo_out(a2_wr[466]));
			radix2 #(.width(width)) rd_st1_211  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[211]), .rdlo_in(a1_wr[467]),  .coef_in(coef[422]), .rdup_out(a2_wr[211]), .rdlo_out(a2_wr[467]));
			radix2 #(.width(width)) rd_st1_212  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[212]), .rdlo_in(a1_wr[468]),  .coef_in(coef[424]), .rdup_out(a2_wr[212]), .rdlo_out(a2_wr[468]));
			radix2 #(.width(width)) rd_st1_213  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[213]), .rdlo_in(a1_wr[469]),  .coef_in(coef[426]), .rdup_out(a2_wr[213]), .rdlo_out(a2_wr[469]));
			radix2 #(.width(width)) rd_st1_214  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[214]), .rdlo_in(a1_wr[470]),  .coef_in(coef[428]), .rdup_out(a2_wr[214]), .rdlo_out(a2_wr[470]));
			radix2 #(.width(width)) rd_st1_215  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[215]), .rdlo_in(a1_wr[471]),  .coef_in(coef[430]), .rdup_out(a2_wr[215]), .rdlo_out(a2_wr[471]));
			radix2 #(.width(width)) rd_st1_216  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[216]), .rdlo_in(a1_wr[472]),  .coef_in(coef[432]), .rdup_out(a2_wr[216]), .rdlo_out(a2_wr[472]));
			radix2 #(.width(width)) rd_st1_217  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[217]), .rdlo_in(a1_wr[473]),  .coef_in(coef[434]), .rdup_out(a2_wr[217]), .rdlo_out(a2_wr[473]));
			radix2 #(.width(width)) rd_st1_218  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[218]), .rdlo_in(a1_wr[474]),  .coef_in(coef[436]), .rdup_out(a2_wr[218]), .rdlo_out(a2_wr[474]));
			radix2 #(.width(width)) rd_st1_219  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[219]), .rdlo_in(a1_wr[475]),  .coef_in(coef[438]), .rdup_out(a2_wr[219]), .rdlo_out(a2_wr[475]));
			radix2 #(.width(width)) rd_st1_220  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[220]), .rdlo_in(a1_wr[476]),  .coef_in(coef[440]), .rdup_out(a2_wr[220]), .rdlo_out(a2_wr[476]));
			radix2 #(.width(width)) rd_st1_221  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[221]), .rdlo_in(a1_wr[477]),  .coef_in(coef[442]), .rdup_out(a2_wr[221]), .rdlo_out(a2_wr[477]));
			radix2 #(.width(width)) rd_st1_222  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[222]), .rdlo_in(a1_wr[478]),  .coef_in(coef[444]), .rdup_out(a2_wr[222]), .rdlo_out(a2_wr[478]));
			radix2 #(.width(width)) rd_st1_223  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[223]), .rdlo_in(a1_wr[479]),  .coef_in(coef[446]), .rdup_out(a2_wr[223]), .rdlo_out(a2_wr[479]));
			radix2 #(.width(width)) rd_st1_224  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[224]), .rdlo_in(a1_wr[480]),  .coef_in(coef[448]), .rdup_out(a2_wr[224]), .rdlo_out(a2_wr[480]));
			radix2 #(.width(width)) rd_st1_225  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[225]), .rdlo_in(a1_wr[481]),  .coef_in(coef[450]), .rdup_out(a2_wr[225]), .rdlo_out(a2_wr[481]));
			radix2 #(.width(width)) rd_st1_226  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[226]), .rdlo_in(a1_wr[482]),  .coef_in(coef[452]), .rdup_out(a2_wr[226]), .rdlo_out(a2_wr[482]));
			radix2 #(.width(width)) rd_st1_227  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[227]), .rdlo_in(a1_wr[483]),  .coef_in(coef[454]), .rdup_out(a2_wr[227]), .rdlo_out(a2_wr[483]));
			radix2 #(.width(width)) rd_st1_228  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[228]), .rdlo_in(a1_wr[484]),  .coef_in(coef[456]), .rdup_out(a2_wr[228]), .rdlo_out(a2_wr[484]));
			radix2 #(.width(width)) rd_st1_229  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[229]), .rdlo_in(a1_wr[485]),  .coef_in(coef[458]), .rdup_out(a2_wr[229]), .rdlo_out(a2_wr[485]));
			radix2 #(.width(width)) rd_st1_230  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[230]), .rdlo_in(a1_wr[486]),  .coef_in(coef[460]), .rdup_out(a2_wr[230]), .rdlo_out(a2_wr[486]));
			radix2 #(.width(width)) rd_st1_231  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[231]), .rdlo_in(a1_wr[487]),  .coef_in(coef[462]), .rdup_out(a2_wr[231]), .rdlo_out(a2_wr[487]));
			radix2 #(.width(width)) rd_st1_232  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[232]), .rdlo_in(a1_wr[488]),  .coef_in(coef[464]), .rdup_out(a2_wr[232]), .rdlo_out(a2_wr[488]));
			radix2 #(.width(width)) rd_st1_233  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[233]), .rdlo_in(a1_wr[489]),  .coef_in(coef[466]), .rdup_out(a2_wr[233]), .rdlo_out(a2_wr[489]));
			radix2 #(.width(width)) rd_st1_234  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[234]), .rdlo_in(a1_wr[490]),  .coef_in(coef[468]), .rdup_out(a2_wr[234]), .rdlo_out(a2_wr[490]));
			radix2 #(.width(width)) rd_st1_235  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[235]), .rdlo_in(a1_wr[491]),  .coef_in(coef[470]), .rdup_out(a2_wr[235]), .rdlo_out(a2_wr[491]));
			radix2 #(.width(width)) rd_st1_236  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[236]), .rdlo_in(a1_wr[492]),  .coef_in(coef[472]), .rdup_out(a2_wr[236]), .rdlo_out(a2_wr[492]));
			radix2 #(.width(width)) rd_st1_237  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[237]), .rdlo_in(a1_wr[493]),  .coef_in(coef[474]), .rdup_out(a2_wr[237]), .rdlo_out(a2_wr[493]));
			radix2 #(.width(width)) rd_st1_238  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[238]), .rdlo_in(a1_wr[494]),  .coef_in(coef[476]), .rdup_out(a2_wr[238]), .rdlo_out(a2_wr[494]));
			radix2 #(.width(width)) rd_st1_239  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[239]), .rdlo_in(a1_wr[495]),  .coef_in(coef[478]), .rdup_out(a2_wr[239]), .rdlo_out(a2_wr[495]));
			radix2 #(.width(width)) rd_st1_240  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[240]), .rdlo_in(a1_wr[496]),  .coef_in(coef[480]), .rdup_out(a2_wr[240]), .rdlo_out(a2_wr[496]));
			radix2 #(.width(width)) rd_st1_241  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[241]), .rdlo_in(a1_wr[497]),  .coef_in(coef[482]), .rdup_out(a2_wr[241]), .rdlo_out(a2_wr[497]));
			radix2 #(.width(width)) rd_st1_242  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[242]), .rdlo_in(a1_wr[498]),  .coef_in(coef[484]), .rdup_out(a2_wr[242]), .rdlo_out(a2_wr[498]));
			radix2 #(.width(width)) rd_st1_243  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[243]), .rdlo_in(a1_wr[499]),  .coef_in(coef[486]), .rdup_out(a2_wr[243]), .rdlo_out(a2_wr[499]));
			radix2 #(.width(width)) rd_st1_244  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[244]), .rdlo_in(a1_wr[500]),  .coef_in(coef[488]), .rdup_out(a2_wr[244]), .rdlo_out(a2_wr[500]));
			radix2 #(.width(width)) rd_st1_245  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[245]), .rdlo_in(a1_wr[501]),  .coef_in(coef[490]), .rdup_out(a2_wr[245]), .rdlo_out(a2_wr[501]));
			radix2 #(.width(width)) rd_st1_246  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[246]), .rdlo_in(a1_wr[502]),  .coef_in(coef[492]), .rdup_out(a2_wr[246]), .rdlo_out(a2_wr[502]));
			radix2 #(.width(width)) rd_st1_247  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[247]), .rdlo_in(a1_wr[503]),  .coef_in(coef[494]), .rdup_out(a2_wr[247]), .rdlo_out(a2_wr[503]));
			radix2 #(.width(width)) rd_st1_248  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[248]), .rdlo_in(a1_wr[504]),  .coef_in(coef[496]), .rdup_out(a2_wr[248]), .rdlo_out(a2_wr[504]));
			radix2 #(.width(width)) rd_st1_249  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[249]), .rdlo_in(a1_wr[505]),  .coef_in(coef[498]), .rdup_out(a2_wr[249]), .rdlo_out(a2_wr[505]));
			radix2 #(.width(width)) rd_st1_250  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[250]), .rdlo_in(a1_wr[506]),  .coef_in(coef[500]), .rdup_out(a2_wr[250]), .rdlo_out(a2_wr[506]));
			radix2 #(.width(width)) rd_st1_251  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[251]), .rdlo_in(a1_wr[507]),  .coef_in(coef[502]), .rdup_out(a2_wr[251]), .rdlo_out(a2_wr[507]));
			radix2 #(.width(width)) rd_st1_252  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[252]), .rdlo_in(a1_wr[508]),  .coef_in(coef[504]), .rdup_out(a2_wr[252]), .rdlo_out(a2_wr[508]));
			radix2 #(.width(width)) rd_st1_253  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[253]), .rdlo_in(a1_wr[509]),  .coef_in(coef[506]), .rdup_out(a2_wr[253]), .rdlo_out(a2_wr[509]));
			radix2 #(.width(width)) rd_st1_254  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[254]), .rdlo_in(a1_wr[510]),  .coef_in(coef[508]), .rdup_out(a2_wr[254]), .rdlo_out(a2_wr[510]));
			radix2 #(.width(width)) rd_st1_255  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[255]), .rdlo_in(a1_wr[511]),  .coef_in(coef[510]), .rdup_out(a2_wr[255]), .rdlo_out(a2_wr[511]));
			radix2 #(.width(width)) rd_st1_512  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[512]), .rdlo_in(a1_wr[768]),  .coef_in(coef[0]), .rdup_out(a2_wr[512]), .rdlo_out(a2_wr[768]));
			radix2 #(.width(width)) rd_st1_513  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[513]), .rdlo_in(a1_wr[769]),  .coef_in(coef[2]), .rdup_out(a2_wr[513]), .rdlo_out(a2_wr[769]));
			radix2 #(.width(width)) rd_st1_514  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[514]), .rdlo_in(a1_wr[770]),  .coef_in(coef[4]), .rdup_out(a2_wr[514]), .rdlo_out(a2_wr[770]));
			radix2 #(.width(width)) rd_st1_515  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[515]), .rdlo_in(a1_wr[771]),  .coef_in(coef[6]), .rdup_out(a2_wr[515]), .rdlo_out(a2_wr[771]));
			radix2 #(.width(width)) rd_st1_516  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[516]), .rdlo_in(a1_wr[772]),  .coef_in(coef[8]), .rdup_out(a2_wr[516]), .rdlo_out(a2_wr[772]));
			radix2 #(.width(width)) rd_st1_517  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[517]), .rdlo_in(a1_wr[773]),  .coef_in(coef[10]), .rdup_out(a2_wr[517]), .rdlo_out(a2_wr[773]));
			radix2 #(.width(width)) rd_st1_518  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[518]), .rdlo_in(a1_wr[774]),  .coef_in(coef[12]), .rdup_out(a2_wr[518]), .rdlo_out(a2_wr[774]));
			radix2 #(.width(width)) rd_st1_519  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[519]), .rdlo_in(a1_wr[775]),  .coef_in(coef[14]), .rdup_out(a2_wr[519]), .rdlo_out(a2_wr[775]));
			radix2 #(.width(width)) rd_st1_520  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[520]), .rdlo_in(a1_wr[776]),  .coef_in(coef[16]), .rdup_out(a2_wr[520]), .rdlo_out(a2_wr[776]));
			radix2 #(.width(width)) rd_st1_521  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[521]), .rdlo_in(a1_wr[777]),  .coef_in(coef[18]), .rdup_out(a2_wr[521]), .rdlo_out(a2_wr[777]));
			radix2 #(.width(width)) rd_st1_522  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[522]), .rdlo_in(a1_wr[778]),  .coef_in(coef[20]), .rdup_out(a2_wr[522]), .rdlo_out(a2_wr[778]));
			radix2 #(.width(width)) rd_st1_523  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[523]), .rdlo_in(a1_wr[779]),  .coef_in(coef[22]), .rdup_out(a2_wr[523]), .rdlo_out(a2_wr[779]));
			radix2 #(.width(width)) rd_st1_524  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[524]), .rdlo_in(a1_wr[780]),  .coef_in(coef[24]), .rdup_out(a2_wr[524]), .rdlo_out(a2_wr[780]));
			radix2 #(.width(width)) rd_st1_525  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[525]), .rdlo_in(a1_wr[781]),  .coef_in(coef[26]), .rdup_out(a2_wr[525]), .rdlo_out(a2_wr[781]));
			radix2 #(.width(width)) rd_st1_526  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[526]), .rdlo_in(a1_wr[782]),  .coef_in(coef[28]), .rdup_out(a2_wr[526]), .rdlo_out(a2_wr[782]));
			radix2 #(.width(width)) rd_st1_527  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[527]), .rdlo_in(a1_wr[783]),  .coef_in(coef[30]), .rdup_out(a2_wr[527]), .rdlo_out(a2_wr[783]));
			radix2 #(.width(width)) rd_st1_528  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[528]), .rdlo_in(a1_wr[784]),  .coef_in(coef[32]), .rdup_out(a2_wr[528]), .rdlo_out(a2_wr[784]));
			radix2 #(.width(width)) rd_st1_529  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[529]), .rdlo_in(a1_wr[785]),  .coef_in(coef[34]), .rdup_out(a2_wr[529]), .rdlo_out(a2_wr[785]));
			radix2 #(.width(width)) rd_st1_530  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[530]), .rdlo_in(a1_wr[786]),  .coef_in(coef[36]), .rdup_out(a2_wr[530]), .rdlo_out(a2_wr[786]));
			radix2 #(.width(width)) rd_st1_531  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[531]), .rdlo_in(a1_wr[787]),  .coef_in(coef[38]), .rdup_out(a2_wr[531]), .rdlo_out(a2_wr[787]));
			radix2 #(.width(width)) rd_st1_532  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[532]), .rdlo_in(a1_wr[788]),  .coef_in(coef[40]), .rdup_out(a2_wr[532]), .rdlo_out(a2_wr[788]));
			radix2 #(.width(width)) rd_st1_533  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[533]), .rdlo_in(a1_wr[789]),  .coef_in(coef[42]), .rdup_out(a2_wr[533]), .rdlo_out(a2_wr[789]));
			radix2 #(.width(width)) rd_st1_534  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[534]), .rdlo_in(a1_wr[790]),  .coef_in(coef[44]), .rdup_out(a2_wr[534]), .rdlo_out(a2_wr[790]));
			radix2 #(.width(width)) rd_st1_535  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[535]), .rdlo_in(a1_wr[791]),  .coef_in(coef[46]), .rdup_out(a2_wr[535]), .rdlo_out(a2_wr[791]));
			radix2 #(.width(width)) rd_st1_536  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[536]), .rdlo_in(a1_wr[792]),  .coef_in(coef[48]), .rdup_out(a2_wr[536]), .rdlo_out(a2_wr[792]));
			radix2 #(.width(width)) rd_st1_537  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[537]), .rdlo_in(a1_wr[793]),  .coef_in(coef[50]), .rdup_out(a2_wr[537]), .rdlo_out(a2_wr[793]));
			radix2 #(.width(width)) rd_st1_538  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[538]), .rdlo_in(a1_wr[794]),  .coef_in(coef[52]), .rdup_out(a2_wr[538]), .rdlo_out(a2_wr[794]));
			radix2 #(.width(width)) rd_st1_539  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[539]), .rdlo_in(a1_wr[795]),  .coef_in(coef[54]), .rdup_out(a2_wr[539]), .rdlo_out(a2_wr[795]));
			radix2 #(.width(width)) rd_st1_540  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[540]), .rdlo_in(a1_wr[796]),  .coef_in(coef[56]), .rdup_out(a2_wr[540]), .rdlo_out(a2_wr[796]));
			radix2 #(.width(width)) rd_st1_541  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[541]), .rdlo_in(a1_wr[797]),  .coef_in(coef[58]), .rdup_out(a2_wr[541]), .rdlo_out(a2_wr[797]));
			radix2 #(.width(width)) rd_st1_542  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[542]), .rdlo_in(a1_wr[798]),  .coef_in(coef[60]), .rdup_out(a2_wr[542]), .rdlo_out(a2_wr[798]));
			radix2 #(.width(width)) rd_st1_543  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[543]), .rdlo_in(a1_wr[799]),  .coef_in(coef[62]), .rdup_out(a2_wr[543]), .rdlo_out(a2_wr[799]));
			radix2 #(.width(width)) rd_st1_544  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[544]), .rdlo_in(a1_wr[800]),  .coef_in(coef[64]), .rdup_out(a2_wr[544]), .rdlo_out(a2_wr[800]));
			radix2 #(.width(width)) rd_st1_545  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[545]), .rdlo_in(a1_wr[801]),  .coef_in(coef[66]), .rdup_out(a2_wr[545]), .rdlo_out(a2_wr[801]));
			radix2 #(.width(width)) rd_st1_546  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[546]), .rdlo_in(a1_wr[802]),  .coef_in(coef[68]), .rdup_out(a2_wr[546]), .rdlo_out(a2_wr[802]));
			radix2 #(.width(width)) rd_st1_547  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[547]), .rdlo_in(a1_wr[803]),  .coef_in(coef[70]), .rdup_out(a2_wr[547]), .rdlo_out(a2_wr[803]));
			radix2 #(.width(width)) rd_st1_548  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[548]), .rdlo_in(a1_wr[804]),  .coef_in(coef[72]), .rdup_out(a2_wr[548]), .rdlo_out(a2_wr[804]));
			radix2 #(.width(width)) rd_st1_549  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[549]), .rdlo_in(a1_wr[805]),  .coef_in(coef[74]), .rdup_out(a2_wr[549]), .rdlo_out(a2_wr[805]));
			radix2 #(.width(width)) rd_st1_550  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[550]), .rdlo_in(a1_wr[806]),  .coef_in(coef[76]), .rdup_out(a2_wr[550]), .rdlo_out(a2_wr[806]));
			radix2 #(.width(width)) rd_st1_551  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[551]), .rdlo_in(a1_wr[807]),  .coef_in(coef[78]), .rdup_out(a2_wr[551]), .rdlo_out(a2_wr[807]));
			radix2 #(.width(width)) rd_st1_552  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[552]), .rdlo_in(a1_wr[808]),  .coef_in(coef[80]), .rdup_out(a2_wr[552]), .rdlo_out(a2_wr[808]));
			radix2 #(.width(width)) rd_st1_553  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[553]), .rdlo_in(a1_wr[809]),  .coef_in(coef[82]), .rdup_out(a2_wr[553]), .rdlo_out(a2_wr[809]));
			radix2 #(.width(width)) rd_st1_554  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[554]), .rdlo_in(a1_wr[810]),  .coef_in(coef[84]), .rdup_out(a2_wr[554]), .rdlo_out(a2_wr[810]));
			radix2 #(.width(width)) rd_st1_555  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[555]), .rdlo_in(a1_wr[811]),  .coef_in(coef[86]), .rdup_out(a2_wr[555]), .rdlo_out(a2_wr[811]));
			radix2 #(.width(width)) rd_st1_556  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[556]), .rdlo_in(a1_wr[812]),  .coef_in(coef[88]), .rdup_out(a2_wr[556]), .rdlo_out(a2_wr[812]));
			radix2 #(.width(width)) rd_st1_557  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[557]), .rdlo_in(a1_wr[813]),  .coef_in(coef[90]), .rdup_out(a2_wr[557]), .rdlo_out(a2_wr[813]));
			radix2 #(.width(width)) rd_st1_558  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[558]), .rdlo_in(a1_wr[814]),  .coef_in(coef[92]), .rdup_out(a2_wr[558]), .rdlo_out(a2_wr[814]));
			radix2 #(.width(width)) rd_st1_559  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[559]), .rdlo_in(a1_wr[815]),  .coef_in(coef[94]), .rdup_out(a2_wr[559]), .rdlo_out(a2_wr[815]));
			radix2 #(.width(width)) rd_st1_560  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[560]), .rdlo_in(a1_wr[816]),  .coef_in(coef[96]), .rdup_out(a2_wr[560]), .rdlo_out(a2_wr[816]));
			radix2 #(.width(width)) rd_st1_561  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[561]), .rdlo_in(a1_wr[817]),  .coef_in(coef[98]), .rdup_out(a2_wr[561]), .rdlo_out(a2_wr[817]));
			radix2 #(.width(width)) rd_st1_562  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[562]), .rdlo_in(a1_wr[818]),  .coef_in(coef[100]), .rdup_out(a2_wr[562]), .rdlo_out(a2_wr[818]));
			radix2 #(.width(width)) rd_st1_563  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[563]), .rdlo_in(a1_wr[819]),  .coef_in(coef[102]), .rdup_out(a2_wr[563]), .rdlo_out(a2_wr[819]));
			radix2 #(.width(width)) rd_st1_564  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[564]), .rdlo_in(a1_wr[820]),  .coef_in(coef[104]), .rdup_out(a2_wr[564]), .rdlo_out(a2_wr[820]));
			radix2 #(.width(width)) rd_st1_565  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[565]), .rdlo_in(a1_wr[821]),  .coef_in(coef[106]), .rdup_out(a2_wr[565]), .rdlo_out(a2_wr[821]));
			radix2 #(.width(width)) rd_st1_566  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[566]), .rdlo_in(a1_wr[822]),  .coef_in(coef[108]), .rdup_out(a2_wr[566]), .rdlo_out(a2_wr[822]));
			radix2 #(.width(width)) rd_st1_567  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[567]), .rdlo_in(a1_wr[823]),  .coef_in(coef[110]), .rdup_out(a2_wr[567]), .rdlo_out(a2_wr[823]));
			radix2 #(.width(width)) rd_st1_568  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[568]), .rdlo_in(a1_wr[824]),  .coef_in(coef[112]), .rdup_out(a2_wr[568]), .rdlo_out(a2_wr[824]));
			radix2 #(.width(width)) rd_st1_569  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[569]), .rdlo_in(a1_wr[825]),  .coef_in(coef[114]), .rdup_out(a2_wr[569]), .rdlo_out(a2_wr[825]));
			radix2 #(.width(width)) rd_st1_570  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[570]), .rdlo_in(a1_wr[826]),  .coef_in(coef[116]), .rdup_out(a2_wr[570]), .rdlo_out(a2_wr[826]));
			radix2 #(.width(width)) rd_st1_571  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[571]), .rdlo_in(a1_wr[827]),  .coef_in(coef[118]), .rdup_out(a2_wr[571]), .rdlo_out(a2_wr[827]));
			radix2 #(.width(width)) rd_st1_572  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[572]), .rdlo_in(a1_wr[828]),  .coef_in(coef[120]), .rdup_out(a2_wr[572]), .rdlo_out(a2_wr[828]));
			radix2 #(.width(width)) rd_st1_573  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[573]), .rdlo_in(a1_wr[829]),  .coef_in(coef[122]), .rdup_out(a2_wr[573]), .rdlo_out(a2_wr[829]));
			radix2 #(.width(width)) rd_st1_574  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[574]), .rdlo_in(a1_wr[830]),  .coef_in(coef[124]), .rdup_out(a2_wr[574]), .rdlo_out(a2_wr[830]));
			radix2 #(.width(width)) rd_st1_575  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[575]), .rdlo_in(a1_wr[831]),  .coef_in(coef[126]), .rdup_out(a2_wr[575]), .rdlo_out(a2_wr[831]));
			radix2 #(.width(width)) rd_st1_576  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[576]), .rdlo_in(a1_wr[832]),  .coef_in(coef[128]), .rdup_out(a2_wr[576]), .rdlo_out(a2_wr[832]));
			radix2 #(.width(width)) rd_st1_577  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[577]), .rdlo_in(a1_wr[833]),  .coef_in(coef[130]), .rdup_out(a2_wr[577]), .rdlo_out(a2_wr[833]));
			radix2 #(.width(width)) rd_st1_578  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[578]), .rdlo_in(a1_wr[834]),  .coef_in(coef[132]), .rdup_out(a2_wr[578]), .rdlo_out(a2_wr[834]));
			radix2 #(.width(width)) rd_st1_579  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[579]), .rdlo_in(a1_wr[835]),  .coef_in(coef[134]), .rdup_out(a2_wr[579]), .rdlo_out(a2_wr[835]));
			radix2 #(.width(width)) rd_st1_580  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[580]), .rdlo_in(a1_wr[836]),  .coef_in(coef[136]), .rdup_out(a2_wr[580]), .rdlo_out(a2_wr[836]));
			radix2 #(.width(width)) rd_st1_581  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[581]), .rdlo_in(a1_wr[837]),  .coef_in(coef[138]), .rdup_out(a2_wr[581]), .rdlo_out(a2_wr[837]));
			radix2 #(.width(width)) rd_st1_582  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[582]), .rdlo_in(a1_wr[838]),  .coef_in(coef[140]), .rdup_out(a2_wr[582]), .rdlo_out(a2_wr[838]));
			radix2 #(.width(width)) rd_st1_583  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[583]), .rdlo_in(a1_wr[839]),  .coef_in(coef[142]), .rdup_out(a2_wr[583]), .rdlo_out(a2_wr[839]));
			radix2 #(.width(width)) rd_st1_584  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[584]), .rdlo_in(a1_wr[840]),  .coef_in(coef[144]), .rdup_out(a2_wr[584]), .rdlo_out(a2_wr[840]));
			radix2 #(.width(width)) rd_st1_585  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[585]), .rdlo_in(a1_wr[841]),  .coef_in(coef[146]), .rdup_out(a2_wr[585]), .rdlo_out(a2_wr[841]));
			radix2 #(.width(width)) rd_st1_586  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[586]), .rdlo_in(a1_wr[842]),  .coef_in(coef[148]), .rdup_out(a2_wr[586]), .rdlo_out(a2_wr[842]));
			radix2 #(.width(width)) rd_st1_587  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[587]), .rdlo_in(a1_wr[843]),  .coef_in(coef[150]), .rdup_out(a2_wr[587]), .rdlo_out(a2_wr[843]));
			radix2 #(.width(width)) rd_st1_588  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[588]), .rdlo_in(a1_wr[844]),  .coef_in(coef[152]), .rdup_out(a2_wr[588]), .rdlo_out(a2_wr[844]));
			radix2 #(.width(width)) rd_st1_589  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[589]), .rdlo_in(a1_wr[845]),  .coef_in(coef[154]), .rdup_out(a2_wr[589]), .rdlo_out(a2_wr[845]));
			radix2 #(.width(width)) rd_st1_590  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[590]), .rdlo_in(a1_wr[846]),  .coef_in(coef[156]), .rdup_out(a2_wr[590]), .rdlo_out(a2_wr[846]));
			radix2 #(.width(width)) rd_st1_591  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[591]), .rdlo_in(a1_wr[847]),  .coef_in(coef[158]), .rdup_out(a2_wr[591]), .rdlo_out(a2_wr[847]));
			radix2 #(.width(width)) rd_st1_592  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[592]), .rdlo_in(a1_wr[848]),  .coef_in(coef[160]), .rdup_out(a2_wr[592]), .rdlo_out(a2_wr[848]));
			radix2 #(.width(width)) rd_st1_593  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[593]), .rdlo_in(a1_wr[849]),  .coef_in(coef[162]), .rdup_out(a2_wr[593]), .rdlo_out(a2_wr[849]));
			radix2 #(.width(width)) rd_st1_594  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[594]), .rdlo_in(a1_wr[850]),  .coef_in(coef[164]), .rdup_out(a2_wr[594]), .rdlo_out(a2_wr[850]));
			radix2 #(.width(width)) rd_st1_595  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[595]), .rdlo_in(a1_wr[851]),  .coef_in(coef[166]), .rdup_out(a2_wr[595]), .rdlo_out(a2_wr[851]));
			radix2 #(.width(width)) rd_st1_596  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[596]), .rdlo_in(a1_wr[852]),  .coef_in(coef[168]), .rdup_out(a2_wr[596]), .rdlo_out(a2_wr[852]));
			radix2 #(.width(width)) rd_st1_597  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[597]), .rdlo_in(a1_wr[853]),  .coef_in(coef[170]), .rdup_out(a2_wr[597]), .rdlo_out(a2_wr[853]));
			radix2 #(.width(width)) rd_st1_598  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[598]), .rdlo_in(a1_wr[854]),  .coef_in(coef[172]), .rdup_out(a2_wr[598]), .rdlo_out(a2_wr[854]));
			radix2 #(.width(width)) rd_st1_599  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[599]), .rdlo_in(a1_wr[855]),  .coef_in(coef[174]), .rdup_out(a2_wr[599]), .rdlo_out(a2_wr[855]));
			radix2 #(.width(width)) rd_st1_600  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[600]), .rdlo_in(a1_wr[856]),  .coef_in(coef[176]), .rdup_out(a2_wr[600]), .rdlo_out(a2_wr[856]));
			radix2 #(.width(width)) rd_st1_601  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[601]), .rdlo_in(a1_wr[857]),  .coef_in(coef[178]), .rdup_out(a2_wr[601]), .rdlo_out(a2_wr[857]));
			radix2 #(.width(width)) rd_st1_602  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[602]), .rdlo_in(a1_wr[858]),  .coef_in(coef[180]), .rdup_out(a2_wr[602]), .rdlo_out(a2_wr[858]));
			radix2 #(.width(width)) rd_st1_603  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[603]), .rdlo_in(a1_wr[859]),  .coef_in(coef[182]), .rdup_out(a2_wr[603]), .rdlo_out(a2_wr[859]));
			radix2 #(.width(width)) rd_st1_604  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[604]), .rdlo_in(a1_wr[860]),  .coef_in(coef[184]), .rdup_out(a2_wr[604]), .rdlo_out(a2_wr[860]));
			radix2 #(.width(width)) rd_st1_605  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[605]), .rdlo_in(a1_wr[861]),  .coef_in(coef[186]), .rdup_out(a2_wr[605]), .rdlo_out(a2_wr[861]));
			radix2 #(.width(width)) rd_st1_606  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[606]), .rdlo_in(a1_wr[862]),  .coef_in(coef[188]), .rdup_out(a2_wr[606]), .rdlo_out(a2_wr[862]));
			radix2 #(.width(width)) rd_st1_607  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[607]), .rdlo_in(a1_wr[863]),  .coef_in(coef[190]), .rdup_out(a2_wr[607]), .rdlo_out(a2_wr[863]));
			radix2 #(.width(width)) rd_st1_608  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[608]), .rdlo_in(a1_wr[864]),  .coef_in(coef[192]), .rdup_out(a2_wr[608]), .rdlo_out(a2_wr[864]));
			radix2 #(.width(width)) rd_st1_609  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[609]), .rdlo_in(a1_wr[865]),  .coef_in(coef[194]), .rdup_out(a2_wr[609]), .rdlo_out(a2_wr[865]));
			radix2 #(.width(width)) rd_st1_610  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[610]), .rdlo_in(a1_wr[866]),  .coef_in(coef[196]), .rdup_out(a2_wr[610]), .rdlo_out(a2_wr[866]));
			radix2 #(.width(width)) rd_st1_611  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[611]), .rdlo_in(a1_wr[867]),  .coef_in(coef[198]), .rdup_out(a2_wr[611]), .rdlo_out(a2_wr[867]));
			radix2 #(.width(width)) rd_st1_612  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[612]), .rdlo_in(a1_wr[868]),  .coef_in(coef[200]), .rdup_out(a2_wr[612]), .rdlo_out(a2_wr[868]));
			radix2 #(.width(width)) rd_st1_613  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[613]), .rdlo_in(a1_wr[869]),  .coef_in(coef[202]), .rdup_out(a2_wr[613]), .rdlo_out(a2_wr[869]));
			radix2 #(.width(width)) rd_st1_614  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[614]), .rdlo_in(a1_wr[870]),  .coef_in(coef[204]), .rdup_out(a2_wr[614]), .rdlo_out(a2_wr[870]));
			radix2 #(.width(width)) rd_st1_615  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[615]), .rdlo_in(a1_wr[871]),  .coef_in(coef[206]), .rdup_out(a2_wr[615]), .rdlo_out(a2_wr[871]));
			radix2 #(.width(width)) rd_st1_616  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[616]), .rdlo_in(a1_wr[872]),  .coef_in(coef[208]), .rdup_out(a2_wr[616]), .rdlo_out(a2_wr[872]));
			radix2 #(.width(width)) rd_st1_617  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[617]), .rdlo_in(a1_wr[873]),  .coef_in(coef[210]), .rdup_out(a2_wr[617]), .rdlo_out(a2_wr[873]));
			radix2 #(.width(width)) rd_st1_618  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[618]), .rdlo_in(a1_wr[874]),  .coef_in(coef[212]), .rdup_out(a2_wr[618]), .rdlo_out(a2_wr[874]));
			radix2 #(.width(width)) rd_st1_619  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[619]), .rdlo_in(a1_wr[875]),  .coef_in(coef[214]), .rdup_out(a2_wr[619]), .rdlo_out(a2_wr[875]));
			radix2 #(.width(width)) rd_st1_620  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[620]), .rdlo_in(a1_wr[876]),  .coef_in(coef[216]), .rdup_out(a2_wr[620]), .rdlo_out(a2_wr[876]));
			radix2 #(.width(width)) rd_st1_621  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[621]), .rdlo_in(a1_wr[877]),  .coef_in(coef[218]), .rdup_out(a2_wr[621]), .rdlo_out(a2_wr[877]));
			radix2 #(.width(width)) rd_st1_622  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[622]), .rdlo_in(a1_wr[878]),  .coef_in(coef[220]), .rdup_out(a2_wr[622]), .rdlo_out(a2_wr[878]));
			radix2 #(.width(width)) rd_st1_623  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[623]), .rdlo_in(a1_wr[879]),  .coef_in(coef[222]), .rdup_out(a2_wr[623]), .rdlo_out(a2_wr[879]));
			radix2 #(.width(width)) rd_st1_624  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[624]), .rdlo_in(a1_wr[880]),  .coef_in(coef[224]), .rdup_out(a2_wr[624]), .rdlo_out(a2_wr[880]));
			radix2 #(.width(width)) rd_st1_625  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[625]), .rdlo_in(a1_wr[881]),  .coef_in(coef[226]), .rdup_out(a2_wr[625]), .rdlo_out(a2_wr[881]));
			radix2 #(.width(width)) rd_st1_626  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[626]), .rdlo_in(a1_wr[882]),  .coef_in(coef[228]), .rdup_out(a2_wr[626]), .rdlo_out(a2_wr[882]));
			radix2 #(.width(width)) rd_st1_627  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[627]), .rdlo_in(a1_wr[883]),  .coef_in(coef[230]), .rdup_out(a2_wr[627]), .rdlo_out(a2_wr[883]));
			radix2 #(.width(width)) rd_st1_628  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[628]), .rdlo_in(a1_wr[884]),  .coef_in(coef[232]), .rdup_out(a2_wr[628]), .rdlo_out(a2_wr[884]));
			radix2 #(.width(width)) rd_st1_629  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[629]), .rdlo_in(a1_wr[885]),  .coef_in(coef[234]), .rdup_out(a2_wr[629]), .rdlo_out(a2_wr[885]));
			radix2 #(.width(width)) rd_st1_630  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[630]), .rdlo_in(a1_wr[886]),  .coef_in(coef[236]), .rdup_out(a2_wr[630]), .rdlo_out(a2_wr[886]));
			radix2 #(.width(width)) rd_st1_631  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[631]), .rdlo_in(a1_wr[887]),  .coef_in(coef[238]), .rdup_out(a2_wr[631]), .rdlo_out(a2_wr[887]));
			radix2 #(.width(width)) rd_st1_632  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[632]), .rdlo_in(a1_wr[888]),  .coef_in(coef[240]), .rdup_out(a2_wr[632]), .rdlo_out(a2_wr[888]));
			radix2 #(.width(width)) rd_st1_633  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[633]), .rdlo_in(a1_wr[889]),  .coef_in(coef[242]), .rdup_out(a2_wr[633]), .rdlo_out(a2_wr[889]));
			radix2 #(.width(width)) rd_st1_634  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[634]), .rdlo_in(a1_wr[890]),  .coef_in(coef[244]), .rdup_out(a2_wr[634]), .rdlo_out(a2_wr[890]));
			radix2 #(.width(width)) rd_st1_635  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[635]), .rdlo_in(a1_wr[891]),  .coef_in(coef[246]), .rdup_out(a2_wr[635]), .rdlo_out(a2_wr[891]));
			radix2 #(.width(width)) rd_st1_636  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[636]), .rdlo_in(a1_wr[892]),  .coef_in(coef[248]), .rdup_out(a2_wr[636]), .rdlo_out(a2_wr[892]));
			radix2 #(.width(width)) rd_st1_637  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[637]), .rdlo_in(a1_wr[893]),  .coef_in(coef[250]), .rdup_out(a2_wr[637]), .rdlo_out(a2_wr[893]));
			radix2 #(.width(width)) rd_st1_638  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[638]), .rdlo_in(a1_wr[894]),  .coef_in(coef[252]), .rdup_out(a2_wr[638]), .rdlo_out(a2_wr[894]));
			radix2 #(.width(width)) rd_st1_639  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[639]), .rdlo_in(a1_wr[895]),  .coef_in(coef[254]), .rdup_out(a2_wr[639]), .rdlo_out(a2_wr[895]));
			radix2 #(.width(width)) rd_st1_640  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[640]), .rdlo_in(a1_wr[896]),  .coef_in(coef[256]), .rdup_out(a2_wr[640]), .rdlo_out(a2_wr[896]));
			radix2 #(.width(width)) rd_st1_641  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[641]), .rdlo_in(a1_wr[897]),  .coef_in(coef[258]), .rdup_out(a2_wr[641]), .rdlo_out(a2_wr[897]));
			radix2 #(.width(width)) rd_st1_642  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[642]), .rdlo_in(a1_wr[898]),  .coef_in(coef[260]), .rdup_out(a2_wr[642]), .rdlo_out(a2_wr[898]));
			radix2 #(.width(width)) rd_st1_643  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[643]), .rdlo_in(a1_wr[899]),  .coef_in(coef[262]), .rdup_out(a2_wr[643]), .rdlo_out(a2_wr[899]));
			radix2 #(.width(width)) rd_st1_644  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[644]), .rdlo_in(a1_wr[900]),  .coef_in(coef[264]), .rdup_out(a2_wr[644]), .rdlo_out(a2_wr[900]));
			radix2 #(.width(width)) rd_st1_645  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[645]), .rdlo_in(a1_wr[901]),  .coef_in(coef[266]), .rdup_out(a2_wr[645]), .rdlo_out(a2_wr[901]));
			radix2 #(.width(width)) rd_st1_646  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[646]), .rdlo_in(a1_wr[902]),  .coef_in(coef[268]), .rdup_out(a2_wr[646]), .rdlo_out(a2_wr[902]));
			radix2 #(.width(width)) rd_st1_647  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[647]), .rdlo_in(a1_wr[903]),  .coef_in(coef[270]), .rdup_out(a2_wr[647]), .rdlo_out(a2_wr[903]));
			radix2 #(.width(width)) rd_st1_648  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[648]), .rdlo_in(a1_wr[904]),  .coef_in(coef[272]), .rdup_out(a2_wr[648]), .rdlo_out(a2_wr[904]));
			radix2 #(.width(width)) rd_st1_649  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[649]), .rdlo_in(a1_wr[905]),  .coef_in(coef[274]), .rdup_out(a2_wr[649]), .rdlo_out(a2_wr[905]));
			radix2 #(.width(width)) rd_st1_650  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[650]), .rdlo_in(a1_wr[906]),  .coef_in(coef[276]), .rdup_out(a2_wr[650]), .rdlo_out(a2_wr[906]));
			radix2 #(.width(width)) rd_st1_651  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[651]), .rdlo_in(a1_wr[907]),  .coef_in(coef[278]), .rdup_out(a2_wr[651]), .rdlo_out(a2_wr[907]));
			radix2 #(.width(width)) rd_st1_652  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[652]), .rdlo_in(a1_wr[908]),  .coef_in(coef[280]), .rdup_out(a2_wr[652]), .rdlo_out(a2_wr[908]));
			radix2 #(.width(width)) rd_st1_653  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[653]), .rdlo_in(a1_wr[909]),  .coef_in(coef[282]), .rdup_out(a2_wr[653]), .rdlo_out(a2_wr[909]));
			radix2 #(.width(width)) rd_st1_654  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[654]), .rdlo_in(a1_wr[910]),  .coef_in(coef[284]), .rdup_out(a2_wr[654]), .rdlo_out(a2_wr[910]));
			radix2 #(.width(width)) rd_st1_655  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[655]), .rdlo_in(a1_wr[911]),  .coef_in(coef[286]), .rdup_out(a2_wr[655]), .rdlo_out(a2_wr[911]));
			radix2 #(.width(width)) rd_st1_656  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[656]), .rdlo_in(a1_wr[912]),  .coef_in(coef[288]), .rdup_out(a2_wr[656]), .rdlo_out(a2_wr[912]));
			radix2 #(.width(width)) rd_st1_657  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[657]), .rdlo_in(a1_wr[913]),  .coef_in(coef[290]), .rdup_out(a2_wr[657]), .rdlo_out(a2_wr[913]));
			radix2 #(.width(width)) rd_st1_658  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[658]), .rdlo_in(a1_wr[914]),  .coef_in(coef[292]), .rdup_out(a2_wr[658]), .rdlo_out(a2_wr[914]));
			radix2 #(.width(width)) rd_st1_659  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[659]), .rdlo_in(a1_wr[915]),  .coef_in(coef[294]), .rdup_out(a2_wr[659]), .rdlo_out(a2_wr[915]));
			radix2 #(.width(width)) rd_st1_660  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[660]), .rdlo_in(a1_wr[916]),  .coef_in(coef[296]), .rdup_out(a2_wr[660]), .rdlo_out(a2_wr[916]));
			radix2 #(.width(width)) rd_st1_661  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[661]), .rdlo_in(a1_wr[917]),  .coef_in(coef[298]), .rdup_out(a2_wr[661]), .rdlo_out(a2_wr[917]));
			radix2 #(.width(width)) rd_st1_662  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[662]), .rdlo_in(a1_wr[918]),  .coef_in(coef[300]), .rdup_out(a2_wr[662]), .rdlo_out(a2_wr[918]));
			radix2 #(.width(width)) rd_st1_663  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[663]), .rdlo_in(a1_wr[919]),  .coef_in(coef[302]), .rdup_out(a2_wr[663]), .rdlo_out(a2_wr[919]));
			radix2 #(.width(width)) rd_st1_664  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[664]), .rdlo_in(a1_wr[920]),  .coef_in(coef[304]), .rdup_out(a2_wr[664]), .rdlo_out(a2_wr[920]));
			radix2 #(.width(width)) rd_st1_665  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[665]), .rdlo_in(a1_wr[921]),  .coef_in(coef[306]), .rdup_out(a2_wr[665]), .rdlo_out(a2_wr[921]));
			radix2 #(.width(width)) rd_st1_666  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[666]), .rdlo_in(a1_wr[922]),  .coef_in(coef[308]), .rdup_out(a2_wr[666]), .rdlo_out(a2_wr[922]));
			radix2 #(.width(width)) rd_st1_667  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[667]), .rdlo_in(a1_wr[923]),  .coef_in(coef[310]), .rdup_out(a2_wr[667]), .rdlo_out(a2_wr[923]));
			radix2 #(.width(width)) rd_st1_668  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[668]), .rdlo_in(a1_wr[924]),  .coef_in(coef[312]), .rdup_out(a2_wr[668]), .rdlo_out(a2_wr[924]));
			radix2 #(.width(width)) rd_st1_669  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[669]), .rdlo_in(a1_wr[925]),  .coef_in(coef[314]), .rdup_out(a2_wr[669]), .rdlo_out(a2_wr[925]));
			radix2 #(.width(width)) rd_st1_670  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[670]), .rdlo_in(a1_wr[926]),  .coef_in(coef[316]), .rdup_out(a2_wr[670]), .rdlo_out(a2_wr[926]));
			radix2 #(.width(width)) rd_st1_671  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[671]), .rdlo_in(a1_wr[927]),  .coef_in(coef[318]), .rdup_out(a2_wr[671]), .rdlo_out(a2_wr[927]));
			radix2 #(.width(width)) rd_st1_672  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[672]), .rdlo_in(a1_wr[928]),  .coef_in(coef[320]), .rdup_out(a2_wr[672]), .rdlo_out(a2_wr[928]));
			radix2 #(.width(width)) rd_st1_673  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[673]), .rdlo_in(a1_wr[929]),  .coef_in(coef[322]), .rdup_out(a2_wr[673]), .rdlo_out(a2_wr[929]));
			radix2 #(.width(width)) rd_st1_674  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[674]), .rdlo_in(a1_wr[930]),  .coef_in(coef[324]), .rdup_out(a2_wr[674]), .rdlo_out(a2_wr[930]));
			radix2 #(.width(width)) rd_st1_675  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[675]), .rdlo_in(a1_wr[931]),  .coef_in(coef[326]), .rdup_out(a2_wr[675]), .rdlo_out(a2_wr[931]));
			radix2 #(.width(width)) rd_st1_676  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[676]), .rdlo_in(a1_wr[932]),  .coef_in(coef[328]), .rdup_out(a2_wr[676]), .rdlo_out(a2_wr[932]));
			radix2 #(.width(width)) rd_st1_677  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[677]), .rdlo_in(a1_wr[933]),  .coef_in(coef[330]), .rdup_out(a2_wr[677]), .rdlo_out(a2_wr[933]));
			radix2 #(.width(width)) rd_st1_678  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[678]), .rdlo_in(a1_wr[934]),  .coef_in(coef[332]), .rdup_out(a2_wr[678]), .rdlo_out(a2_wr[934]));
			radix2 #(.width(width)) rd_st1_679  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[679]), .rdlo_in(a1_wr[935]),  .coef_in(coef[334]), .rdup_out(a2_wr[679]), .rdlo_out(a2_wr[935]));
			radix2 #(.width(width)) rd_st1_680  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[680]), .rdlo_in(a1_wr[936]),  .coef_in(coef[336]), .rdup_out(a2_wr[680]), .rdlo_out(a2_wr[936]));
			radix2 #(.width(width)) rd_st1_681  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[681]), .rdlo_in(a1_wr[937]),  .coef_in(coef[338]), .rdup_out(a2_wr[681]), .rdlo_out(a2_wr[937]));
			radix2 #(.width(width)) rd_st1_682  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[682]), .rdlo_in(a1_wr[938]),  .coef_in(coef[340]), .rdup_out(a2_wr[682]), .rdlo_out(a2_wr[938]));
			radix2 #(.width(width)) rd_st1_683  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[683]), .rdlo_in(a1_wr[939]),  .coef_in(coef[342]), .rdup_out(a2_wr[683]), .rdlo_out(a2_wr[939]));
			radix2 #(.width(width)) rd_st1_684  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[684]), .rdlo_in(a1_wr[940]),  .coef_in(coef[344]), .rdup_out(a2_wr[684]), .rdlo_out(a2_wr[940]));
			radix2 #(.width(width)) rd_st1_685  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[685]), .rdlo_in(a1_wr[941]),  .coef_in(coef[346]), .rdup_out(a2_wr[685]), .rdlo_out(a2_wr[941]));
			radix2 #(.width(width)) rd_st1_686  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[686]), .rdlo_in(a1_wr[942]),  .coef_in(coef[348]), .rdup_out(a2_wr[686]), .rdlo_out(a2_wr[942]));
			radix2 #(.width(width)) rd_st1_687  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[687]), .rdlo_in(a1_wr[943]),  .coef_in(coef[350]), .rdup_out(a2_wr[687]), .rdlo_out(a2_wr[943]));
			radix2 #(.width(width)) rd_st1_688  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[688]), .rdlo_in(a1_wr[944]),  .coef_in(coef[352]), .rdup_out(a2_wr[688]), .rdlo_out(a2_wr[944]));
			radix2 #(.width(width)) rd_st1_689  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[689]), .rdlo_in(a1_wr[945]),  .coef_in(coef[354]), .rdup_out(a2_wr[689]), .rdlo_out(a2_wr[945]));
			radix2 #(.width(width)) rd_st1_690  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[690]), .rdlo_in(a1_wr[946]),  .coef_in(coef[356]), .rdup_out(a2_wr[690]), .rdlo_out(a2_wr[946]));
			radix2 #(.width(width)) rd_st1_691  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[691]), .rdlo_in(a1_wr[947]),  .coef_in(coef[358]), .rdup_out(a2_wr[691]), .rdlo_out(a2_wr[947]));
			radix2 #(.width(width)) rd_st1_692  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[692]), .rdlo_in(a1_wr[948]),  .coef_in(coef[360]), .rdup_out(a2_wr[692]), .rdlo_out(a2_wr[948]));
			radix2 #(.width(width)) rd_st1_693  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[693]), .rdlo_in(a1_wr[949]),  .coef_in(coef[362]), .rdup_out(a2_wr[693]), .rdlo_out(a2_wr[949]));
			radix2 #(.width(width)) rd_st1_694  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[694]), .rdlo_in(a1_wr[950]),  .coef_in(coef[364]), .rdup_out(a2_wr[694]), .rdlo_out(a2_wr[950]));
			radix2 #(.width(width)) rd_st1_695  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[695]), .rdlo_in(a1_wr[951]),  .coef_in(coef[366]), .rdup_out(a2_wr[695]), .rdlo_out(a2_wr[951]));
			radix2 #(.width(width)) rd_st1_696  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[696]), .rdlo_in(a1_wr[952]),  .coef_in(coef[368]), .rdup_out(a2_wr[696]), .rdlo_out(a2_wr[952]));
			radix2 #(.width(width)) rd_st1_697  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[697]), .rdlo_in(a1_wr[953]),  .coef_in(coef[370]), .rdup_out(a2_wr[697]), .rdlo_out(a2_wr[953]));
			radix2 #(.width(width)) rd_st1_698  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[698]), .rdlo_in(a1_wr[954]),  .coef_in(coef[372]), .rdup_out(a2_wr[698]), .rdlo_out(a2_wr[954]));
			radix2 #(.width(width)) rd_st1_699  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[699]), .rdlo_in(a1_wr[955]),  .coef_in(coef[374]), .rdup_out(a2_wr[699]), .rdlo_out(a2_wr[955]));
			radix2 #(.width(width)) rd_st1_700  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[700]), .rdlo_in(a1_wr[956]),  .coef_in(coef[376]), .rdup_out(a2_wr[700]), .rdlo_out(a2_wr[956]));
			radix2 #(.width(width)) rd_st1_701  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[701]), .rdlo_in(a1_wr[957]),  .coef_in(coef[378]), .rdup_out(a2_wr[701]), .rdlo_out(a2_wr[957]));
			radix2 #(.width(width)) rd_st1_702  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[702]), .rdlo_in(a1_wr[958]),  .coef_in(coef[380]), .rdup_out(a2_wr[702]), .rdlo_out(a2_wr[958]));
			radix2 #(.width(width)) rd_st1_703  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[703]), .rdlo_in(a1_wr[959]),  .coef_in(coef[382]), .rdup_out(a2_wr[703]), .rdlo_out(a2_wr[959]));
			radix2 #(.width(width)) rd_st1_704  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[704]), .rdlo_in(a1_wr[960]),  .coef_in(coef[384]), .rdup_out(a2_wr[704]), .rdlo_out(a2_wr[960]));
			radix2 #(.width(width)) rd_st1_705  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[705]), .rdlo_in(a1_wr[961]),  .coef_in(coef[386]), .rdup_out(a2_wr[705]), .rdlo_out(a2_wr[961]));
			radix2 #(.width(width)) rd_st1_706  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[706]), .rdlo_in(a1_wr[962]),  .coef_in(coef[388]), .rdup_out(a2_wr[706]), .rdlo_out(a2_wr[962]));
			radix2 #(.width(width)) rd_st1_707  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[707]), .rdlo_in(a1_wr[963]),  .coef_in(coef[390]), .rdup_out(a2_wr[707]), .rdlo_out(a2_wr[963]));
			radix2 #(.width(width)) rd_st1_708  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[708]), .rdlo_in(a1_wr[964]),  .coef_in(coef[392]), .rdup_out(a2_wr[708]), .rdlo_out(a2_wr[964]));
			radix2 #(.width(width)) rd_st1_709  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[709]), .rdlo_in(a1_wr[965]),  .coef_in(coef[394]), .rdup_out(a2_wr[709]), .rdlo_out(a2_wr[965]));
			radix2 #(.width(width)) rd_st1_710  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[710]), .rdlo_in(a1_wr[966]),  .coef_in(coef[396]), .rdup_out(a2_wr[710]), .rdlo_out(a2_wr[966]));
			radix2 #(.width(width)) rd_st1_711  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[711]), .rdlo_in(a1_wr[967]),  .coef_in(coef[398]), .rdup_out(a2_wr[711]), .rdlo_out(a2_wr[967]));
			radix2 #(.width(width)) rd_st1_712  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[712]), .rdlo_in(a1_wr[968]),  .coef_in(coef[400]), .rdup_out(a2_wr[712]), .rdlo_out(a2_wr[968]));
			radix2 #(.width(width)) rd_st1_713  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[713]), .rdlo_in(a1_wr[969]),  .coef_in(coef[402]), .rdup_out(a2_wr[713]), .rdlo_out(a2_wr[969]));
			radix2 #(.width(width)) rd_st1_714  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[714]), .rdlo_in(a1_wr[970]),  .coef_in(coef[404]), .rdup_out(a2_wr[714]), .rdlo_out(a2_wr[970]));
			radix2 #(.width(width)) rd_st1_715  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[715]), .rdlo_in(a1_wr[971]),  .coef_in(coef[406]), .rdup_out(a2_wr[715]), .rdlo_out(a2_wr[971]));
			radix2 #(.width(width)) rd_st1_716  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[716]), .rdlo_in(a1_wr[972]),  .coef_in(coef[408]), .rdup_out(a2_wr[716]), .rdlo_out(a2_wr[972]));
			radix2 #(.width(width)) rd_st1_717  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[717]), .rdlo_in(a1_wr[973]),  .coef_in(coef[410]), .rdup_out(a2_wr[717]), .rdlo_out(a2_wr[973]));
			radix2 #(.width(width)) rd_st1_718  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[718]), .rdlo_in(a1_wr[974]),  .coef_in(coef[412]), .rdup_out(a2_wr[718]), .rdlo_out(a2_wr[974]));
			radix2 #(.width(width)) rd_st1_719  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[719]), .rdlo_in(a1_wr[975]),  .coef_in(coef[414]), .rdup_out(a2_wr[719]), .rdlo_out(a2_wr[975]));
			radix2 #(.width(width)) rd_st1_720  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[720]), .rdlo_in(a1_wr[976]),  .coef_in(coef[416]), .rdup_out(a2_wr[720]), .rdlo_out(a2_wr[976]));
			radix2 #(.width(width)) rd_st1_721  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[721]), .rdlo_in(a1_wr[977]),  .coef_in(coef[418]), .rdup_out(a2_wr[721]), .rdlo_out(a2_wr[977]));
			radix2 #(.width(width)) rd_st1_722  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[722]), .rdlo_in(a1_wr[978]),  .coef_in(coef[420]), .rdup_out(a2_wr[722]), .rdlo_out(a2_wr[978]));
			radix2 #(.width(width)) rd_st1_723  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[723]), .rdlo_in(a1_wr[979]),  .coef_in(coef[422]), .rdup_out(a2_wr[723]), .rdlo_out(a2_wr[979]));
			radix2 #(.width(width)) rd_st1_724  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[724]), .rdlo_in(a1_wr[980]),  .coef_in(coef[424]), .rdup_out(a2_wr[724]), .rdlo_out(a2_wr[980]));
			radix2 #(.width(width)) rd_st1_725  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[725]), .rdlo_in(a1_wr[981]),  .coef_in(coef[426]), .rdup_out(a2_wr[725]), .rdlo_out(a2_wr[981]));
			radix2 #(.width(width)) rd_st1_726  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[726]), .rdlo_in(a1_wr[982]),  .coef_in(coef[428]), .rdup_out(a2_wr[726]), .rdlo_out(a2_wr[982]));
			radix2 #(.width(width)) rd_st1_727  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[727]), .rdlo_in(a1_wr[983]),  .coef_in(coef[430]), .rdup_out(a2_wr[727]), .rdlo_out(a2_wr[983]));
			radix2 #(.width(width)) rd_st1_728  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[728]), .rdlo_in(a1_wr[984]),  .coef_in(coef[432]), .rdup_out(a2_wr[728]), .rdlo_out(a2_wr[984]));
			radix2 #(.width(width)) rd_st1_729  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[729]), .rdlo_in(a1_wr[985]),  .coef_in(coef[434]), .rdup_out(a2_wr[729]), .rdlo_out(a2_wr[985]));
			radix2 #(.width(width)) rd_st1_730  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[730]), .rdlo_in(a1_wr[986]),  .coef_in(coef[436]), .rdup_out(a2_wr[730]), .rdlo_out(a2_wr[986]));
			radix2 #(.width(width)) rd_st1_731  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[731]), .rdlo_in(a1_wr[987]),  .coef_in(coef[438]), .rdup_out(a2_wr[731]), .rdlo_out(a2_wr[987]));
			radix2 #(.width(width)) rd_st1_732  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[732]), .rdlo_in(a1_wr[988]),  .coef_in(coef[440]), .rdup_out(a2_wr[732]), .rdlo_out(a2_wr[988]));
			radix2 #(.width(width)) rd_st1_733  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[733]), .rdlo_in(a1_wr[989]),  .coef_in(coef[442]), .rdup_out(a2_wr[733]), .rdlo_out(a2_wr[989]));
			radix2 #(.width(width)) rd_st1_734  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[734]), .rdlo_in(a1_wr[990]),  .coef_in(coef[444]), .rdup_out(a2_wr[734]), .rdlo_out(a2_wr[990]));
			radix2 #(.width(width)) rd_st1_735  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[735]), .rdlo_in(a1_wr[991]),  .coef_in(coef[446]), .rdup_out(a2_wr[735]), .rdlo_out(a2_wr[991]));
			radix2 #(.width(width)) rd_st1_736  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[736]), .rdlo_in(a1_wr[992]),  .coef_in(coef[448]), .rdup_out(a2_wr[736]), .rdlo_out(a2_wr[992]));
			radix2 #(.width(width)) rd_st1_737  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[737]), .rdlo_in(a1_wr[993]),  .coef_in(coef[450]), .rdup_out(a2_wr[737]), .rdlo_out(a2_wr[993]));
			radix2 #(.width(width)) rd_st1_738  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[738]), .rdlo_in(a1_wr[994]),  .coef_in(coef[452]), .rdup_out(a2_wr[738]), .rdlo_out(a2_wr[994]));
			radix2 #(.width(width)) rd_st1_739  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[739]), .rdlo_in(a1_wr[995]),  .coef_in(coef[454]), .rdup_out(a2_wr[739]), .rdlo_out(a2_wr[995]));
			radix2 #(.width(width)) rd_st1_740  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[740]), .rdlo_in(a1_wr[996]),  .coef_in(coef[456]), .rdup_out(a2_wr[740]), .rdlo_out(a2_wr[996]));
			radix2 #(.width(width)) rd_st1_741  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[741]), .rdlo_in(a1_wr[997]),  .coef_in(coef[458]), .rdup_out(a2_wr[741]), .rdlo_out(a2_wr[997]));
			radix2 #(.width(width)) rd_st1_742  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[742]), .rdlo_in(a1_wr[998]),  .coef_in(coef[460]), .rdup_out(a2_wr[742]), .rdlo_out(a2_wr[998]));
			radix2 #(.width(width)) rd_st1_743  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[743]), .rdlo_in(a1_wr[999]),  .coef_in(coef[462]), .rdup_out(a2_wr[743]), .rdlo_out(a2_wr[999]));
			radix2 #(.width(width)) rd_st1_744  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[744]), .rdlo_in(a1_wr[1000]),  .coef_in(coef[464]), .rdup_out(a2_wr[744]), .rdlo_out(a2_wr[1000]));
			radix2 #(.width(width)) rd_st1_745  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[745]), .rdlo_in(a1_wr[1001]),  .coef_in(coef[466]), .rdup_out(a2_wr[745]), .rdlo_out(a2_wr[1001]));
			radix2 #(.width(width)) rd_st1_746  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[746]), .rdlo_in(a1_wr[1002]),  .coef_in(coef[468]), .rdup_out(a2_wr[746]), .rdlo_out(a2_wr[1002]));
			radix2 #(.width(width)) rd_st1_747  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[747]), .rdlo_in(a1_wr[1003]),  .coef_in(coef[470]), .rdup_out(a2_wr[747]), .rdlo_out(a2_wr[1003]));
			radix2 #(.width(width)) rd_st1_748  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[748]), .rdlo_in(a1_wr[1004]),  .coef_in(coef[472]), .rdup_out(a2_wr[748]), .rdlo_out(a2_wr[1004]));
			radix2 #(.width(width)) rd_st1_749  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[749]), .rdlo_in(a1_wr[1005]),  .coef_in(coef[474]), .rdup_out(a2_wr[749]), .rdlo_out(a2_wr[1005]));
			radix2 #(.width(width)) rd_st1_750  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[750]), .rdlo_in(a1_wr[1006]),  .coef_in(coef[476]), .rdup_out(a2_wr[750]), .rdlo_out(a2_wr[1006]));
			radix2 #(.width(width)) rd_st1_751  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[751]), .rdlo_in(a1_wr[1007]),  .coef_in(coef[478]), .rdup_out(a2_wr[751]), .rdlo_out(a2_wr[1007]));
			radix2 #(.width(width)) rd_st1_752  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[752]), .rdlo_in(a1_wr[1008]),  .coef_in(coef[480]), .rdup_out(a2_wr[752]), .rdlo_out(a2_wr[1008]));
			radix2 #(.width(width)) rd_st1_753  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[753]), .rdlo_in(a1_wr[1009]),  .coef_in(coef[482]), .rdup_out(a2_wr[753]), .rdlo_out(a2_wr[1009]));
			radix2 #(.width(width)) rd_st1_754  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[754]), .rdlo_in(a1_wr[1010]),  .coef_in(coef[484]), .rdup_out(a2_wr[754]), .rdlo_out(a2_wr[1010]));
			radix2 #(.width(width)) rd_st1_755  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[755]), .rdlo_in(a1_wr[1011]),  .coef_in(coef[486]), .rdup_out(a2_wr[755]), .rdlo_out(a2_wr[1011]));
			radix2 #(.width(width)) rd_st1_756  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[756]), .rdlo_in(a1_wr[1012]),  .coef_in(coef[488]), .rdup_out(a2_wr[756]), .rdlo_out(a2_wr[1012]));
			radix2 #(.width(width)) rd_st1_757  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[757]), .rdlo_in(a1_wr[1013]),  .coef_in(coef[490]), .rdup_out(a2_wr[757]), .rdlo_out(a2_wr[1013]));
			radix2 #(.width(width)) rd_st1_758  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[758]), .rdlo_in(a1_wr[1014]),  .coef_in(coef[492]), .rdup_out(a2_wr[758]), .rdlo_out(a2_wr[1014]));
			radix2 #(.width(width)) rd_st1_759  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[759]), .rdlo_in(a1_wr[1015]),  .coef_in(coef[494]), .rdup_out(a2_wr[759]), .rdlo_out(a2_wr[1015]));
			radix2 #(.width(width)) rd_st1_760  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[760]), .rdlo_in(a1_wr[1016]),  .coef_in(coef[496]), .rdup_out(a2_wr[760]), .rdlo_out(a2_wr[1016]));
			radix2 #(.width(width)) rd_st1_761  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[761]), .rdlo_in(a1_wr[1017]),  .coef_in(coef[498]), .rdup_out(a2_wr[761]), .rdlo_out(a2_wr[1017]));
			radix2 #(.width(width)) rd_st1_762  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[762]), .rdlo_in(a1_wr[1018]),  .coef_in(coef[500]), .rdup_out(a2_wr[762]), .rdlo_out(a2_wr[1018]));
			radix2 #(.width(width)) rd_st1_763  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[763]), .rdlo_in(a1_wr[1019]),  .coef_in(coef[502]), .rdup_out(a2_wr[763]), .rdlo_out(a2_wr[1019]));
			radix2 #(.width(width)) rd_st1_764  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[764]), .rdlo_in(a1_wr[1020]),  .coef_in(coef[504]), .rdup_out(a2_wr[764]), .rdlo_out(a2_wr[1020]));
			radix2 #(.width(width)) rd_st1_765  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[765]), .rdlo_in(a1_wr[1021]),  .coef_in(coef[506]), .rdup_out(a2_wr[765]), .rdlo_out(a2_wr[1021]));
			radix2 #(.width(width)) rd_st1_766  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[766]), .rdlo_in(a1_wr[1022]),  .coef_in(coef[508]), .rdup_out(a2_wr[766]), .rdlo_out(a2_wr[1022]));
			radix2 #(.width(width)) rd_st1_767  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[767]), .rdlo_in(a1_wr[1023]),  .coef_in(coef[510]), .rdup_out(a2_wr[767]), .rdlo_out(a2_wr[1023]));

		//--- radix stage 2
			radix2 #(.width(width)) rd_st2_0   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[0]), .rdlo_in(a2_wr[128]),  .coef_in(coef[0]), .rdup_out(a3_wr[0]), .rdlo_out(a3_wr[128]));
			radix2 #(.width(width)) rd_st2_1   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1]), .rdlo_in(a2_wr[129]),  .coef_in(coef[4]), .rdup_out(a3_wr[1]), .rdlo_out(a3_wr[129]));
			radix2 #(.width(width)) rd_st2_2   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[2]), .rdlo_in(a2_wr[130]),  .coef_in(coef[8]), .rdup_out(a3_wr[2]), .rdlo_out(a3_wr[130]));
			radix2 #(.width(width)) rd_st2_3   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[3]), .rdlo_in(a2_wr[131]),  .coef_in(coef[12]), .rdup_out(a3_wr[3]), .rdlo_out(a3_wr[131]));
			radix2 #(.width(width)) rd_st2_4   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[4]), .rdlo_in(a2_wr[132]),  .coef_in(coef[16]), .rdup_out(a3_wr[4]), .rdlo_out(a3_wr[132]));
			radix2 #(.width(width)) rd_st2_5   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[5]), .rdlo_in(a2_wr[133]),  .coef_in(coef[20]), .rdup_out(a3_wr[5]), .rdlo_out(a3_wr[133]));
			radix2 #(.width(width)) rd_st2_6   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[6]), .rdlo_in(a2_wr[134]),  .coef_in(coef[24]), .rdup_out(a3_wr[6]), .rdlo_out(a3_wr[134]));
			radix2 #(.width(width)) rd_st2_7   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[7]), .rdlo_in(a2_wr[135]),  .coef_in(coef[28]), .rdup_out(a3_wr[7]), .rdlo_out(a3_wr[135]));
			radix2 #(.width(width)) rd_st2_8   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[8]), .rdlo_in(a2_wr[136]),  .coef_in(coef[32]), .rdup_out(a3_wr[8]), .rdlo_out(a3_wr[136]));
			radix2 #(.width(width)) rd_st2_9   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[9]), .rdlo_in(a2_wr[137]),  .coef_in(coef[36]), .rdup_out(a3_wr[9]), .rdlo_out(a3_wr[137]));
			radix2 #(.width(width)) rd_st2_10  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[10]), .rdlo_in(a2_wr[138]),  .coef_in(coef[40]), .rdup_out(a3_wr[10]), .rdlo_out(a3_wr[138]));
			radix2 #(.width(width)) rd_st2_11  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[11]), .rdlo_in(a2_wr[139]),  .coef_in(coef[44]), .rdup_out(a3_wr[11]), .rdlo_out(a3_wr[139]));
			radix2 #(.width(width)) rd_st2_12  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[12]), .rdlo_in(a2_wr[140]),  .coef_in(coef[48]), .rdup_out(a3_wr[12]), .rdlo_out(a3_wr[140]));
			radix2 #(.width(width)) rd_st2_13  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[13]), .rdlo_in(a2_wr[141]),  .coef_in(coef[52]), .rdup_out(a3_wr[13]), .rdlo_out(a3_wr[141]));
			radix2 #(.width(width)) rd_st2_14  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[14]), .rdlo_in(a2_wr[142]),  .coef_in(coef[56]), .rdup_out(a3_wr[14]), .rdlo_out(a3_wr[142]));
			radix2 #(.width(width)) rd_st2_15  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[15]), .rdlo_in(a2_wr[143]),  .coef_in(coef[60]), .rdup_out(a3_wr[15]), .rdlo_out(a3_wr[143]));
			radix2 #(.width(width)) rd_st2_16  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[16]), .rdlo_in(a2_wr[144]),  .coef_in(coef[64]), .rdup_out(a3_wr[16]), .rdlo_out(a3_wr[144]));
			radix2 #(.width(width)) rd_st2_17  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[17]), .rdlo_in(a2_wr[145]),  .coef_in(coef[68]), .rdup_out(a3_wr[17]), .rdlo_out(a3_wr[145]));
			radix2 #(.width(width)) rd_st2_18  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[18]), .rdlo_in(a2_wr[146]),  .coef_in(coef[72]), .rdup_out(a3_wr[18]), .rdlo_out(a3_wr[146]));
			radix2 #(.width(width)) rd_st2_19  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[19]), .rdlo_in(a2_wr[147]),  .coef_in(coef[76]), .rdup_out(a3_wr[19]), .rdlo_out(a3_wr[147]));
			radix2 #(.width(width)) rd_st2_20  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[20]), .rdlo_in(a2_wr[148]),  .coef_in(coef[80]), .rdup_out(a3_wr[20]), .rdlo_out(a3_wr[148]));
			radix2 #(.width(width)) rd_st2_21  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[21]), .rdlo_in(a2_wr[149]),  .coef_in(coef[84]), .rdup_out(a3_wr[21]), .rdlo_out(a3_wr[149]));
			radix2 #(.width(width)) rd_st2_22  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[22]), .rdlo_in(a2_wr[150]),  .coef_in(coef[88]), .rdup_out(a3_wr[22]), .rdlo_out(a3_wr[150]));
			radix2 #(.width(width)) rd_st2_23  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[23]), .rdlo_in(a2_wr[151]),  .coef_in(coef[92]), .rdup_out(a3_wr[23]), .rdlo_out(a3_wr[151]));
			radix2 #(.width(width)) rd_st2_24  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[24]), .rdlo_in(a2_wr[152]),  .coef_in(coef[96]), .rdup_out(a3_wr[24]), .rdlo_out(a3_wr[152]));
			radix2 #(.width(width)) rd_st2_25  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[25]), .rdlo_in(a2_wr[153]),  .coef_in(coef[100]), .rdup_out(a3_wr[25]), .rdlo_out(a3_wr[153]));
			radix2 #(.width(width)) rd_st2_26  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[26]), .rdlo_in(a2_wr[154]),  .coef_in(coef[104]), .rdup_out(a3_wr[26]), .rdlo_out(a3_wr[154]));
			radix2 #(.width(width)) rd_st2_27  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[27]), .rdlo_in(a2_wr[155]),  .coef_in(coef[108]), .rdup_out(a3_wr[27]), .rdlo_out(a3_wr[155]));
			radix2 #(.width(width)) rd_st2_28  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[28]), .rdlo_in(a2_wr[156]),  .coef_in(coef[112]), .rdup_out(a3_wr[28]), .rdlo_out(a3_wr[156]));
			radix2 #(.width(width)) rd_st2_29  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[29]), .rdlo_in(a2_wr[157]),  .coef_in(coef[116]), .rdup_out(a3_wr[29]), .rdlo_out(a3_wr[157]));
			radix2 #(.width(width)) rd_st2_30  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[30]), .rdlo_in(a2_wr[158]),  .coef_in(coef[120]), .rdup_out(a3_wr[30]), .rdlo_out(a3_wr[158]));
			radix2 #(.width(width)) rd_st2_31  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[31]), .rdlo_in(a2_wr[159]),  .coef_in(coef[124]), .rdup_out(a3_wr[31]), .rdlo_out(a3_wr[159]));
			radix2 #(.width(width)) rd_st2_32  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[32]), .rdlo_in(a2_wr[160]),  .coef_in(coef[128]), .rdup_out(a3_wr[32]), .rdlo_out(a3_wr[160]));
			radix2 #(.width(width)) rd_st2_33  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[33]), .rdlo_in(a2_wr[161]),  .coef_in(coef[132]), .rdup_out(a3_wr[33]), .rdlo_out(a3_wr[161]));
			radix2 #(.width(width)) rd_st2_34  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[34]), .rdlo_in(a2_wr[162]),  .coef_in(coef[136]), .rdup_out(a3_wr[34]), .rdlo_out(a3_wr[162]));
			radix2 #(.width(width)) rd_st2_35  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[35]), .rdlo_in(a2_wr[163]),  .coef_in(coef[140]), .rdup_out(a3_wr[35]), .rdlo_out(a3_wr[163]));
			radix2 #(.width(width)) rd_st2_36  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[36]), .rdlo_in(a2_wr[164]),  .coef_in(coef[144]), .rdup_out(a3_wr[36]), .rdlo_out(a3_wr[164]));
			radix2 #(.width(width)) rd_st2_37  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[37]), .rdlo_in(a2_wr[165]),  .coef_in(coef[148]), .rdup_out(a3_wr[37]), .rdlo_out(a3_wr[165]));
			radix2 #(.width(width)) rd_st2_38  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[38]), .rdlo_in(a2_wr[166]),  .coef_in(coef[152]), .rdup_out(a3_wr[38]), .rdlo_out(a3_wr[166]));
			radix2 #(.width(width)) rd_st2_39  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[39]), .rdlo_in(a2_wr[167]),  .coef_in(coef[156]), .rdup_out(a3_wr[39]), .rdlo_out(a3_wr[167]));
			radix2 #(.width(width)) rd_st2_40  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[40]), .rdlo_in(a2_wr[168]),  .coef_in(coef[160]), .rdup_out(a3_wr[40]), .rdlo_out(a3_wr[168]));
			radix2 #(.width(width)) rd_st2_41  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[41]), .rdlo_in(a2_wr[169]),  .coef_in(coef[164]), .rdup_out(a3_wr[41]), .rdlo_out(a3_wr[169]));
			radix2 #(.width(width)) rd_st2_42  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[42]), .rdlo_in(a2_wr[170]),  .coef_in(coef[168]), .rdup_out(a3_wr[42]), .rdlo_out(a3_wr[170]));
			radix2 #(.width(width)) rd_st2_43  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[43]), .rdlo_in(a2_wr[171]),  .coef_in(coef[172]), .rdup_out(a3_wr[43]), .rdlo_out(a3_wr[171]));
			radix2 #(.width(width)) rd_st2_44  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[44]), .rdlo_in(a2_wr[172]),  .coef_in(coef[176]), .rdup_out(a3_wr[44]), .rdlo_out(a3_wr[172]));
			radix2 #(.width(width)) rd_st2_45  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[45]), .rdlo_in(a2_wr[173]),  .coef_in(coef[180]), .rdup_out(a3_wr[45]), .rdlo_out(a3_wr[173]));
			radix2 #(.width(width)) rd_st2_46  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[46]), .rdlo_in(a2_wr[174]),  .coef_in(coef[184]), .rdup_out(a3_wr[46]), .rdlo_out(a3_wr[174]));
			radix2 #(.width(width)) rd_st2_47  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[47]), .rdlo_in(a2_wr[175]),  .coef_in(coef[188]), .rdup_out(a3_wr[47]), .rdlo_out(a3_wr[175]));
			radix2 #(.width(width)) rd_st2_48  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[48]), .rdlo_in(a2_wr[176]),  .coef_in(coef[192]), .rdup_out(a3_wr[48]), .rdlo_out(a3_wr[176]));
			radix2 #(.width(width)) rd_st2_49  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[49]), .rdlo_in(a2_wr[177]),  .coef_in(coef[196]), .rdup_out(a3_wr[49]), .rdlo_out(a3_wr[177]));
			radix2 #(.width(width)) rd_st2_50  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[50]), .rdlo_in(a2_wr[178]),  .coef_in(coef[200]), .rdup_out(a3_wr[50]), .rdlo_out(a3_wr[178]));
			radix2 #(.width(width)) rd_st2_51  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[51]), .rdlo_in(a2_wr[179]),  .coef_in(coef[204]), .rdup_out(a3_wr[51]), .rdlo_out(a3_wr[179]));
			radix2 #(.width(width)) rd_st2_52  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[52]), .rdlo_in(a2_wr[180]),  .coef_in(coef[208]), .rdup_out(a3_wr[52]), .rdlo_out(a3_wr[180]));
			radix2 #(.width(width)) rd_st2_53  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[53]), .rdlo_in(a2_wr[181]),  .coef_in(coef[212]), .rdup_out(a3_wr[53]), .rdlo_out(a3_wr[181]));
			radix2 #(.width(width)) rd_st2_54  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[54]), .rdlo_in(a2_wr[182]),  .coef_in(coef[216]), .rdup_out(a3_wr[54]), .rdlo_out(a3_wr[182]));
			radix2 #(.width(width)) rd_st2_55  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[55]), .rdlo_in(a2_wr[183]),  .coef_in(coef[220]), .rdup_out(a3_wr[55]), .rdlo_out(a3_wr[183]));
			radix2 #(.width(width)) rd_st2_56  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[56]), .rdlo_in(a2_wr[184]),  .coef_in(coef[224]), .rdup_out(a3_wr[56]), .rdlo_out(a3_wr[184]));
			radix2 #(.width(width)) rd_st2_57  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[57]), .rdlo_in(a2_wr[185]),  .coef_in(coef[228]), .rdup_out(a3_wr[57]), .rdlo_out(a3_wr[185]));
			radix2 #(.width(width)) rd_st2_58  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[58]), .rdlo_in(a2_wr[186]),  .coef_in(coef[232]), .rdup_out(a3_wr[58]), .rdlo_out(a3_wr[186]));
			radix2 #(.width(width)) rd_st2_59  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[59]), .rdlo_in(a2_wr[187]),  .coef_in(coef[236]), .rdup_out(a3_wr[59]), .rdlo_out(a3_wr[187]));
			radix2 #(.width(width)) rd_st2_60  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[60]), .rdlo_in(a2_wr[188]),  .coef_in(coef[240]), .rdup_out(a3_wr[60]), .rdlo_out(a3_wr[188]));
			radix2 #(.width(width)) rd_st2_61  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[61]), .rdlo_in(a2_wr[189]),  .coef_in(coef[244]), .rdup_out(a3_wr[61]), .rdlo_out(a3_wr[189]));
			radix2 #(.width(width)) rd_st2_62  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[62]), .rdlo_in(a2_wr[190]),  .coef_in(coef[248]), .rdup_out(a3_wr[62]), .rdlo_out(a3_wr[190]));
			radix2 #(.width(width)) rd_st2_63  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[63]), .rdlo_in(a2_wr[191]),  .coef_in(coef[252]), .rdup_out(a3_wr[63]), .rdlo_out(a3_wr[191]));
			radix2 #(.width(width)) rd_st2_64  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[64]), .rdlo_in(a2_wr[192]),  .coef_in(coef[256]), .rdup_out(a3_wr[64]), .rdlo_out(a3_wr[192]));
			radix2 #(.width(width)) rd_st2_65  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[65]), .rdlo_in(a2_wr[193]),  .coef_in(coef[260]), .rdup_out(a3_wr[65]), .rdlo_out(a3_wr[193]));
			radix2 #(.width(width)) rd_st2_66  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[66]), .rdlo_in(a2_wr[194]),  .coef_in(coef[264]), .rdup_out(a3_wr[66]), .rdlo_out(a3_wr[194]));
			radix2 #(.width(width)) rd_st2_67  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[67]), .rdlo_in(a2_wr[195]),  .coef_in(coef[268]), .rdup_out(a3_wr[67]), .rdlo_out(a3_wr[195]));
			radix2 #(.width(width)) rd_st2_68  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[68]), .rdlo_in(a2_wr[196]),  .coef_in(coef[272]), .rdup_out(a3_wr[68]), .rdlo_out(a3_wr[196]));
			radix2 #(.width(width)) rd_st2_69  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[69]), .rdlo_in(a2_wr[197]),  .coef_in(coef[276]), .rdup_out(a3_wr[69]), .rdlo_out(a3_wr[197]));
			radix2 #(.width(width)) rd_st2_70  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[70]), .rdlo_in(a2_wr[198]),  .coef_in(coef[280]), .rdup_out(a3_wr[70]), .rdlo_out(a3_wr[198]));
			radix2 #(.width(width)) rd_st2_71  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[71]), .rdlo_in(a2_wr[199]),  .coef_in(coef[284]), .rdup_out(a3_wr[71]), .rdlo_out(a3_wr[199]));
			radix2 #(.width(width)) rd_st2_72  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[72]), .rdlo_in(a2_wr[200]),  .coef_in(coef[288]), .rdup_out(a3_wr[72]), .rdlo_out(a3_wr[200]));
			radix2 #(.width(width)) rd_st2_73  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[73]), .rdlo_in(a2_wr[201]),  .coef_in(coef[292]), .rdup_out(a3_wr[73]), .rdlo_out(a3_wr[201]));
			radix2 #(.width(width)) rd_st2_74  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[74]), .rdlo_in(a2_wr[202]),  .coef_in(coef[296]), .rdup_out(a3_wr[74]), .rdlo_out(a3_wr[202]));
			radix2 #(.width(width)) rd_st2_75  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[75]), .rdlo_in(a2_wr[203]),  .coef_in(coef[300]), .rdup_out(a3_wr[75]), .rdlo_out(a3_wr[203]));
			radix2 #(.width(width)) rd_st2_76  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[76]), .rdlo_in(a2_wr[204]),  .coef_in(coef[304]), .rdup_out(a3_wr[76]), .rdlo_out(a3_wr[204]));
			radix2 #(.width(width)) rd_st2_77  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[77]), .rdlo_in(a2_wr[205]),  .coef_in(coef[308]), .rdup_out(a3_wr[77]), .rdlo_out(a3_wr[205]));
			radix2 #(.width(width)) rd_st2_78  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[78]), .rdlo_in(a2_wr[206]),  .coef_in(coef[312]), .rdup_out(a3_wr[78]), .rdlo_out(a3_wr[206]));
			radix2 #(.width(width)) rd_st2_79  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[79]), .rdlo_in(a2_wr[207]),  .coef_in(coef[316]), .rdup_out(a3_wr[79]), .rdlo_out(a3_wr[207]));
			radix2 #(.width(width)) rd_st2_80  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[80]), .rdlo_in(a2_wr[208]),  .coef_in(coef[320]), .rdup_out(a3_wr[80]), .rdlo_out(a3_wr[208]));
			radix2 #(.width(width)) rd_st2_81  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[81]), .rdlo_in(a2_wr[209]),  .coef_in(coef[324]), .rdup_out(a3_wr[81]), .rdlo_out(a3_wr[209]));
			radix2 #(.width(width)) rd_st2_82  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[82]), .rdlo_in(a2_wr[210]),  .coef_in(coef[328]), .rdup_out(a3_wr[82]), .rdlo_out(a3_wr[210]));
			radix2 #(.width(width)) rd_st2_83  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[83]), .rdlo_in(a2_wr[211]),  .coef_in(coef[332]), .rdup_out(a3_wr[83]), .rdlo_out(a3_wr[211]));
			radix2 #(.width(width)) rd_st2_84  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[84]), .rdlo_in(a2_wr[212]),  .coef_in(coef[336]), .rdup_out(a3_wr[84]), .rdlo_out(a3_wr[212]));
			radix2 #(.width(width)) rd_st2_85  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[85]), .rdlo_in(a2_wr[213]),  .coef_in(coef[340]), .rdup_out(a3_wr[85]), .rdlo_out(a3_wr[213]));
			radix2 #(.width(width)) rd_st2_86  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[86]), .rdlo_in(a2_wr[214]),  .coef_in(coef[344]), .rdup_out(a3_wr[86]), .rdlo_out(a3_wr[214]));
			radix2 #(.width(width)) rd_st2_87  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[87]), .rdlo_in(a2_wr[215]),  .coef_in(coef[348]), .rdup_out(a3_wr[87]), .rdlo_out(a3_wr[215]));
			radix2 #(.width(width)) rd_st2_88  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[88]), .rdlo_in(a2_wr[216]),  .coef_in(coef[352]), .rdup_out(a3_wr[88]), .rdlo_out(a3_wr[216]));
			radix2 #(.width(width)) rd_st2_89  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[89]), .rdlo_in(a2_wr[217]),  .coef_in(coef[356]), .rdup_out(a3_wr[89]), .rdlo_out(a3_wr[217]));
			radix2 #(.width(width)) rd_st2_90  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[90]), .rdlo_in(a2_wr[218]),  .coef_in(coef[360]), .rdup_out(a3_wr[90]), .rdlo_out(a3_wr[218]));
			radix2 #(.width(width)) rd_st2_91  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[91]), .rdlo_in(a2_wr[219]),  .coef_in(coef[364]), .rdup_out(a3_wr[91]), .rdlo_out(a3_wr[219]));
			radix2 #(.width(width)) rd_st2_92  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[92]), .rdlo_in(a2_wr[220]),  .coef_in(coef[368]), .rdup_out(a3_wr[92]), .rdlo_out(a3_wr[220]));
			radix2 #(.width(width)) rd_st2_93  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[93]), .rdlo_in(a2_wr[221]),  .coef_in(coef[372]), .rdup_out(a3_wr[93]), .rdlo_out(a3_wr[221]));
			radix2 #(.width(width)) rd_st2_94  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[94]), .rdlo_in(a2_wr[222]),  .coef_in(coef[376]), .rdup_out(a3_wr[94]), .rdlo_out(a3_wr[222]));
			radix2 #(.width(width)) rd_st2_95  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[95]), .rdlo_in(a2_wr[223]),  .coef_in(coef[380]), .rdup_out(a3_wr[95]), .rdlo_out(a3_wr[223]));
			radix2 #(.width(width)) rd_st2_96  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[96]), .rdlo_in(a2_wr[224]),  .coef_in(coef[384]), .rdup_out(a3_wr[96]), .rdlo_out(a3_wr[224]));
			radix2 #(.width(width)) rd_st2_97  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[97]), .rdlo_in(a2_wr[225]),  .coef_in(coef[388]), .rdup_out(a3_wr[97]), .rdlo_out(a3_wr[225]));
			radix2 #(.width(width)) rd_st2_98  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[98]), .rdlo_in(a2_wr[226]),  .coef_in(coef[392]), .rdup_out(a3_wr[98]), .rdlo_out(a3_wr[226]));
			radix2 #(.width(width)) rd_st2_99  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[99]), .rdlo_in(a2_wr[227]),  .coef_in(coef[396]), .rdup_out(a3_wr[99]), .rdlo_out(a3_wr[227]));
			radix2 #(.width(width)) rd_st2_100  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[100]), .rdlo_in(a2_wr[228]),  .coef_in(coef[400]), .rdup_out(a3_wr[100]), .rdlo_out(a3_wr[228]));
			radix2 #(.width(width)) rd_st2_101  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[101]), .rdlo_in(a2_wr[229]),  .coef_in(coef[404]), .rdup_out(a3_wr[101]), .rdlo_out(a3_wr[229]));
			radix2 #(.width(width)) rd_st2_102  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[102]), .rdlo_in(a2_wr[230]),  .coef_in(coef[408]), .rdup_out(a3_wr[102]), .rdlo_out(a3_wr[230]));
			radix2 #(.width(width)) rd_st2_103  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[103]), .rdlo_in(a2_wr[231]),  .coef_in(coef[412]), .rdup_out(a3_wr[103]), .rdlo_out(a3_wr[231]));
			radix2 #(.width(width)) rd_st2_104  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[104]), .rdlo_in(a2_wr[232]),  .coef_in(coef[416]), .rdup_out(a3_wr[104]), .rdlo_out(a3_wr[232]));
			radix2 #(.width(width)) rd_st2_105  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[105]), .rdlo_in(a2_wr[233]),  .coef_in(coef[420]), .rdup_out(a3_wr[105]), .rdlo_out(a3_wr[233]));
			radix2 #(.width(width)) rd_st2_106  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[106]), .rdlo_in(a2_wr[234]),  .coef_in(coef[424]), .rdup_out(a3_wr[106]), .rdlo_out(a3_wr[234]));
			radix2 #(.width(width)) rd_st2_107  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[107]), .rdlo_in(a2_wr[235]),  .coef_in(coef[428]), .rdup_out(a3_wr[107]), .rdlo_out(a3_wr[235]));
			radix2 #(.width(width)) rd_st2_108  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[108]), .rdlo_in(a2_wr[236]),  .coef_in(coef[432]), .rdup_out(a3_wr[108]), .rdlo_out(a3_wr[236]));
			radix2 #(.width(width)) rd_st2_109  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[109]), .rdlo_in(a2_wr[237]),  .coef_in(coef[436]), .rdup_out(a3_wr[109]), .rdlo_out(a3_wr[237]));
			radix2 #(.width(width)) rd_st2_110  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[110]), .rdlo_in(a2_wr[238]),  .coef_in(coef[440]), .rdup_out(a3_wr[110]), .rdlo_out(a3_wr[238]));
			radix2 #(.width(width)) rd_st2_111  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[111]), .rdlo_in(a2_wr[239]),  .coef_in(coef[444]), .rdup_out(a3_wr[111]), .rdlo_out(a3_wr[239]));
			radix2 #(.width(width)) rd_st2_112  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[112]), .rdlo_in(a2_wr[240]),  .coef_in(coef[448]), .rdup_out(a3_wr[112]), .rdlo_out(a3_wr[240]));
			radix2 #(.width(width)) rd_st2_113  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[113]), .rdlo_in(a2_wr[241]),  .coef_in(coef[452]), .rdup_out(a3_wr[113]), .rdlo_out(a3_wr[241]));
			radix2 #(.width(width)) rd_st2_114  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[114]), .rdlo_in(a2_wr[242]),  .coef_in(coef[456]), .rdup_out(a3_wr[114]), .rdlo_out(a3_wr[242]));
			radix2 #(.width(width)) rd_st2_115  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[115]), .rdlo_in(a2_wr[243]),  .coef_in(coef[460]), .rdup_out(a3_wr[115]), .rdlo_out(a3_wr[243]));
			radix2 #(.width(width)) rd_st2_116  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[116]), .rdlo_in(a2_wr[244]),  .coef_in(coef[464]), .rdup_out(a3_wr[116]), .rdlo_out(a3_wr[244]));
			radix2 #(.width(width)) rd_st2_117  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[117]), .rdlo_in(a2_wr[245]),  .coef_in(coef[468]), .rdup_out(a3_wr[117]), .rdlo_out(a3_wr[245]));
			radix2 #(.width(width)) rd_st2_118  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[118]), .rdlo_in(a2_wr[246]),  .coef_in(coef[472]), .rdup_out(a3_wr[118]), .rdlo_out(a3_wr[246]));
			radix2 #(.width(width)) rd_st2_119  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[119]), .rdlo_in(a2_wr[247]),  .coef_in(coef[476]), .rdup_out(a3_wr[119]), .rdlo_out(a3_wr[247]));
			radix2 #(.width(width)) rd_st2_120  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[120]), .rdlo_in(a2_wr[248]),  .coef_in(coef[480]), .rdup_out(a3_wr[120]), .rdlo_out(a3_wr[248]));
			radix2 #(.width(width)) rd_st2_121  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[121]), .rdlo_in(a2_wr[249]),  .coef_in(coef[484]), .rdup_out(a3_wr[121]), .rdlo_out(a3_wr[249]));
			radix2 #(.width(width)) rd_st2_122  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[122]), .rdlo_in(a2_wr[250]),  .coef_in(coef[488]), .rdup_out(a3_wr[122]), .rdlo_out(a3_wr[250]));
			radix2 #(.width(width)) rd_st2_123  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[123]), .rdlo_in(a2_wr[251]),  .coef_in(coef[492]), .rdup_out(a3_wr[123]), .rdlo_out(a3_wr[251]));
			radix2 #(.width(width)) rd_st2_124  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[124]), .rdlo_in(a2_wr[252]),  .coef_in(coef[496]), .rdup_out(a3_wr[124]), .rdlo_out(a3_wr[252]));
			radix2 #(.width(width)) rd_st2_125  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[125]), .rdlo_in(a2_wr[253]),  .coef_in(coef[500]), .rdup_out(a3_wr[125]), .rdlo_out(a3_wr[253]));
			radix2 #(.width(width)) rd_st2_126  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[126]), .rdlo_in(a2_wr[254]),  .coef_in(coef[504]), .rdup_out(a3_wr[126]), .rdlo_out(a3_wr[254]));
			radix2 #(.width(width)) rd_st2_127  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[127]), .rdlo_in(a2_wr[255]),  .coef_in(coef[508]), .rdup_out(a3_wr[127]), .rdlo_out(a3_wr[255]));
			radix2 #(.width(width)) rd_st2_256  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[256]), .rdlo_in(a2_wr[384]),  .coef_in(coef[0]), .rdup_out(a3_wr[256]), .rdlo_out(a3_wr[384]));
			radix2 #(.width(width)) rd_st2_257  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[257]), .rdlo_in(a2_wr[385]),  .coef_in(coef[4]), .rdup_out(a3_wr[257]), .rdlo_out(a3_wr[385]));
			radix2 #(.width(width)) rd_st2_258  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[258]), .rdlo_in(a2_wr[386]),  .coef_in(coef[8]), .rdup_out(a3_wr[258]), .rdlo_out(a3_wr[386]));
			radix2 #(.width(width)) rd_st2_259  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[259]), .rdlo_in(a2_wr[387]),  .coef_in(coef[12]), .rdup_out(a3_wr[259]), .rdlo_out(a3_wr[387]));
			radix2 #(.width(width)) rd_st2_260  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[260]), .rdlo_in(a2_wr[388]),  .coef_in(coef[16]), .rdup_out(a3_wr[260]), .rdlo_out(a3_wr[388]));
			radix2 #(.width(width)) rd_st2_261  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[261]), .rdlo_in(a2_wr[389]),  .coef_in(coef[20]), .rdup_out(a3_wr[261]), .rdlo_out(a3_wr[389]));
			radix2 #(.width(width)) rd_st2_262  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[262]), .rdlo_in(a2_wr[390]),  .coef_in(coef[24]), .rdup_out(a3_wr[262]), .rdlo_out(a3_wr[390]));
			radix2 #(.width(width)) rd_st2_263  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[263]), .rdlo_in(a2_wr[391]),  .coef_in(coef[28]), .rdup_out(a3_wr[263]), .rdlo_out(a3_wr[391]));
			radix2 #(.width(width)) rd_st2_264  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[264]), .rdlo_in(a2_wr[392]),  .coef_in(coef[32]), .rdup_out(a3_wr[264]), .rdlo_out(a3_wr[392]));
			radix2 #(.width(width)) rd_st2_265  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[265]), .rdlo_in(a2_wr[393]),  .coef_in(coef[36]), .rdup_out(a3_wr[265]), .rdlo_out(a3_wr[393]));
			radix2 #(.width(width)) rd_st2_266  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[266]), .rdlo_in(a2_wr[394]),  .coef_in(coef[40]), .rdup_out(a3_wr[266]), .rdlo_out(a3_wr[394]));
			radix2 #(.width(width)) rd_st2_267  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[267]), .rdlo_in(a2_wr[395]),  .coef_in(coef[44]), .rdup_out(a3_wr[267]), .rdlo_out(a3_wr[395]));
			radix2 #(.width(width)) rd_st2_268  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[268]), .rdlo_in(a2_wr[396]),  .coef_in(coef[48]), .rdup_out(a3_wr[268]), .rdlo_out(a3_wr[396]));
			radix2 #(.width(width)) rd_st2_269  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[269]), .rdlo_in(a2_wr[397]),  .coef_in(coef[52]), .rdup_out(a3_wr[269]), .rdlo_out(a3_wr[397]));
			radix2 #(.width(width)) rd_st2_270  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[270]), .rdlo_in(a2_wr[398]),  .coef_in(coef[56]), .rdup_out(a3_wr[270]), .rdlo_out(a3_wr[398]));
			radix2 #(.width(width)) rd_st2_271  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[271]), .rdlo_in(a2_wr[399]),  .coef_in(coef[60]), .rdup_out(a3_wr[271]), .rdlo_out(a3_wr[399]));
			radix2 #(.width(width)) rd_st2_272  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[272]), .rdlo_in(a2_wr[400]),  .coef_in(coef[64]), .rdup_out(a3_wr[272]), .rdlo_out(a3_wr[400]));
			radix2 #(.width(width)) rd_st2_273  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[273]), .rdlo_in(a2_wr[401]),  .coef_in(coef[68]), .rdup_out(a3_wr[273]), .rdlo_out(a3_wr[401]));
			radix2 #(.width(width)) rd_st2_274  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[274]), .rdlo_in(a2_wr[402]),  .coef_in(coef[72]), .rdup_out(a3_wr[274]), .rdlo_out(a3_wr[402]));
			radix2 #(.width(width)) rd_st2_275  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[275]), .rdlo_in(a2_wr[403]),  .coef_in(coef[76]), .rdup_out(a3_wr[275]), .rdlo_out(a3_wr[403]));
			radix2 #(.width(width)) rd_st2_276  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[276]), .rdlo_in(a2_wr[404]),  .coef_in(coef[80]), .rdup_out(a3_wr[276]), .rdlo_out(a3_wr[404]));
			radix2 #(.width(width)) rd_st2_277  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[277]), .rdlo_in(a2_wr[405]),  .coef_in(coef[84]), .rdup_out(a3_wr[277]), .rdlo_out(a3_wr[405]));
			radix2 #(.width(width)) rd_st2_278  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[278]), .rdlo_in(a2_wr[406]),  .coef_in(coef[88]), .rdup_out(a3_wr[278]), .rdlo_out(a3_wr[406]));
			radix2 #(.width(width)) rd_st2_279  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[279]), .rdlo_in(a2_wr[407]),  .coef_in(coef[92]), .rdup_out(a3_wr[279]), .rdlo_out(a3_wr[407]));
			radix2 #(.width(width)) rd_st2_280  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[280]), .rdlo_in(a2_wr[408]),  .coef_in(coef[96]), .rdup_out(a3_wr[280]), .rdlo_out(a3_wr[408]));
			radix2 #(.width(width)) rd_st2_281  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[281]), .rdlo_in(a2_wr[409]),  .coef_in(coef[100]), .rdup_out(a3_wr[281]), .rdlo_out(a3_wr[409]));
			radix2 #(.width(width)) rd_st2_282  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[282]), .rdlo_in(a2_wr[410]),  .coef_in(coef[104]), .rdup_out(a3_wr[282]), .rdlo_out(a3_wr[410]));
			radix2 #(.width(width)) rd_st2_283  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[283]), .rdlo_in(a2_wr[411]),  .coef_in(coef[108]), .rdup_out(a3_wr[283]), .rdlo_out(a3_wr[411]));
			radix2 #(.width(width)) rd_st2_284  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[284]), .rdlo_in(a2_wr[412]),  .coef_in(coef[112]), .rdup_out(a3_wr[284]), .rdlo_out(a3_wr[412]));
			radix2 #(.width(width)) rd_st2_285  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[285]), .rdlo_in(a2_wr[413]),  .coef_in(coef[116]), .rdup_out(a3_wr[285]), .rdlo_out(a3_wr[413]));
			radix2 #(.width(width)) rd_st2_286  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[286]), .rdlo_in(a2_wr[414]),  .coef_in(coef[120]), .rdup_out(a3_wr[286]), .rdlo_out(a3_wr[414]));
			radix2 #(.width(width)) rd_st2_287  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[287]), .rdlo_in(a2_wr[415]),  .coef_in(coef[124]), .rdup_out(a3_wr[287]), .rdlo_out(a3_wr[415]));
			radix2 #(.width(width)) rd_st2_288  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[288]), .rdlo_in(a2_wr[416]),  .coef_in(coef[128]), .rdup_out(a3_wr[288]), .rdlo_out(a3_wr[416]));
			radix2 #(.width(width)) rd_st2_289  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[289]), .rdlo_in(a2_wr[417]),  .coef_in(coef[132]), .rdup_out(a3_wr[289]), .rdlo_out(a3_wr[417]));
			radix2 #(.width(width)) rd_st2_290  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[290]), .rdlo_in(a2_wr[418]),  .coef_in(coef[136]), .rdup_out(a3_wr[290]), .rdlo_out(a3_wr[418]));
			radix2 #(.width(width)) rd_st2_291  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[291]), .rdlo_in(a2_wr[419]),  .coef_in(coef[140]), .rdup_out(a3_wr[291]), .rdlo_out(a3_wr[419]));
			radix2 #(.width(width)) rd_st2_292  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[292]), .rdlo_in(a2_wr[420]),  .coef_in(coef[144]), .rdup_out(a3_wr[292]), .rdlo_out(a3_wr[420]));
			radix2 #(.width(width)) rd_st2_293  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[293]), .rdlo_in(a2_wr[421]),  .coef_in(coef[148]), .rdup_out(a3_wr[293]), .rdlo_out(a3_wr[421]));
			radix2 #(.width(width)) rd_st2_294  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[294]), .rdlo_in(a2_wr[422]),  .coef_in(coef[152]), .rdup_out(a3_wr[294]), .rdlo_out(a3_wr[422]));
			radix2 #(.width(width)) rd_st2_295  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[295]), .rdlo_in(a2_wr[423]),  .coef_in(coef[156]), .rdup_out(a3_wr[295]), .rdlo_out(a3_wr[423]));
			radix2 #(.width(width)) rd_st2_296  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[296]), .rdlo_in(a2_wr[424]),  .coef_in(coef[160]), .rdup_out(a3_wr[296]), .rdlo_out(a3_wr[424]));
			radix2 #(.width(width)) rd_st2_297  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[297]), .rdlo_in(a2_wr[425]),  .coef_in(coef[164]), .rdup_out(a3_wr[297]), .rdlo_out(a3_wr[425]));
			radix2 #(.width(width)) rd_st2_298  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[298]), .rdlo_in(a2_wr[426]),  .coef_in(coef[168]), .rdup_out(a3_wr[298]), .rdlo_out(a3_wr[426]));
			radix2 #(.width(width)) rd_st2_299  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[299]), .rdlo_in(a2_wr[427]),  .coef_in(coef[172]), .rdup_out(a3_wr[299]), .rdlo_out(a3_wr[427]));
			radix2 #(.width(width)) rd_st2_300  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[300]), .rdlo_in(a2_wr[428]),  .coef_in(coef[176]), .rdup_out(a3_wr[300]), .rdlo_out(a3_wr[428]));
			radix2 #(.width(width)) rd_st2_301  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[301]), .rdlo_in(a2_wr[429]),  .coef_in(coef[180]), .rdup_out(a3_wr[301]), .rdlo_out(a3_wr[429]));
			radix2 #(.width(width)) rd_st2_302  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[302]), .rdlo_in(a2_wr[430]),  .coef_in(coef[184]), .rdup_out(a3_wr[302]), .rdlo_out(a3_wr[430]));
			radix2 #(.width(width)) rd_st2_303  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[303]), .rdlo_in(a2_wr[431]),  .coef_in(coef[188]), .rdup_out(a3_wr[303]), .rdlo_out(a3_wr[431]));
			radix2 #(.width(width)) rd_st2_304  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[304]), .rdlo_in(a2_wr[432]),  .coef_in(coef[192]), .rdup_out(a3_wr[304]), .rdlo_out(a3_wr[432]));
			radix2 #(.width(width)) rd_st2_305  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[305]), .rdlo_in(a2_wr[433]),  .coef_in(coef[196]), .rdup_out(a3_wr[305]), .rdlo_out(a3_wr[433]));
			radix2 #(.width(width)) rd_st2_306  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[306]), .rdlo_in(a2_wr[434]),  .coef_in(coef[200]), .rdup_out(a3_wr[306]), .rdlo_out(a3_wr[434]));
			radix2 #(.width(width)) rd_st2_307  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[307]), .rdlo_in(a2_wr[435]),  .coef_in(coef[204]), .rdup_out(a3_wr[307]), .rdlo_out(a3_wr[435]));
			radix2 #(.width(width)) rd_st2_308  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[308]), .rdlo_in(a2_wr[436]),  .coef_in(coef[208]), .rdup_out(a3_wr[308]), .rdlo_out(a3_wr[436]));
			radix2 #(.width(width)) rd_st2_309  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[309]), .rdlo_in(a2_wr[437]),  .coef_in(coef[212]), .rdup_out(a3_wr[309]), .rdlo_out(a3_wr[437]));
			radix2 #(.width(width)) rd_st2_310  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[310]), .rdlo_in(a2_wr[438]),  .coef_in(coef[216]), .rdup_out(a3_wr[310]), .rdlo_out(a3_wr[438]));
			radix2 #(.width(width)) rd_st2_311  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[311]), .rdlo_in(a2_wr[439]),  .coef_in(coef[220]), .rdup_out(a3_wr[311]), .rdlo_out(a3_wr[439]));
			radix2 #(.width(width)) rd_st2_312  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[312]), .rdlo_in(a2_wr[440]),  .coef_in(coef[224]), .rdup_out(a3_wr[312]), .rdlo_out(a3_wr[440]));
			radix2 #(.width(width)) rd_st2_313  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[313]), .rdlo_in(a2_wr[441]),  .coef_in(coef[228]), .rdup_out(a3_wr[313]), .rdlo_out(a3_wr[441]));
			radix2 #(.width(width)) rd_st2_314  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[314]), .rdlo_in(a2_wr[442]),  .coef_in(coef[232]), .rdup_out(a3_wr[314]), .rdlo_out(a3_wr[442]));
			radix2 #(.width(width)) rd_st2_315  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[315]), .rdlo_in(a2_wr[443]),  .coef_in(coef[236]), .rdup_out(a3_wr[315]), .rdlo_out(a3_wr[443]));
			radix2 #(.width(width)) rd_st2_316  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[316]), .rdlo_in(a2_wr[444]),  .coef_in(coef[240]), .rdup_out(a3_wr[316]), .rdlo_out(a3_wr[444]));
			radix2 #(.width(width)) rd_st2_317  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[317]), .rdlo_in(a2_wr[445]),  .coef_in(coef[244]), .rdup_out(a3_wr[317]), .rdlo_out(a3_wr[445]));
			radix2 #(.width(width)) rd_st2_318  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[318]), .rdlo_in(a2_wr[446]),  .coef_in(coef[248]), .rdup_out(a3_wr[318]), .rdlo_out(a3_wr[446]));
			radix2 #(.width(width)) rd_st2_319  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[319]), .rdlo_in(a2_wr[447]),  .coef_in(coef[252]), .rdup_out(a3_wr[319]), .rdlo_out(a3_wr[447]));
			radix2 #(.width(width)) rd_st2_320  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[320]), .rdlo_in(a2_wr[448]),  .coef_in(coef[256]), .rdup_out(a3_wr[320]), .rdlo_out(a3_wr[448]));
			radix2 #(.width(width)) rd_st2_321  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[321]), .rdlo_in(a2_wr[449]),  .coef_in(coef[260]), .rdup_out(a3_wr[321]), .rdlo_out(a3_wr[449]));
			radix2 #(.width(width)) rd_st2_322  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[322]), .rdlo_in(a2_wr[450]),  .coef_in(coef[264]), .rdup_out(a3_wr[322]), .rdlo_out(a3_wr[450]));
			radix2 #(.width(width)) rd_st2_323  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[323]), .rdlo_in(a2_wr[451]),  .coef_in(coef[268]), .rdup_out(a3_wr[323]), .rdlo_out(a3_wr[451]));
			radix2 #(.width(width)) rd_st2_324  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[324]), .rdlo_in(a2_wr[452]),  .coef_in(coef[272]), .rdup_out(a3_wr[324]), .rdlo_out(a3_wr[452]));
			radix2 #(.width(width)) rd_st2_325  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[325]), .rdlo_in(a2_wr[453]),  .coef_in(coef[276]), .rdup_out(a3_wr[325]), .rdlo_out(a3_wr[453]));
			radix2 #(.width(width)) rd_st2_326  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[326]), .rdlo_in(a2_wr[454]),  .coef_in(coef[280]), .rdup_out(a3_wr[326]), .rdlo_out(a3_wr[454]));
			radix2 #(.width(width)) rd_st2_327  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[327]), .rdlo_in(a2_wr[455]),  .coef_in(coef[284]), .rdup_out(a3_wr[327]), .rdlo_out(a3_wr[455]));
			radix2 #(.width(width)) rd_st2_328  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[328]), .rdlo_in(a2_wr[456]),  .coef_in(coef[288]), .rdup_out(a3_wr[328]), .rdlo_out(a3_wr[456]));
			radix2 #(.width(width)) rd_st2_329  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[329]), .rdlo_in(a2_wr[457]),  .coef_in(coef[292]), .rdup_out(a3_wr[329]), .rdlo_out(a3_wr[457]));
			radix2 #(.width(width)) rd_st2_330  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[330]), .rdlo_in(a2_wr[458]),  .coef_in(coef[296]), .rdup_out(a3_wr[330]), .rdlo_out(a3_wr[458]));
			radix2 #(.width(width)) rd_st2_331  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[331]), .rdlo_in(a2_wr[459]),  .coef_in(coef[300]), .rdup_out(a3_wr[331]), .rdlo_out(a3_wr[459]));
			radix2 #(.width(width)) rd_st2_332  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[332]), .rdlo_in(a2_wr[460]),  .coef_in(coef[304]), .rdup_out(a3_wr[332]), .rdlo_out(a3_wr[460]));
			radix2 #(.width(width)) rd_st2_333  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[333]), .rdlo_in(a2_wr[461]),  .coef_in(coef[308]), .rdup_out(a3_wr[333]), .rdlo_out(a3_wr[461]));
			radix2 #(.width(width)) rd_st2_334  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[334]), .rdlo_in(a2_wr[462]),  .coef_in(coef[312]), .rdup_out(a3_wr[334]), .rdlo_out(a3_wr[462]));
			radix2 #(.width(width)) rd_st2_335  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[335]), .rdlo_in(a2_wr[463]),  .coef_in(coef[316]), .rdup_out(a3_wr[335]), .rdlo_out(a3_wr[463]));
			radix2 #(.width(width)) rd_st2_336  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[336]), .rdlo_in(a2_wr[464]),  .coef_in(coef[320]), .rdup_out(a3_wr[336]), .rdlo_out(a3_wr[464]));
			radix2 #(.width(width)) rd_st2_337  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[337]), .rdlo_in(a2_wr[465]),  .coef_in(coef[324]), .rdup_out(a3_wr[337]), .rdlo_out(a3_wr[465]));
			radix2 #(.width(width)) rd_st2_338  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[338]), .rdlo_in(a2_wr[466]),  .coef_in(coef[328]), .rdup_out(a3_wr[338]), .rdlo_out(a3_wr[466]));
			radix2 #(.width(width)) rd_st2_339  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[339]), .rdlo_in(a2_wr[467]),  .coef_in(coef[332]), .rdup_out(a3_wr[339]), .rdlo_out(a3_wr[467]));
			radix2 #(.width(width)) rd_st2_340  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[340]), .rdlo_in(a2_wr[468]),  .coef_in(coef[336]), .rdup_out(a3_wr[340]), .rdlo_out(a3_wr[468]));
			radix2 #(.width(width)) rd_st2_341  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[341]), .rdlo_in(a2_wr[469]),  .coef_in(coef[340]), .rdup_out(a3_wr[341]), .rdlo_out(a3_wr[469]));
			radix2 #(.width(width)) rd_st2_342  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[342]), .rdlo_in(a2_wr[470]),  .coef_in(coef[344]), .rdup_out(a3_wr[342]), .rdlo_out(a3_wr[470]));
			radix2 #(.width(width)) rd_st2_343  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[343]), .rdlo_in(a2_wr[471]),  .coef_in(coef[348]), .rdup_out(a3_wr[343]), .rdlo_out(a3_wr[471]));
			radix2 #(.width(width)) rd_st2_344  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[344]), .rdlo_in(a2_wr[472]),  .coef_in(coef[352]), .rdup_out(a3_wr[344]), .rdlo_out(a3_wr[472]));
			radix2 #(.width(width)) rd_st2_345  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[345]), .rdlo_in(a2_wr[473]),  .coef_in(coef[356]), .rdup_out(a3_wr[345]), .rdlo_out(a3_wr[473]));
			radix2 #(.width(width)) rd_st2_346  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[346]), .rdlo_in(a2_wr[474]),  .coef_in(coef[360]), .rdup_out(a3_wr[346]), .rdlo_out(a3_wr[474]));
			radix2 #(.width(width)) rd_st2_347  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[347]), .rdlo_in(a2_wr[475]),  .coef_in(coef[364]), .rdup_out(a3_wr[347]), .rdlo_out(a3_wr[475]));
			radix2 #(.width(width)) rd_st2_348  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[348]), .rdlo_in(a2_wr[476]),  .coef_in(coef[368]), .rdup_out(a3_wr[348]), .rdlo_out(a3_wr[476]));
			radix2 #(.width(width)) rd_st2_349  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[349]), .rdlo_in(a2_wr[477]),  .coef_in(coef[372]), .rdup_out(a3_wr[349]), .rdlo_out(a3_wr[477]));
			radix2 #(.width(width)) rd_st2_350  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[350]), .rdlo_in(a2_wr[478]),  .coef_in(coef[376]), .rdup_out(a3_wr[350]), .rdlo_out(a3_wr[478]));
			radix2 #(.width(width)) rd_st2_351  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[351]), .rdlo_in(a2_wr[479]),  .coef_in(coef[380]), .rdup_out(a3_wr[351]), .rdlo_out(a3_wr[479]));
			radix2 #(.width(width)) rd_st2_352  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[352]), .rdlo_in(a2_wr[480]),  .coef_in(coef[384]), .rdup_out(a3_wr[352]), .rdlo_out(a3_wr[480]));
			radix2 #(.width(width)) rd_st2_353  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[353]), .rdlo_in(a2_wr[481]),  .coef_in(coef[388]), .rdup_out(a3_wr[353]), .rdlo_out(a3_wr[481]));
			radix2 #(.width(width)) rd_st2_354  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[354]), .rdlo_in(a2_wr[482]),  .coef_in(coef[392]), .rdup_out(a3_wr[354]), .rdlo_out(a3_wr[482]));
			radix2 #(.width(width)) rd_st2_355  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[355]), .rdlo_in(a2_wr[483]),  .coef_in(coef[396]), .rdup_out(a3_wr[355]), .rdlo_out(a3_wr[483]));
			radix2 #(.width(width)) rd_st2_356  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[356]), .rdlo_in(a2_wr[484]),  .coef_in(coef[400]), .rdup_out(a3_wr[356]), .rdlo_out(a3_wr[484]));
			radix2 #(.width(width)) rd_st2_357  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[357]), .rdlo_in(a2_wr[485]),  .coef_in(coef[404]), .rdup_out(a3_wr[357]), .rdlo_out(a3_wr[485]));
			radix2 #(.width(width)) rd_st2_358  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[358]), .rdlo_in(a2_wr[486]),  .coef_in(coef[408]), .rdup_out(a3_wr[358]), .rdlo_out(a3_wr[486]));
			radix2 #(.width(width)) rd_st2_359  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[359]), .rdlo_in(a2_wr[487]),  .coef_in(coef[412]), .rdup_out(a3_wr[359]), .rdlo_out(a3_wr[487]));
			radix2 #(.width(width)) rd_st2_360  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[360]), .rdlo_in(a2_wr[488]),  .coef_in(coef[416]), .rdup_out(a3_wr[360]), .rdlo_out(a3_wr[488]));
			radix2 #(.width(width)) rd_st2_361  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[361]), .rdlo_in(a2_wr[489]),  .coef_in(coef[420]), .rdup_out(a3_wr[361]), .rdlo_out(a3_wr[489]));
			radix2 #(.width(width)) rd_st2_362  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[362]), .rdlo_in(a2_wr[490]),  .coef_in(coef[424]), .rdup_out(a3_wr[362]), .rdlo_out(a3_wr[490]));
			radix2 #(.width(width)) rd_st2_363  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[363]), .rdlo_in(a2_wr[491]),  .coef_in(coef[428]), .rdup_out(a3_wr[363]), .rdlo_out(a3_wr[491]));
			radix2 #(.width(width)) rd_st2_364  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[364]), .rdlo_in(a2_wr[492]),  .coef_in(coef[432]), .rdup_out(a3_wr[364]), .rdlo_out(a3_wr[492]));
			radix2 #(.width(width)) rd_st2_365  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[365]), .rdlo_in(a2_wr[493]),  .coef_in(coef[436]), .rdup_out(a3_wr[365]), .rdlo_out(a3_wr[493]));
			radix2 #(.width(width)) rd_st2_366  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[366]), .rdlo_in(a2_wr[494]),  .coef_in(coef[440]), .rdup_out(a3_wr[366]), .rdlo_out(a3_wr[494]));
			radix2 #(.width(width)) rd_st2_367  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[367]), .rdlo_in(a2_wr[495]),  .coef_in(coef[444]), .rdup_out(a3_wr[367]), .rdlo_out(a3_wr[495]));
			radix2 #(.width(width)) rd_st2_368  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[368]), .rdlo_in(a2_wr[496]),  .coef_in(coef[448]), .rdup_out(a3_wr[368]), .rdlo_out(a3_wr[496]));
			radix2 #(.width(width)) rd_st2_369  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[369]), .rdlo_in(a2_wr[497]),  .coef_in(coef[452]), .rdup_out(a3_wr[369]), .rdlo_out(a3_wr[497]));
			radix2 #(.width(width)) rd_st2_370  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[370]), .rdlo_in(a2_wr[498]),  .coef_in(coef[456]), .rdup_out(a3_wr[370]), .rdlo_out(a3_wr[498]));
			radix2 #(.width(width)) rd_st2_371  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[371]), .rdlo_in(a2_wr[499]),  .coef_in(coef[460]), .rdup_out(a3_wr[371]), .rdlo_out(a3_wr[499]));
			radix2 #(.width(width)) rd_st2_372  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[372]), .rdlo_in(a2_wr[500]),  .coef_in(coef[464]), .rdup_out(a3_wr[372]), .rdlo_out(a3_wr[500]));
			radix2 #(.width(width)) rd_st2_373  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[373]), .rdlo_in(a2_wr[501]),  .coef_in(coef[468]), .rdup_out(a3_wr[373]), .rdlo_out(a3_wr[501]));
			radix2 #(.width(width)) rd_st2_374  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[374]), .rdlo_in(a2_wr[502]),  .coef_in(coef[472]), .rdup_out(a3_wr[374]), .rdlo_out(a3_wr[502]));
			radix2 #(.width(width)) rd_st2_375  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[375]), .rdlo_in(a2_wr[503]),  .coef_in(coef[476]), .rdup_out(a3_wr[375]), .rdlo_out(a3_wr[503]));
			radix2 #(.width(width)) rd_st2_376  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[376]), .rdlo_in(a2_wr[504]),  .coef_in(coef[480]), .rdup_out(a3_wr[376]), .rdlo_out(a3_wr[504]));
			radix2 #(.width(width)) rd_st2_377  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[377]), .rdlo_in(a2_wr[505]),  .coef_in(coef[484]), .rdup_out(a3_wr[377]), .rdlo_out(a3_wr[505]));
			radix2 #(.width(width)) rd_st2_378  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[378]), .rdlo_in(a2_wr[506]),  .coef_in(coef[488]), .rdup_out(a3_wr[378]), .rdlo_out(a3_wr[506]));
			radix2 #(.width(width)) rd_st2_379  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[379]), .rdlo_in(a2_wr[507]),  .coef_in(coef[492]), .rdup_out(a3_wr[379]), .rdlo_out(a3_wr[507]));
			radix2 #(.width(width)) rd_st2_380  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[380]), .rdlo_in(a2_wr[508]),  .coef_in(coef[496]), .rdup_out(a3_wr[380]), .rdlo_out(a3_wr[508]));
			radix2 #(.width(width)) rd_st2_381  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[381]), .rdlo_in(a2_wr[509]),  .coef_in(coef[500]), .rdup_out(a3_wr[381]), .rdlo_out(a3_wr[509]));
			radix2 #(.width(width)) rd_st2_382  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[382]), .rdlo_in(a2_wr[510]),  .coef_in(coef[504]), .rdup_out(a3_wr[382]), .rdlo_out(a3_wr[510]));
			radix2 #(.width(width)) rd_st2_383  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[383]), .rdlo_in(a2_wr[511]),  .coef_in(coef[508]), .rdup_out(a3_wr[383]), .rdlo_out(a3_wr[511]));
			radix2 #(.width(width)) rd_st2_512  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[512]), .rdlo_in(a2_wr[640]),  .coef_in(coef[0]), .rdup_out(a3_wr[512]), .rdlo_out(a3_wr[640]));
			radix2 #(.width(width)) rd_st2_513  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[513]), .rdlo_in(a2_wr[641]),  .coef_in(coef[4]), .rdup_out(a3_wr[513]), .rdlo_out(a3_wr[641]));
			radix2 #(.width(width)) rd_st2_514  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[514]), .rdlo_in(a2_wr[642]),  .coef_in(coef[8]), .rdup_out(a3_wr[514]), .rdlo_out(a3_wr[642]));
			radix2 #(.width(width)) rd_st2_515  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[515]), .rdlo_in(a2_wr[643]),  .coef_in(coef[12]), .rdup_out(a3_wr[515]), .rdlo_out(a3_wr[643]));
			radix2 #(.width(width)) rd_st2_516  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[516]), .rdlo_in(a2_wr[644]),  .coef_in(coef[16]), .rdup_out(a3_wr[516]), .rdlo_out(a3_wr[644]));
			radix2 #(.width(width)) rd_st2_517  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[517]), .rdlo_in(a2_wr[645]),  .coef_in(coef[20]), .rdup_out(a3_wr[517]), .rdlo_out(a3_wr[645]));
			radix2 #(.width(width)) rd_st2_518  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[518]), .rdlo_in(a2_wr[646]),  .coef_in(coef[24]), .rdup_out(a3_wr[518]), .rdlo_out(a3_wr[646]));
			radix2 #(.width(width)) rd_st2_519  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[519]), .rdlo_in(a2_wr[647]),  .coef_in(coef[28]), .rdup_out(a3_wr[519]), .rdlo_out(a3_wr[647]));
			radix2 #(.width(width)) rd_st2_520  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[520]), .rdlo_in(a2_wr[648]),  .coef_in(coef[32]), .rdup_out(a3_wr[520]), .rdlo_out(a3_wr[648]));
			radix2 #(.width(width)) rd_st2_521  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[521]), .rdlo_in(a2_wr[649]),  .coef_in(coef[36]), .rdup_out(a3_wr[521]), .rdlo_out(a3_wr[649]));
			radix2 #(.width(width)) rd_st2_522  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[522]), .rdlo_in(a2_wr[650]),  .coef_in(coef[40]), .rdup_out(a3_wr[522]), .rdlo_out(a3_wr[650]));
			radix2 #(.width(width)) rd_st2_523  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[523]), .rdlo_in(a2_wr[651]),  .coef_in(coef[44]), .rdup_out(a3_wr[523]), .rdlo_out(a3_wr[651]));
			radix2 #(.width(width)) rd_st2_524  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[524]), .rdlo_in(a2_wr[652]),  .coef_in(coef[48]), .rdup_out(a3_wr[524]), .rdlo_out(a3_wr[652]));
			radix2 #(.width(width)) rd_st2_525  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[525]), .rdlo_in(a2_wr[653]),  .coef_in(coef[52]), .rdup_out(a3_wr[525]), .rdlo_out(a3_wr[653]));
			radix2 #(.width(width)) rd_st2_526  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[526]), .rdlo_in(a2_wr[654]),  .coef_in(coef[56]), .rdup_out(a3_wr[526]), .rdlo_out(a3_wr[654]));
			radix2 #(.width(width)) rd_st2_527  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[527]), .rdlo_in(a2_wr[655]),  .coef_in(coef[60]), .rdup_out(a3_wr[527]), .rdlo_out(a3_wr[655]));
			radix2 #(.width(width)) rd_st2_528  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[528]), .rdlo_in(a2_wr[656]),  .coef_in(coef[64]), .rdup_out(a3_wr[528]), .rdlo_out(a3_wr[656]));
			radix2 #(.width(width)) rd_st2_529  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[529]), .rdlo_in(a2_wr[657]),  .coef_in(coef[68]), .rdup_out(a3_wr[529]), .rdlo_out(a3_wr[657]));
			radix2 #(.width(width)) rd_st2_530  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[530]), .rdlo_in(a2_wr[658]),  .coef_in(coef[72]), .rdup_out(a3_wr[530]), .rdlo_out(a3_wr[658]));
			radix2 #(.width(width)) rd_st2_531  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[531]), .rdlo_in(a2_wr[659]),  .coef_in(coef[76]), .rdup_out(a3_wr[531]), .rdlo_out(a3_wr[659]));
			radix2 #(.width(width)) rd_st2_532  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[532]), .rdlo_in(a2_wr[660]),  .coef_in(coef[80]), .rdup_out(a3_wr[532]), .rdlo_out(a3_wr[660]));
			radix2 #(.width(width)) rd_st2_533  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[533]), .rdlo_in(a2_wr[661]),  .coef_in(coef[84]), .rdup_out(a3_wr[533]), .rdlo_out(a3_wr[661]));
			radix2 #(.width(width)) rd_st2_534  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[534]), .rdlo_in(a2_wr[662]),  .coef_in(coef[88]), .rdup_out(a3_wr[534]), .rdlo_out(a3_wr[662]));
			radix2 #(.width(width)) rd_st2_535  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[535]), .rdlo_in(a2_wr[663]),  .coef_in(coef[92]), .rdup_out(a3_wr[535]), .rdlo_out(a3_wr[663]));
			radix2 #(.width(width)) rd_st2_536  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[536]), .rdlo_in(a2_wr[664]),  .coef_in(coef[96]), .rdup_out(a3_wr[536]), .rdlo_out(a3_wr[664]));
			radix2 #(.width(width)) rd_st2_537  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[537]), .rdlo_in(a2_wr[665]),  .coef_in(coef[100]), .rdup_out(a3_wr[537]), .rdlo_out(a3_wr[665]));
			radix2 #(.width(width)) rd_st2_538  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[538]), .rdlo_in(a2_wr[666]),  .coef_in(coef[104]), .rdup_out(a3_wr[538]), .rdlo_out(a3_wr[666]));
			radix2 #(.width(width)) rd_st2_539  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[539]), .rdlo_in(a2_wr[667]),  .coef_in(coef[108]), .rdup_out(a3_wr[539]), .rdlo_out(a3_wr[667]));
			radix2 #(.width(width)) rd_st2_540  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[540]), .rdlo_in(a2_wr[668]),  .coef_in(coef[112]), .rdup_out(a3_wr[540]), .rdlo_out(a3_wr[668]));
			radix2 #(.width(width)) rd_st2_541  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[541]), .rdlo_in(a2_wr[669]),  .coef_in(coef[116]), .rdup_out(a3_wr[541]), .rdlo_out(a3_wr[669]));
			radix2 #(.width(width)) rd_st2_542  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[542]), .rdlo_in(a2_wr[670]),  .coef_in(coef[120]), .rdup_out(a3_wr[542]), .rdlo_out(a3_wr[670]));
			radix2 #(.width(width)) rd_st2_543  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[543]), .rdlo_in(a2_wr[671]),  .coef_in(coef[124]), .rdup_out(a3_wr[543]), .rdlo_out(a3_wr[671]));
			radix2 #(.width(width)) rd_st2_544  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[544]), .rdlo_in(a2_wr[672]),  .coef_in(coef[128]), .rdup_out(a3_wr[544]), .rdlo_out(a3_wr[672]));
			radix2 #(.width(width)) rd_st2_545  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[545]), .rdlo_in(a2_wr[673]),  .coef_in(coef[132]), .rdup_out(a3_wr[545]), .rdlo_out(a3_wr[673]));
			radix2 #(.width(width)) rd_st2_546  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[546]), .rdlo_in(a2_wr[674]),  .coef_in(coef[136]), .rdup_out(a3_wr[546]), .rdlo_out(a3_wr[674]));
			radix2 #(.width(width)) rd_st2_547  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[547]), .rdlo_in(a2_wr[675]),  .coef_in(coef[140]), .rdup_out(a3_wr[547]), .rdlo_out(a3_wr[675]));
			radix2 #(.width(width)) rd_st2_548  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[548]), .rdlo_in(a2_wr[676]),  .coef_in(coef[144]), .rdup_out(a3_wr[548]), .rdlo_out(a3_wr[676]));
			radix2 #(.width(width)) rd_st2_549  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[549]), .rdlo_in(a2_wr[677]),  .coef_in(coef[148]), .rdup_out(a3_wr[549]), .rdlo_out(a3_wr[677]));
			radix2 #(.width(width)) rd_st2_550  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[550]), .rdlo_in(a2_wr[678]),  .coef_in(coef[152]), .rdup_out(a3_wr[550]), .rdlo_out(a3_wr[678]));
			radix2 #(.width(width)) rd_st2_551  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[551]), .rdlo_in(a2_wr[679]),  .coef_in(coef[156]), .rdup_out(a3_wr[551]), .rdlo_out(a3_wr[679]));
			radix2 #(.width(width)) rd_st2_552  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[552]), .rdlo_in(a2_wr[680]),  .coef_in(coef[160]), .rdup_out(a3_wr[552]), .rdlo_out(a3_wr[680]));
			radix2 #(.width(width)) rd_st2_553  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[553]), .rdlo_in(a2_wr[681]),  .coef_in(coef[164]), .rdup_out(a3_wr[553]), .rdlo_out(a3_wr[681]));
			radix2 #(.width(width)) rd_st2_554  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[554]), .rdlo_in(a2_wr[682]),  .coef_in(coef[168]), .rdup_out(a3_wr[554]), .rdlo_out(a3_wr[682]));
			radix2 #(.width(width)) rd_st2_555  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[555]), .rdlo_in(a2_wr[683]),  .coef_in(coef[172]), .rdup_out(a3_wr[555]), .rdlo_out(a3_wr[683]));
			radix2 #(.width(width)) rd_st2_556  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[556]), .rdlo_in(a2_wr[684]),  .coef_in(coef[176]), .rdup_out(a3_wr[556]), .rdlo_out(a3_wr[684]));
			radix2 #(.width(width)) rd_st2_557  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[557]), .rdlo_in(a2_wr[685]),  .coef_in(coef[180]), .rdup_out(a3_wr[557]), .rdlo_out(a3_wr[685]));
			radix2 #(.width(width)) rd_st2_558  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[558]), .rdlo_in(a2_wr[686]),  .coef_in(coef[184]), .rdup_out(a3_wr[558]), .rdlo_out(a3_wr[686]));
			radix2 #(.width(width)) rd_st2_559  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[559]), .rdlo_in(a2_wr[687]),  .coef_in(coef[188]), .rdup_out(a3_wr[559]), .rdlo_out(a3_wr[687]));
			radix2 #(.width(width)) rd_st2_560  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[560]), .rdlo_in(a2_wr[688]),  .coef_in(coef[192]), .rdup_out(a3_wr[560]), .rdlo_out(a3_wr[688]));
			radix2 #(.width(width)) rd_st2_561  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[561]), .rdlo_in(a2_wr[689]),  .coef_in(coef[196]), .rdup_out(a3_wr[561]), .rdlo_out(a3_wr[689]));
			radix2 #(.width(width)) rd_st2_562  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[562]), .rdlo_in(a2_wr[690]),  .coef_in(coef[200]), .rdup_out(a3_wr[562]), .rdlo_out(a3_wr[690]));
			radix2 #(.width(width)) rd_st2_563  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[563]), .rdlo_in(a2_wr[691]),  .coef_in(coef[204]), .rdup_out(a3_wr[563]), .rdlo_out(a3_wr[691]));
			radix2 #(.width(width)) rd_st2_564  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[564]), .rdlo_in(a2_wr[692]),  .coef_in(coef[208]), .rdup_out(a3_wr[564]), .rdlo_out(a3_wr[692]));
			radix2 #(.width(width)) rd_st2_565  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[565]), .rdlo_in(a2_wr[693]),  .coef_in(coef[212]), .rdup_out(a3_wr[565]), .rdlo_out(a3_wr[693]));
			radix2 #(.width(width)) rd_st2_566  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[566]), .rdlo_in(a2_wr[694]),  .coef_in(coef[216]), .rdup_out(a3_wr[566]), .rdlo_out(a3_wr[694]));
			radix2 #(.width(width)) rd_st2_567  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[567]), .rdlo_in(a2_wr[695]),  .coef_in(coef[220]), .rdup_out(a3_wr[567]), .rdlo_out(a3_wr[695]));
			radix2 #(.width(width)) rd_st2_568  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[568]), .rdlo_in(a2_wr[696]),  .coef_in(coef[224]), .rdup_out(a3_wr[568]), .rdlo_out(a3_wr[696]));
			radix2 #(.width(width)) rd_st2_569  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[569]), .rdlo_in(a2_wr[697]),  .coef_in(coef[228]), .rdup_out(a3_wr[569]), .rdlo_out(a3_wr[697]));
			radix2 #(.width(width)) rd_st2_570  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[570]), .rdlo_in(a2_wr[698]),  .coef_in(coef[232]), .rdup_out(a3_wr[570]), .rdlo_out(a3_wr[698]));
			radix2 #(.width(width)) rd_st2_571  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[571]), .rdlo_in(a2_wr[699]),  .coef_in(coef[236]), .rdup_out(a3_wr[571]), .rdlo_out(a3_wr[699]));
			radix2 #(.width(width)) rd_st2_572  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[572]), .rdlo_in(a2_wr[700]),  .coef_in(coef[240]), .rdup_out(a3_wr[572]), .rdlo_out(a3_wr[700]));
			radix2 #(.width(width)) rd_st2_573  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[573]), .rdlo_in(a2_wr[701]),  .coef_in(coef[244]), .rdup_out(a3_wr[573]), .rdlo_out(a3_wr[701]));
			radix2 #(.width(width)) rd_st2_574  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[574]), .rdlo_in(a2_wr[702]),  .coef_in(coef[248]), .rdup_out(a3_wr[574]), .rdlo_out(a3_wr[702]));
			radix2 #(.width(width)) rd_st2_575  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[575]), .rdlo_in(a2_wr[703]),  .coef_in(coef[252]), .rdup_out(a3_wr[575]), .rdlo_out(a3_wr[703]));
			radix2 #(.width(width)) rd_st2_576  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[576]), .rdlo_in(a2_wr[704]),  .coef_in(coef[256]), .rdup_out(a3_wr[576]), .rdlo_out(a3_wr[704]));
			radix2 #(.width(width)) rd_st2_577  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[577]), .rdlo_in(a2_wr[705]),  .coef_in(coef[260]), .rdup_out(a3_wr[577]), .rdlo_out(a3_wr[705]));
			radix2 #(.width(width)) rd_st2_578  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[578]), .rdlo_in(a2_wr[706]),  .coef_in(coef[264]), .rdup_out(a3_wr[578]), .rdlo_out(a3_wr[706]));
			radix2 #(.width(width)) rd_st2_579  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[579]), .rdlo_in(a2_wr[707]),  .coef_in(coef[268]), .rdup_out(a3_wr[579]), .rdlo_out(a3_wr[707]));
			radix2 #(.width(width)) rd_st2_580  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[580]), .rdlo_in(a2_wr[708]),  .coef_in(coef[272]), .rdup_out(a3_wr[580]), .rdlo_out(a3_wr[708]));
			radix2 #(.width(width)) rd_st2_581  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[581]), .rdlo_in(a2_wr[709]),  .coef_in(coef[276]), .rdup_out(a3_wr[581]), .rdlo_out(a3_wr[709]));
			radix2 #(.width(width)) rd_st2_582  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[582]), .rdlo_in(a2_wr[710]),  .coef_in(coef[280]), .rdup_out(a3_wr[582]), .rdlo_out(a3_wr[710]));
			radix2 #(.width(width)) rd_st2_583  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[583]), .rdlo_in(a2_wr[711]),  .coef_in(coef[284]), .rdup_out(a3_wr[583]), .rdlo_out(a3_wr[711]));
			radix2 #(.width(width)) rd_st2_584  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[584]), .rdlo_in(a2_wr[712]),  .coef_in(coef[288]), .rdup_out(a3_wr[584]), .rdlo_out(a3_wr[712]));
			radix2 #(.width(width)) rd_st2_585  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[585]), .rdlo_in(a2_wr[713]),  .coef_in(coef[292]), .rdup_out(a3_wr[585]), .rdlo_out(a3_wr[713]));
			radix2 #(.width(width)) rd_st2_586  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[586]), .rdlo_in(a2_wr[714]),  .coef_in(coef[296]), .rdup_out(a3_wr[586]), .rdlo_out(a3_wr[714]));
			radix2 #(.width(width)) rd_st2_587  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[587]), .rdlo_in(a2_wr[715]),  .coef_in(coef[300]), .rdup_out(a3_wr[587]), .rdlo_out(a3_wr[715]));
			radix2 #(.width(width)) rd_st2_588  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[588]), .rdlo_in(a2_wr[716]),  .coef_in(coef[304]), .rdup_out(a3_wr[588]), .rdlo_out(a3_wr[716]));
			radix2 #(.width(width)) rd_st2_589  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[589]), .rdlo_in(a2_wr[717]),  .coef_in(coef[308]), .rdup_out(a3_wr[589]), .rdlo_out(a3_wr[717]));
			radix2 #(.width(width)) rd_st2_590  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[590]), .rdlo_in(a2_wr[718]),  .coef_in(coef[312]), .rdup_out(a3_wr[590]), .rdlo_out(a3_wr[718]));
			radix2 #(.width(width)) rd_st2_591  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[591]), .rdlo_in(a2_wr[719]),  .coef_in(coef[316]), .rdup_out(a3_wr[591]), .rdlo_out(a3_wr[719]));
			radix2 #(.width(width)) rd_st2_592  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[592]), .rdlo_in(a2_wr[720]),  .coef_in(coef[320]), .rdup_out(a3_wr[592]), .rdlo_out(a3_wr[720]));
			radix2 #(.width(width)) rd_st2_593  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[593]), .rdlo_in(a2_wr[721]),  .coef_in(coef[324]), .rdup_out(a3_wr[593]), .rdlo_out(a3_wr[721]));
			radix2 #(.width(width)) rd_st2_594  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[594]), .rdlo_in(a2_wr[722]),  .coef_in(coef[328]), .rdup_out(a3_wr[594]), .rdlo_out(a3_wr[722]));
			radix2 #(.width(width)) rd_st2_595  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[595]), .rdlo_in(a2_wr[723]),  .coef_in(coef[332]), .rdup_out(a3_wr[595]), .rdlo_out(a3_wr[723]));
			radix2 #(.width(width)) rd_st2_596  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[596]), .rdlo_in(a2_wr[724]),  .coef_in(coef[336]), .rdup_out(a3_wr[596]), .rdlo_out(a3_wr[724]));
			radix2 #(.width(width)) rd_st2_597  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[597]), .rdlo_in(a2_wr[725]),  .coef_in(coef[340]), .rdup_out(a3_wr[597]), .rdlo_out(a3_wr[725]));
			radix2 #(.width(width)) rd_st2_598  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[598]), .rdlo_in(a2_wr[726]),  .coef_in(coef[344]), .rdup_out(a3_wr[598]), .rdlo_out(a3_wr[726]));
			radix2 #(.width(width)) rd_st2_599  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[599]), .rdlo_in(a2_wr[727]),  .coef_in(coef[348]), .rdup_out(a3_wr[599]), .rdlo_out(a3_wr[727]));
			radix2 #(.width(width)) rd_st2_600  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[600]), .rdlo_in(a2_wr[728]),  .coef_in(coef[352]), .rdup_out(a3_wr[600]), .rdlo_out(a3_wr[728]));
			radix2 #(.width(width)) rd_st2_601  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[601]), .rdlo_in(a2_wr[729]),  .coef_in(coef[356]), .rdup_out(a3_wr[601]), .rdlo_out(a3_wr[729]));
			radix2 #(.width(width)) rd_st2_602  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[602]), .rdlo_in(a2_wr[730]),  .coef_in(coef[360]), .rdup_out(a3_wr[602]), .rdlo_out(a3_wr[730]));
			radix2 #(.width(width)) rd_st2_603  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[603]), .rdlo_in(a2_wr[731]),  .coef_in(coef[364]), .rdup_out(a3_wr[603]), .rdlo_out(a3_wr[731]));
			radix2 #(.width(width)) rd_st2_604  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[604]), .rdlo_in(a2_wr[732]),  .coef_in(coef[368]), .rdup_out(a3_wr[604]), .rdlo_out(a3_wr[732]));
			radix2 #(.width(width)) rd_st2_605  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[605]), .rdlo_in(a2_wr[733]),  .coef_in(coef[372]), .rdup_out(a3_wr[605]), .rdlo_out(a3_wr[733]));
			radix2 #(.width(width)) rd_st2_606  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[606]), .rdlo_in(a2_wr[734]),  .coef_in(coef[376]), .rdup_out(a3_wr[606]), .rdlo_out(a3_wr[734]));
			radix2 #(.width(width)) rd_st2_607  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[607]), .rdlo_in(a2_wr[735]),  .coef_in(coef[380]), .rdup_out(a3_wr[607]), .rdlo_out(a3_wr[735]));
			radix2 #(.width(width)) rd_st2_608  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[608]), .rdlo_in(a2_wr[736]),  .coef_in(coef[384]), .rdup_out(a3_wr[608]), .rdlo_out(a3_wr[736]));
			radix2 #(.width(width)) rd_st2_609  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[609]), .rdlo_in(a2_wr[737]),  .coef_in(coef[388]), .rdup_out(a3_wr[609]), .rdlo_out(a3_wr[737]));
			radix2 #(.width(width)) rd_st2_610  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[610]), .rdlo_in(a2_wr[738]),  .coef_in(coef[392]), .rdup_out(a3_wr[610]), .rdlo_out(a3_wr[738]));
			radix2 #(.width(width)) rd_st2_611  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[611]), .rdlo_in(a2_wr[739]),  .coef_in(coef[396]), .rdup_out(a3_wr[611]), .rdlo_out(a3_wr[739]));
			radix2 #(.width(width)) rd_st2_612  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[612]), .rdlo_in(a2_wr[740]),  .coef_in(coef[400]), .rdup_out(a3_wr[612]), .rdlo_out(a3_wr[740]));
			radix2 #(.width(width)) rd_st2_613  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[613]), .rdlo_in(a2_wr[741]),  .coef_in(coef[404]), .rdup_out(a3_wr[613]), .rdlo_out(a3_wr[741]));
			radix2 #(.width(width)) rd_st2_614  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[614]), .rdlo_in(a2_wr[742]),  .coef_in(coef[408]), .rdup_out(a3_wr[614]), .rdlo_out(a3_wr[742]));
			radix2 #(.width(width)) rd_st2_615  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[615]), .rdlo_in(a2_wr[743]),  .coef_in(coef[412]), .rdup_out(a3_wr[615]), .rdlo_out(a3_wr[743]));
			radix2 #(.width(width)) rd_st2_616  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[616]), .rdlo_in(a2_wr[744]),  .coef_in(coef[416]), .rdup_out(a3_wr[616]), .rdlo_out(a3_wr[744]));
			radix2 #(.width(width)) rd_st2_617  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[617]), .rdlo_in(a2_wr[745]),  .coef_in(coef[420]), .rdup_out(a3_wr[617]), .rdlo_out(a3_wr[745]));
			radix2 #(.width(width)) rd_st2_618  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[618]), .rdlo_in(a2_wr[746]),  .coef_in(coef[424]), .rdup_out(a3_wr[618]), .rdlo_out(a3_wr[746]));
			radix2 #(.width(width)) rd_st2_619  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[619]), .rdlo_in(a2_wr[747]),  .coef_in(coef[428]), .rdup_out(a3_wr[619]), .rdlo_out(a3_wr[747]));
			radix2 #(.width(width)) rd_st2_620  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[620]), .rdlo_in(a2_wr[748]),  .coef_in(coef[432]), .rdup_out(a3_wr[620]), .rdlo_out(a3_wr[748]));
			radix2 #(.width(width)) rd_st2_621  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[621]), .rdlo_in(a2_wr[749]),  .coef_in(coef[436]), .rdup_out(a3_wr[621]), .rdlo_out(a3_wr[749]));
			radix2 #(.width(width)) rd_st2_622  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[622]), .rdlo_in(a2_wr[750]),  .coef_in(coef[440]), .rdup_out(a3_wr[622]), .rdlo_out(a3_wr[750]));
			radix2 #(.width(width)) rd_st2_623  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[623]), .rdlo_in(a2_wr[751]),  .coef_in(coef[444]), .rdup_out(a3_wr[623]), .rdlo_out(a3_wr[751]));
			radix2 #(.width(width)) rd_st2_624  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[624]), .rdlo_in(a2_wr[752]),  .coef_in(coef[448]), .rdup_out(a3_wr[624]), .rdlo_out(a3_wr[752]));
			radix2 #(.width(width)) rd_st2_625  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[625]), .rdlo_in(a2_wr[753]),  .coef_in(coef[452]), .rdup_out(a3_wr[625]), .rdlo_out(a3_wr[753]));
			radix2 #(.width(width)) rd_st2_626  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[626]), .rdlo_in(a2_wr[754]),  .coef_in(coef[456]), .rdup_out(a3_wr[626]), .rdlo_out(a3_wr[754]));
			radix2 #(.width(width)) rd_st2_627  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[627]), .rdlo_in(a2_wr[755]),  .coef_in(coef[460]), .rdup_out(a3_wr[627]), .rdlo_out(a3_wr[755]));
			radix2 #(.width(width)) rd_st2_628  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[628]), .rdlo_in(a2_wr[756]),  .coef_in(coef[464]), .rdup_out(a3_wr[628]), .rdlo_out(a3_wr[756]));
			radix2 #(.width(width)) rd_st2_629  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[629]), .rdlo_in(a2_wr[757]),  .coef_in(coef[468]), .rdup_out(a3_wr[629]), .rdlo_out(a3_wr[757]));
			radix2 #(.width(width)) rd_st2_630  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[630]), .rdlo_in(a2_wr[758]),  .coef_in(coef[472]), .rdup_out(a3_wr[630]), .rdlo_out(a3_wr[758]));
			radix2 #(.width(width)) rd_st2_631  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[631]), .rdlo_in(a2_wr[759]),  .coef_in(coef[476]), .rdup_out(a3_wr[631]), .rdlo_out(a3_wr[759]));
			radix2 #(.width(width)) rd_st2_632  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[632]), .rdlo_in(a2_wr[760]),  .coef_in(coef[480]), .rdup_out(a3_wr[632]), .rdlo_out(a3_wr[760]));
			radix2 #(.width(width)) rd_st2_633  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[633]), .rdlo_in(a2_wr[761]),  .coef_in(coef[484]), .rdup_out(a3_wr[633]), .rdlo_out(a3_wr[761]));
			radix2 #(.width(width)) rd_st2_634  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[634]), .rdlo_in(a2_wr[762]),  .coef_in(coef[488]), .rdup_out(a3_wr[634]), .rdlo_out(a3_wr[762]));
			radix2 #(.width(width)) rd_st2_635  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[635]), .rdlo_in(a2_wr[763]),  .coef_in(coef[492]), .rdup_out(a3_wr[635]), .rdlo_out(a3_wr[763]));
			radix2 #(.width(width)) rd_st2_636  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[636]), .rdlo_in(a2_wr[764]),  .coef_in(coef[496]), .rdup_out(a3_wr[636]), .rdlo_out(a3_wr[764]));
			radix2 #(.width(width)) rd_st2_637  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[637]), .rdlo_in(a2_wr[765]),  .coef_in(coef[500]), .rdup_out(a3_wr[637]), .rdlo_out(a3_wr[765]));
			radix2 #(.width(width)) rd_st2_638  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[638]), .rdlo_in(a2_wr[766]),  .coef_in(coef[504]), .rdup_out(a3_wr[638]), .rdlo_out(a3_wr[766]));
			radix2 #(.width(width)) rd_st2_639  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[639]), .rdlo_in(a2_wr[767]),  .coef_in(coef[508]), .rdup_out(a3_wr[639]), .rdlo_out(a3_wr[767]));
			radix2 #(.width(width)) rd_st2_768  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[768]), .rdlo_in(a2_wr[896]),  .coef_in(coef[0]), .rdup_out(a3_wr[768]), .rdlo_out(a3_wr[896]));
			radix2 #(.width(width)) rd_st2_769  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[769]), .rdlo_in(a2_wr[897]),  .coef_in(coef[4]), .rdup_out(a3_wr[769]), .rdlo_out(a3_wr[897]));
			radix2 #(.width(width)) rd_st2_770  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[770]), .rdlo_in(a2_wr[898]),  .coef_in(coef[8]), .rdup_out(a3_wr[770]), .rdlo_out(a3_wr[898]));
			radix2 #(.width(width)) rd_st2_771  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[771]), .rdlo_in(a2_wr[899]),  .coef_in(coef[12]), .rdup_out(a3_wr[771]), .rdlo_out(a3_wr[899]));
			radix2 #(.width(width)) rd_st2_772  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[772]), .rdlo_in(a2_wr[900]),  .coef_in(coef[16]), .rdup_out(a3_wr[772]), .rdlo_out(a3_wr[900]));
			radix2 #(.width(width)) rd_st2_773  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[773]), .rdlo_in(a2_wr[901]),  .coef_in(coef[20]), .rdup_out(a3_wr[773]), .rdlo_out(a3_wr[901]));
			radix2 #(.width(width)) rd_st2_774  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[774]), .rdlo_in(a2_wr[902]),  .coef_in(coef[24]), .rdup_out(a3_wr[774]), .rdlo_out(a3_wr[902]));
			radix2 #(.width(width)) rd_st2_775  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[775]), .rdlo_in(a2_wr[903]),  .coef_in(coef[28]), .rdup_out(a3_wr[775]), .rdlo_out(a3_wr[903]));
			radix2 #(.width(width)) rd_st2_776  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[776]), .rdlo_in(a2_wr[904]),  .coef_in(coef[32]), .rdup_out(a3_wr[776]), .rdlo_out(a3_wr[904]));
			radix2 #(.width(width)) rd_st2_777  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[777]), .rdlo_in(a2_wr[905]),  .coef_in(coef[36]), .rdup_out(a3_wr[777]), .rdlo_out(a3_wr[905]));
			radix2 #(.width(width)) rd_st2_778  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[778]), .rdlo_in(a2_wr[906]),  .coef_in(coef[40]), .rdup_out(a3_wr[778]), .rdlo_out(a3_wr[906]));
			radix2 #(.width(width)) rd_st2_779  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[779]), .rdlo_in(a2_wr[907]),  .coef_in(coef[44]), .rdup_out(a3_wr[779]), .rdlo_out(a3_wr[907]));
			radix2 #(.width(width)) rd_st2_780  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[780]), .rdlo_in(a2_wr[908]),  .coef_in(coef[48]), .rdup_out(a3_wr[780]), .rdlo_out(a3_wr[908]));
			radix2 #(.width(width)) rd_st2_781  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[781]), .rdlo_in(a2_wr[909]),  .coef_in(coef[52]), .rdup_out(a3_wr[781]), .rdlo_out(a3_wr[909]));
			radix2 #(.width(width)) rd_st2_782  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[782]), .rdlo_in(a2_wr[910]),  .coef_in(coef[56]), .rdup_out(a3_wr[782]), .rdlo_out(a3_wr[910]));
			radix2 #(.width(width)) rd_st2_783  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[783]), .rdlo_in(a2_wr[911]),  .coef_in(coef[60]), .rdup_out(a3_wr[783]), .rdlo_out(a3_wr[911]));
			radix2 #(.width(width)) rd_st2_784  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[784]), .rdlo_in(a2_wr[912]),  .coef_in(coef[64]), .rdup_out(a3_wr[784]), .rdlo_out(a3_wr[912]));
			radix2 #(.width(width)) rd_st2_785  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[785]), .rdlo_in(a2_wr[913]),  .coef_in(coef[68]), .rdup_out(a3_wr[785]), .rdlo_out(a3_wr[913]));
			radix2 #(.width(width)) rd_st2_786  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[786]), .rdlo_in(a2_wr[914]),  .coef_in(coef[72]), .rdup_out(a3_wr[786]), .rdlo_out(a3_wr[914]));
			radix2 #(.width(width)) rd_st2_787  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[787]), .rdlo_in(a2_wr[915]),  .coef_in(coef[76]), .rdup_out(a3_wr[787]), .rdlo_out(a3_wr[915]));
			radix2 #(.width(width)) rd_st2_788  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[788]), .rdlo_in(a2_wr[916]),  .coef_in(coef[80]), .rdup_out(a3_wr[788]), .rdlo_out(a3_wr[916]));
			radix2 #(.width(width)) rd_st2_789  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[789]), .rdlo_in(a2_wr[917]),  .coef_in(coef[84]), .rdup_out(a3_wr[789]), .rdlo_out(a3_wr[917]));
			radix2 #(.width(width)) rd_st2_790  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[790]), .rdlo_in(a2_wr[918]),  .coef_in(coef[88]), .rdup_out(a3_wr[790]), .rdlo_out(a3_wr[918]));
			radix2 #(.width(width)) rd_st2_791  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[791]), .rdlo_in(a2_wr[919]),  .coef_in(coef[92]), .rdup_out(a3_wr[791]), .rdlo_out(a3_wr[919]));
			radix2 #(.width(width)) rd_st2_792  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[792]), .rdlo_in(a2_wr[920]),  .coef_in(coef[96]), .rdup_out(a3_wr[792]), .rdlo_out(a3_wr[920]));
			radix2 #(.width(width)) rd_st2_793  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[793]), .rdlo_in(a2_wr[921]),  .coef_in(coef[100]), .rdup_out(a3_wr[793]), .rdlo_out(a3_wr[921]));
			radix2 #(.width(width)) rd_st2_794  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[794]), .rdlo_in(a2_wr[922]),  .coef_in(coef[104]), .rdup_out(a3_wr[794]), .rdlo_out(a3_wr[922]));
			radix2 #(.width(width)) rd_st2_795  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[795]), .rdlo_in(a2_wr[923]),  .coef_in(coef[108]), .rdup_out(a3_wr[795]), .rdlo_out(a3_wr[923]));
			radix2 #(.width(width)) rd_st2_796  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[796]), .rdlo_in(a2_wr[924]),  .coef_in(coef[112]), .rdup_out(a3_wr[796]), .rdlo_out(a3_wr[924]));
			radix2 #(.width(width)) rd_st2_797  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[797]), .rdlo_in(a2_wr[925]),  .coef_in(coef[116]), .rdup_out(a3_wr[797]), .rdlo_out(a3_wr[925]));
			radix2 #(.width(width)) rd_st2_798  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[798]), .rdlo_in(a2_wr[926]),  .coef_in(coef[120]), .rdup_out(a3_wr[798]), .rdlo_out(a3_wr[926]));
			radix2 #(.width(width)) rd_st2_799  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[799]), .rdlo_in(a2_wr[927]),  .coef_in(coef[124]), .rdup_out(a3_wr[799]), .rdlo_out(a3_wr[927]));
			radix2 #(.width(width)) rd_st2_800  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[800]), .rdlo_in(a2_wr[928]),  .coef_in(coef[128]), .rdup_out(a3_wr[800]), .rdlo_out(a3_wr[928]));
			radix2 #(.width(width)) rd_st2_801  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[801]), .rdlo_in(a2_wr[929]),  .coef_in(coef[132]), .rdup_out(a3_wr[801]), .rdlo_out(a3_wr[929]));
			radix2 #(.width(width)) rd_st2_802  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[802]), .rdlo_in(a2_wr[930]),  .coef_in(coef[136]), .rdup_out(a3_wr[802]), .rdlo_out(a3_wr[930]));
			radix2 #(.width(width)) rd_st2_803  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[803]), .rdlo_in(a2_wr[931]),  .coef_in(coef[140]), .rdup_out(a3_wr[803]), .rdlo_out(a3_wr[931]));
			radix2 #(.width(width)) rd_st2_804  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[804]), .rdlo_in(a2_wr[932]),  .coef_in(coef[144]), .rdup_out(a3_wr[804]), .rdlo_out(a3_wr[932]));
			radix2 #(.width(width)) rd_st2_805  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[805]), .rdlo_in(a2_wr[933]),  .coef_in(coef[148]), .rdup_out(a3_wr[805]), .rdlo_out(a3_wr[933]));
			radix2 #(.width(width)) rd_st2_806  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[806]), .rdlo_in(a2_wr[934]),  .coef_in(coef[152]), .rdup_out(a3_wr[806]), .rdlo_out(a3_wr[934]));
			radix2 #(.width(width)) rd_st2_807  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[807]), .rdlo_in(a2_wr[935]),  .coef_in(coef[156]), .rdup_out(a3_wr[807]), .rdlo_out(a3_wr[935]));
			radix2 #(.width(width)) rd_st2_808  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[808]), .rdlo_in(a2_wr[936]),  .coef_in(coef[160]), .rdup_out(a3_wr[808]), .rdlo_out(a3_wr[936]));
			radix2 #(.width(width)) rd_st2_809  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[809]), .rdlo_in(a2_wr[937]),  .coef_in(coef[164]), .rdup_out(a3_wr[809]), .rdlo_out(a3_wr[937]));
			radix2 #(.width(width)) rd_st2_810  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[810]), .rdlo_in(a2_wr[938]),  .coef_in(coef[168]), .rdup_out(a3_wr[810]), .rdlo_out(a3_wr[938]));
			radix2 #(.width(width)) rd_st2_811  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[811]), .rdlo_in(a2_wr[939]),  .coef_in(coef[172]), .rdup_out(a3_wr[811]), .rdlo_out(a3_wr[939]));
			radix2 #(.width(width)) rd_st2_812  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[812]), .rdlo_in(a2_wr[940]),  .coef_in(coef[176]), .rdup_out(a3_wr[812]), .rdlo_out(a3_wr[940]));
			radix2 #(.width(width)) rd_st2_813  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[813]), .rdlo_in(a2_wr[941]),  .coef_in(coef[180]), .rdup_out(a3_wr[813]), .rdlo_out(a3_wr[941]));
			radix2 #(.width(width)) rd_st2_814  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[814]), .rdlo_in(a2_wr[942]),  .coef_in(coef[184]), .rdup_out(a3_wr[814]), .rdlo_out(a3_wr[942]));
			radix2 #(.width(width)) rd_st2_815  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[815]), .rdlo_in(a2_wr[943]),  .coef_in(coef[188]), .rdup_out(a3_wr[815]), .rdlo_out(a3_wr[943]));
			radix2 #(.width(width)) rd_st2_816  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[816]), .rdlo_in(a2_wr[944]),  .coef_in(coef[192]), .rdup_out(a3_wr[816]), .rdlo_out(a3_wr[944]));
			radix2 #(.width(width)) rd_st2_817  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[817]), .rdlo_in(a2_wr[945]),  .coef_in(coef[196]), .rdup_out(a3_wr[817]), .rdlo_out(a3_wr[945]));
			radix2 #(.width(width)) rd_st2_818  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[818]), .rdlo_in(a2_wr[946]),  .coef_in(coef[200]), .rdup_out(a3_wr[818]), .rdlo_out(a3_wr[946]));
			radix2 #(.width(width)) rd_st2_819  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[819]), .rdlo_in(a2_wr[947]),  .coef_in(coef[204]), .rdup_out(a3_wr[819]), .rdlo_out(a3_wr[947]));
			radix2 #(.width(width)) rd_st2_820  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[820]), .rdlo_in(a2_wr[948]),  .coef_in(coef[208]), .rdup_out(a3_wr[820]), .rdlo_out(a3_wr[948]));
			radix2 #(.width(width)) rd_st2_821  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[821]), .rdlo_in(a2_wr[949]),  .coef_in(coef[212]), .rdup_out(a3_wr[821]), .rdlo_out(a3_wr[949]));
			radix2 #(.width(width)) rd_st2_822  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[822]), .rdlo_in(a2_wr[950]),  .coef_in(coef[216]), .rdup_out(a3_wr[822]), .rdlo_out(a3_wr[950]));
			radix2 #(.width(width)) rd_st2_823  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[823]), .rdlo_in(a2_wr[951]),  .coef_in(coef[220]), .rdup_out(a3_wr[823]), .rdlo_out(a3_wr[951]));
			radix2 #(.width(width)) rd_st2_824  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[824]), .rdlo_in(a2_wr[952]),  .coef_in(coef[224]), .rdup_out(a3_wr[824]), .rdlo_out(a3_wr[952]));
			radix2 #(.width(width)) rd_st2_825  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[825]), .rdlo_in(a2_wr[953]),  .coef_in(coef[228]), .rdup_out(a3_wr[825]), .rdlo_out(a3_wr[953]));
			radix2 #(.width(width)) rd_st2_826  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[826]), .rdlo_in(a2_wr[954]),  .coef_in(coef[232]), .rdup_out(a3_wr[826]), .rdlo_out(a3_wr[954]));
			radix2 #(.width(width)) rd_st2_827  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[827]), .rdlo_in(a2_wr[955]),  .coef_in(coef[236]), .rdup_out(a3_wr[827]), .rdlo_out(a3_wr[955]));
			radix2 #(.width(width)) rd_st2_828  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[828]), .rdlo_in(a2_wr[956]),  .coef_in(coef[240]), .rdup_out(a3_wr[828]), .rdlo_out(a3_wr[956]));
			radix2 #(.width(width)) rd_st2_829  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[829]), .rdlo_in(a2_wr[957]),  .coef_in(coef[244]), .rdup_out(a3_wr[829]), .rdlo_out(a3_wr[957]));
			radix2 #(.width(width)) rd_st2_830  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[830]), .rdlo_in(a2_wr[958]),  .coef_in(coef[248]), .rdup_out(a3_wr[830]), .rdlo_out(a3_wr[958]));
			radix2 #(.width(width)) rd_st2_831  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[831]), .rdlo_in(a2_wr[959]),  .coef_in(coef[252]), .rdup_out(a3_wr[831]), .rdlo_out(a3_wr[959]));
			radix2 #(.width(width)) rd_st2_832  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[832]), .rdlo_in(a2_wr[960]),  .coef_in(coef[256]), .rdup_out(a3_wr[832]), .rdlo_out(a3_wr[960]));
			radix2 #(.width(width)) rd_st2_833  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[833]), .rdlo_in(a2_wr[961]),  .coef_in(coef[260]), .rdup_out(a3_wr[833]), .rdlo_out(a3_wr[961]));
			radix2 #(.width(width)) rd_st2_834  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[834]), .rdlo_in(a2_wr[962]),  .coef_in(coef[264]), .rdup_out(a3_wr[834]), .rdlo_out(a3_wr[962]));
			radix2 #(.width(width)) rd_st2_835  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[835]), .rdlo_in(a2_wr[963]),  .coef_in(coef[268]), .rdup_out(a3_wr[835]), .rdlo_out(a3_wr[963]));
			radix2 #(.width(width)) rd_st2_836  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[836]), .rdlo_in(a2_wr[964]),  .coef_in(coef[272]), .rdup_out(a3_wr[836]), .rdlo_out(a3_wr[964]));
			radix2 #(.width(width)) rd_st2_837  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[837]), .rdlo_in(a2_wr[965]),  .coef_in(coef[276]), .rdup_out(a3_wr[837]), .rdlo_out(a3_wr[965]));
			radix2 #(.width(width)) rd_st2_838  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[838]), .rdlo_in(a2_wr[966]),  .coef_in(coef[280]), .rdup_out(a3_wr[838]), .rdlo_out(a3_wr[966]));
			radix2 #(.width(width)) rd_st2_839  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[839]), .rdlo_in(a2_wr[967]),  .coef_in(coef[284]), .rdup_out(a3_wr[839]), .rdlo_out(a3_wr[967]));
			radix2 #(.width(width)) rd_st2_840  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[840]), .rdlo_in(a2_wr[968]),  .coef_in(coef[288]), .rdup_out(a3_wr[840]), .rdlo_out(a3_wr[968]));
			radix2 #(.width(width)) rd_st2_841  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[841]), .rdlo_in(a2_wr[969]),  .coef_in(coef[292]), .rdup_out(a3_wr[841]), .rdlo_out(a3_wr[969]));
			radix2 #(.width(width)) rd_st2_842  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[842]), .rdlo_in(a2_wr[970]),  .coef_in(coef[296]), .rdup_out(a3_wr[842]), .rdlo_out(a3_wr[970]));
			radix2 #(.width(width)) rd_st2_843  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[843]), .rdlo_in(a2_wr[971]),  .coef_in(coef[300]), .rdup_out(a3_wr[843]), .rdlo_out(a3_wr[971]));
			radix2 #(.width(width)) rd_st2_844  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[844]), .rdlo_in(a2_wr[972]),  .coef_in(coef[304]), .rdup_out(a3_wr[844]), .rdlo_out(a3_wr[972]));
			radix2 #(.width(width)) rd_st2_845  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[845]), .rdlo_in(a2_wr[973]),  .coef_in(coef[308]), .rdup_out(a3_wr[845]), .rdlo_out(a3_wr[973]));
			radix2 #(.width(width)) rd_st2_846  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[846]), .rdlo_in(a2_wr[974]),  .coef_in(coef[312]), .rdup_out(a3_wr[846]), .rdlo_out(a3_wr[974]));
			radix2 #(.width(width)) rd_st2_847  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[847]), .rdlo_in(a2_wr[975]),  .coef_in(coef[316]), .rdup_out(a3_wr[847]), .rdlo_out(a3_wr[975]));
			radix2 #(.width(width)) rd_st2_848  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[848]), .rdlo_in(a2_wr[976]),  .coef_in(coef[320]), .rdup_out(a3_wr[848]), .rdlo_out(a3_wr[976]));
			radix2 #(.width(width)) rd_st2_849  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[849]), .rdlo_in(a2_wr[977]),  .coef_in(coef[324]), .rdup_out(a3_wr[849]), .rdlo_out(a3_wr[977]));
			radix2 #(.width(width)) rd_st2_850  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[850]), .rdlo_in(a2_wr[978]),  .coef_in(coef[328]), .rdup_out(a3_wr[850]), .rdlo_out(a3_wr[978]));
			radix2 #(.width(width)) rd_st2_851  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[851]), .rdlo_in(a2_wr[979]),  .coef_in(coef[332]), .rdup_out(a3_wr[851]), .rdlo_out(a3_wr[979]));
			radix2 #(.width(width)) rd_st2_852  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[852]), .rdlo_in(a2_wr[980]),  .coef_in(coef[336]), .rdup_out(a3_wr[852]), .rdlo_out(a3_wr[980]));
			radix2 #(.width(width)) rd_st2_853  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[853]), .rdlo_in(a2_wr[981]),  .coef_in(coef[340]), .rdup_out(a3_wr[853]), .rdlo_out(a3_wr[981]));
			radix2 #(.width(width)) rd_st2_854  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[854]), .rdlo_in(a2_wr[982]),  .coef_in(coef[344]), .rdup_out(a3_wr[854]), .rdlo_out(a3_wr[982]));
			radix2 #(.width(width)) rd_st2_855  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[855]), .rdlo_in(a2_wr[983]),  .coef_in(coef[348]), .rdup_out(a3_wr[855]), .rdlo_out(a3_wr[983]));
			radix2 #(.width(width)) rd_st2_856  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[856]), .rdlo_in(a2_wr[984]),  .coef_in(coef[352]), .rdup_out(a3_wr[856]), .rdlo_out(a3_wr[984]));
			radix2 #(.width(width)) rd_st2_857  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[857]), .rdlo_in(a2_wr[985]),  .coef_in(coef[356]), .rdup_out(a3_wr[857]), .rdlo_out(a3_wr[985]));
			radix2 #(.width(width)) rd_st2_858  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[858]), .rdlo_in(a2_wr[986]),  .coef_in(coef[360]), .rdup_out(a3_wr[858]), .rdlo_out(a3_wr[986]));
			radix2 #(.width(width)) rd_st2_859  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[859]), .rdlo_in(a2_wr[987]),  .coef_in(coef[364]), .rdup_out(a3_wr[859]), .rdlo_out(a3_wr[987]));
			radix2 #(.width(width)) rd_st2_860  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[860]), .rdlo_in(a2_wr[988]),  .coef_in(coef[368]), .rdup_out(a3_wr[860]), .rdlo_out(a3_wr[988]));
			radix2 #(.width(width)) rd_st2_861  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[861]), .rdlo_in(a2_wr[989]),  .coef_in(coef[372]), .rdup_out(a3_wr[861]), .rdlo_out(a3_wr[989]));
			radix2 #(.width(width)) rd_st2_862  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[862]), .rdlo_in(a2_wr[990]),  .coef_in(coef[376]), .rdup_out(a3_wr[862]), .rdlo_out(a3_wr[990]));
			radix2 #(.width(width)) rd_st2_863  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[863]), .rdlo_in(a2_wr[991]),  .coef_in(coef[380]), .rdup_out(a3_wr[863]), .rdlo_out(a3_wr[991]));
			radix2 #(.width(width)) rd_st2_864  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[864]), .rdlo_in(a2_wr[992]),  .coef_in(coef[384]), .rdup_out(a3_wr[864]), .rdlo_out(a3_wr[992]));
			radix2 #(.width(width)) rd_st2_865  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[865]), .rdlo_in(a2_wr[993]),  .coef_in(coef[388]), .rdup_out(a3_wr[865]), .rdlo_out(a3_wr[993]));
			radix2 #(.width(width)) rd_st2_866  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[866]), .rdlo_in(a2_wr[994]),  .coef_in(coef[392]), .rdup_out(a3_wr[866]), .rdlo_out(a3_wr[994]));
			radix2 #(.width(width)) rd_st2_867  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[867]), .rdlo_in(a2_wr[995]),  .coef_in(coef[396]), .rdup_out(a3_wr[867]), .rdlo_out(a3_wr[995]));
			radix2 #(.width(width)) rd_st2_868  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[868]), .rdlo_in(a2_wr[996]),  .coef_in(coef[400]), .rdup_out(a3_wr[868]), .rdlo_out(a3_wr[996]));
			radix2 #(.width(width)) rd_st2_869  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[869]), .rdlo_in(a2_wr[997]),  .coef_in(coef[404]), .rdup_out(a3_wr[869]), .rdlo_out(a3_wr[997]));
			radix2 #(.width(width)) rd_st2_870  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[870]), .rdlo_in(a2_wr[998]),  .coef_in(coef[408]), .rdup_out(a3_wr[870]), .rdlo_out(a3_wr[998]));
			radix2 #(.width(width)) rd_st2_871  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[871]), .rdlo_in(a2_wr[999]),  .coef_in(coef[412]), .rdup_out(a3_wr[871]), .rdlo_out(a3_wr[999]));
			radix2 #(.width(width)) rd_st2_872  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[872]), .rdlo_in(a2_wr[1000]),  .coef_in(coef[416]), .rdup_out(a3_wr[872]), .rdlo_out(a3_wr[1000]));
			radix2 #(.width(width)) rd_st2_873  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[873]), .rdlo_in(a2_wr[1001]),  .coef_in(coef[420]), .rdup_out(a3_wr[873]), .rdlo_out(a3_wr[1001]));
			radix2 #(.width(width)) rd_st2_874  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[874]), .rdlo_in(a2_wr[1002]),  .coef_in(coef[424]), .rdup_out(a3_wr[874]), .rdlo_out(a3_wr[1002]));
			radix2 #(.width(width)) rd_st2_875  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[875]), .rdlo_in(a2_wr[1003]),  .coef_in(coef[428]), .rdup_out(a3_wr[875]), .rdlo_out(a3_wr[1003]));
			radix2 #(.width(width)) rd_st2_876  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[876]), .rdlo_in(a2_wr[1004]),  .coef_in(coef[432]), .rdup_out(a3_wr[876]), .rdlo_out(a3_wr[1004]));
			radix2 #(.width(width)) rd_st2_877  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[877]), .rdlo_in(a2_wr[1005]),  .coef_in(coef[436]), .rdup_out(a3_wr[877]), .rdlo_out(a3_wr[1005]));
			radix2 #(.width(width)) rd_st2_878  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[878]), .rdlo_in(a2_wr[1006]),  .coef_in(coef[440]), .rdup_out(a3_wr[878]), .rdlo_out(a3_wr[1006]));
			radix2 #(.width(width)) rd_st2_879  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[879]), .rdlo_in(a2_wr[1007]),  .coef_in(coef[444]), .rdup_out(a3_wr[879]), .rdlo_out(a3_wr[1007]));
			radix2 #(.width(width)) rd_st2_880  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[880]), .rdlo_in(a2_wr[1008]),  .coef_in(coef[448]), .rdup_out(a3_wr[880]), .rdlo_out(a3_wr[1008]));
			radix2 #(.width(width)) rd_st2_881  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[881]), .rdlo_in(a2_wr[1009]),  .coef_in(coef[452]), .rdup_out(a3_wr[881]), .rdlo_out(a3_wr[1009]));
			radix2 #(.width(width)) rd_st2_882  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[882]), .rdlo_in(a2_wr[1010]),  .coef_in(coef[456]), .rdup_out(a3_wr[882]), .rdlo_out(a3_wr[1010]));
			radix2 #(.width(width)) rd_st2_883  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[883]), .rdlo_in(a2_wr[1011]),  .coef_in(coef[460]), .rdup_out(a3_wr[883]), .rdlo_out(a3_wr[1011]));
			radix2 #(.width(width)) rd_st2_884  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[884]), .rdlo_in(a2_wr[1012]),  .coef_in(coef[464]), .rdup_out(a3_wr[884]), .rdlo_out(a3_wr[1012]));
			radix2 #(.width(width)) rd_st2_885  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[885]), .rdlo_in(a2_wr[1013]),  .coef_in(coef[468]), .rdup_out(a3_wr[885]), .rdlo_out(a3_wr[1013]));
			radix2 #(.width(width)) rd_st2_886  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[886]), .rdlo_in(a2_wr[1014]),  .coef_in(coef[472]), .rdup_out(a3_wr[886]), .rdlo_out(a3_wr[1014]));
			radix2 #(.width(width)) rd_st2_887  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[887]), .rdlo_in(a2_wr[1015]),  .coef_in(coef[476]), .rdup_out(a3_wr[887]), .rdlo_out(a3_wr[1015]));
			radix2 #(.width(width)) rd_st2_888  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[888]), .rdlo_in(a2_wr[1016]),  .coef_in(coef[480]), .rdup_out(a3_wr[888]), .rdlo_out(a3_wr[1016]));
			radix2 #(.width(width)) rd_st2_889  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[889]), .rdlo_in(a2_wr[1017]),  .coef_in(coef[484]), .rdup_out(a3_wr[889]), .rdlo_out(a3_wr[1017]));
			radix2 #(.width(width)) rd_st2_890  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[890]), .rdlo_in(a2_wr[1018]),  .coef_in(coef[488]), .rdup_out(a3_wr[890]), .rdlo_out(a3_wr[1018]));
			radix2 #(.width(width)) rd_st2_891  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[891]), .rdlo_in(a2_wr[1019]),  .coef_in(coef[492]), .rdup_out(a3_wr[891]), .rdlo_out(a3_wr[1019]));
			radix2 #(.width(width)) rd_st2_892  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[892]), .rdlo_in(a2_wr[1020]),  .coef_in(coef[496]), .rdup_out(a3_wr[892]), .rdlo_out(a3_wr[1020]));
			radix2 #(.width(width)) rd_st2_893  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[893]), .rdlo_in(a2_wr[1021]),  .coef_in(coef[500]), .rdup_out(a3_wr[893]), .rdlo_out(a3_wr[1021]));
			radix2 #(.width(width)) rd_st2_894  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[894]), .rdlo_in(a2_wr[1022]),  .coef_in(coef[504]), .rdup_out(a3_wr[894]), .rdlo_out(a3_wr[1022]));
			radix2 #(.width(width)) rd_st2_895  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[895]), .rdlo_in(a2_wr[1023]),  .coef_in(coef[508]), .rdup_out(a3_wr[895]), .rdlo_out(a3_wr[1023]));

		//--- radix stage 3
			radix2 #(.width(width)) rd_st3_0   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[0]), .rdlo_in(a3_wr[64]),  .coef_in(coef[0]), .rdup_out(a4_wr[0]), .rdlo_out(a4_wr[64]));
			radix2 #(.width(width)) rd_st3_1   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1]), .rdlo_in(a3_wr[65]),  .coef_in(coef[8]), .rdup_out(a4_wr[1]), .rdlo_out(a4_wr[65]));
			radix2 #(.width(width)) rd_st3_2   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[2]), .rdlo_in(a3_wr[66]),  .coef_in(coef[16]), .rdup_out(a4_wr[2]), .rdlo_out(a4_wr[66]));
			radix2 #(.width(width)) rd_st3_3   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[3]), .rdlo_in(a3_wr[67]),  .coef_in(coef[24]), .rdup_out(a4_wr[3]), .rdlo_out(a4_wr[67]));
			radix2 #(.width(width)) rd_st3_4   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[4]), .rdlo_in(a3_wr[68]),  .coef_in(coef[32]), .rdup_out(a4_wr[4]), .rdlo_out(a4_wr[68]));
			radix2 #(.width(width)) rd_st3_5   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[5]), .rdlo_in(a3_wr[69]),  .coef_in(coef[40]), .rdup_out(a4_wr[5]), .rdlo_out(a4_wr[69]));
			radix2 #(.width(width)) rd_st3_6   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[6]), .rdlo_in(a3_wr[70]),  .coef_in(coef[48]), .rdup_out(a4_wr[6]), .rdlo_out(a4_wr[70]));
			radix2 #(.width(width)) rd_st3_7   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[7]), .rdlo_in(a3_wr[71]),  .coef_in(coef[56]), .rdup_out(a4_wr[7]), .rdlo_out(a4_wr[71]));
			radix2 #(.width(width)) rd_st3_8   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[8]), .rdlo_in(a3_wr[72]),  .coef_in(coef[64]), .rdup_out(a4_wr[8]), .rdlo_out(a4_wr[72]));
			radix2 #(.width(width)) rd_st3_9   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[9]), .rdlo_in(a3_wr[73]),  .coef_in(coef[72]), .rdup_out(a4_wr[9]), .rdlo_out(a4_wr[73]));
			radix2 #(.width(width)) rd_st3_10  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[10]), .rdlo_in(a3_wr[74]),  .coef_in(coef[80]), .rdup_out(a4_wr[10]), .rdlo_out(a4_wr[74]));
			radix2 #(.width(width)) rd_st3_11  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[11]), .rdlo_in(a3_wr[75]),  .coef_in(coef[88]), .rdup_out(a4_wr[11]), .rdlo_out(a4_wr[75]));
			radix2 #(.width(width)) rd_st3_12  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[12]), .rdlo_in(a3_wr[76]),  .coef_in(coef[96]), .rdup_out(a4_wr[12]), .rdlo_out(a4_wr[76]));
			radix2 #(.width(width)) rd_st3_13  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[13]), .rdlo_in(a3_wr[77]),  .coef_in(coef[104]), .rdup_out(a4_wr[13]), .rdlo_out(a4_wr[77]));
			radix2 #(.width(width)) rd_st3_14  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[14]), .rdlo_in(a3_wr[78]),  .coef_in(coef[112]), .rdup_out(a4_wr[14]), .rdlo_out(a4_wr[78]));
			radix2 #(.width(width)) rd_st3_15  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[15]), .rdlo_in(a3_wr[79]),  .coef_in(coef[120]), .rdup_out(a4_wr[15]), .rdlo_out(a4_wr[79]));
			radix2 #(.width(width)) rd_st3_16  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[16]), .rdlo_in(a3_wr[80]),  .coef_in(coef[128]), .rdup_out(a4_wr[16]), .rdlo_out(a4_wr[80]));
			radix2 #(.width(width)) rd_st3_17  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[17]), .rdlo_in(a3_wr[81]),  .coef_in(coef[136]), .rdup_out(a4_wr[17]), .rdlo_out(a4_wr[81]));
			radix2 #(.width(width)) rd_st3_18  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[18]), .rdlo_in(a3_wr[82]),  .coef_in(coef[144]), .rdup_out(a4_wr[18]), .rdlo_out(a4_wr[82]));
			radix2 #(.width(width)) rd_st3_19  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[19]), .rdlo_in(a3_wr[83]),  .coef_in(coef[152]), .rdup_out(a4_wr[19]), .rdlo_out(a4_wr[83]));
			radix2 #(.width(width)) rd_st3_20  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[20]), .rdlo_in(a3_wr[84]),  .coef_in(coef[160]), .rdup_out(a4_wr[20]), .rdlo_out(a4_wr[84]));
			radix2 #(.width(width)) rd_st3_21  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[21]), .rdlo_in(a3_wr[85]),  .coef_in(coef[168]), .rdup_out(a4_wr[21]), .rdlo_out(a4_wr[85]));
			radix2 #(.width(width)) rd_st3_22  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[22]), .rdlo_in(a3_wr[86]),  .coef_in(coef[176]), .rdup_out(a4_wr[22]), .rdlo_out(a4_wr[86]));
			radix2 #(.width(width)) rd_st3_23  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[23]), .rdlo_in(a3_wr[87]),  .coef_in(coef[184]), .rdup_out(a4_wr[23]), .rdlo_out(a4_wr[87]));
			radix2 #(.width(width)) rd_st3_24  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[24]), .rdlo_in(a3_wr[88]),  .coef_in(coef[192]), .rdup_out(a4_wr[24]), .rdlo_out(a4_wr[88]));
			radix2 #(.width(width)) rd_st3_25  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[25]), .rdlo_in(a3_wr[89]),  .coef_in(coef[200]), .rdup_out(a4_wr[25]), .rdlo_out(a4_wr[89]));
			radix2 #(.width(width)) rd_st3_26  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[26]), .rdlo_in(a3_wr[90]),  .coef_in(coef[208]), .rdup_out(a4_wr[26]), .rdlo_out(a4_wr[90]));
			radix2 #(.width(width)) rd_st3_27  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[27]), .rdlo_in(a3_wr[91]),  .coef_in(coef[216]), .rdup_out(a4_wr[27]), .rdlo_out(a4_wr[91]));
			radix2 #(.width(width)) rd_st3_28  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[28]), .rdlo_in(a3_wr[92]),  .coef_in(coef[224]), .rdup_out(a4_wr[28]), .rdlo_out(a4_wr[92]));
			radix2 #(.width(width)) rd_st3_29  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[29]), .rdlo_in(a3_wr[93]),  .coef_in(coef[232]), .rdup_out(a4_wr[29]), .rdlo_out(a4_wr[93]));
			radix2 #(.width(width)) rd_st3_30  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[30]), .rdlo_in(a3_wr[94]),  .coef_in(coef[240]), .rdup_out(a4_wr[30]), .rdlo_out(a4_wr[94]));
			radix2 #(.width(width)) rd_st3_31  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[31]), .rdlo_in(a3_wr[95]),  .coef_in(coef[248]), .rdup_out(a4_wr[31]), .rdlo_out(a4_wr[95]));
			radix2 #(.width(width)) rd_st3_32  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[32]), .rdlo_in(a3_wr[96]),  .coef_in(coef[256]), .rdup_out(a4_wr[32]), .rdlo_out(a4_wr[96]));
			radix2 #(.width(width)) rd_st3_33  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[33]), .rdlo_in(a3_wr[97]),  .coef_in(coef[264]), .rdup_out(a4_wr[33]), .rdlo_out(a4_wr[97]));
			radix2 #(.width(width)) rd_st3_34  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[34]), .rdlo_in(a3_wr[98]),  .coef_in(coef[272]), .rdup_out(a4_wr[34]), .rdlo_out(a4_wr[98]));
			radix2 #(.width(width)) rd_st3_35  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[35]), .rdlo_in(a3_wr[99]),  .coef_in(coef[280]), .rdup_out(a4_wr[35]), .rdlo_out(a4_wr[99]));
			radix2 #(.width(width)) rd_st3_36  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[36]), .rdlo_in(a3_wr[100]),  .coef_in(coef[288]), .rdup_out(a4_wr[36]), .rdlo_out(a4_wr[100]));
			radix2 #(.width(width)) rd_st3_37  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[37]), .rdlo_in(a3_wr[101]),  .coef_in(coef[296]), .rdup_out(a4_wr[37]), .rdlo_out(a4_wr[101]));
			radix2 #(.width(width)) rd_st3_38  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[38]), .rdlo_in(a3_wr[102]),  .coef_in(coef[304]), .rdup_out(a4_wr[38]), .rdlo_out(a4_wr[102]));
			radix2 #(.width(width)) rd_st3_39  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[39]), .rdlo_in(a3_wr[103]),  .coef_in(coef[312]), .rdup_out(a4_wr[39]), .rdlo_out(a4_wr[103]));
			radix2 #(.width(width)) rd_st3_40  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[40]), .rdlo_in(a3_wr[104]),  .coef_in(coef[320]), .rdup_out(a4_wr[40]), .rdlo_out(a4_wr[104]));
			radix2 #(.width(width)) rd_st3_41  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[41]), .rdlo_in(a3_wr[105]),  .coef_in(coef[328]), .rdup_out(a4_wr[41]), .rdlo_out(a4_wr[105]));
			radix2 #(.width(width)) rd_st3_42  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[42]), .rdlo_in(a3_wr[106]),  .coef_in(coef[336]), .rdup_out(a4_wr[42]), .rdlo_out(a4_wr[106]));
			radix2 #(.width(width)) rd_st3_43  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[43]), .rdlo_in(a3_wr[107]),  .coef_in(coef[344]), .rdup_out(a4_wr[43]), .rdlo_out(a4_wr[107]));
			radix2 #(.width(width)) rd_st3_44  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[44]), .rdlo_in(a3_wr[108]),  .coef_in(coef[352]), .rdup_out(a4_wr[44]), .rdlo_out(a4_wr[108]));
			radix2 #(.width(width)) rd_st3_45  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[45]), .rdlo_in(a3_wr[109]),  .coef_in(coef[360]), .rdup_out(a4_wr[45]), .rdlo_out(a4_wr[109]));
			radix2 #(.width(width)) rd_st3_46  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[46]), .rdlo_in(a3_wr[110]),  .coef_in(coef[368]), .rdup_out(a4_wr[46]), .rdlo_out(a4_wr[110]));
			radix2 #(.width(width)) rd_st3_47  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[47]), .rdlo_in(a3_wr[111]),  .coef_in(coef[376]), .rdup_out(a4_wr[47]), .rdlo_out(a4_wr[111]));
			radix2 #(.width(width)) rd_st3_48  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[48]), .rdlo_in(a3_wr[112]),  .coef_in(coef[384]), .rdup_out(a4_wr[48]), .rdlo_out(a4_wr[112]));
			radix2 #(.width(width)) rd_st3_49  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[49]), .rdlo_in(a3_wr[113]),  .coef_in(coef[392]), .rdup_out(a4_wr[49]), .rdlo_out(a4_wr[113]));
			radix2 #(.width(width)) rd_st3_50  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[50]), .rdlo_in(a3_wr[114]),  .coef_in(coef[400]), .rdup_out(a4_wr[50]), .rdlo_out(a4_wr[114]));
			radix2 #(.width(width)) rd_st3_51  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[51]), .rdlo_in(a3_wr[115]),  .coef_in(coef[408]), .rdup_out(a4_wr[51]), .rdlo_out(a4_wr[115]));
			radix2 #(.width(width)) rd_st3_52  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[52]), .rdlo_in(a3_wr[116]),  .coef_in(coef[416]), .rdup_out(a4_wr[52]), .rdlo_out(a4_wr[116]));
			radix2 #(.width(width)) rd_st3_53  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[53]), .rdlo_in(a3_wr[117]),  .coef_in(coef[424]), .rdup_out(a4_wr[53]), .rdlo_out(a4_wr[117]));
			radix2 #(.width(width)) rd_st3_54  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[54]), .rdlo_in(a3_wr[118]),  .coef_in(coef[432]), .rdup_out(a4_wr[54]), .rdlo_out(a4_wr[118]));
			radix2 #(.width(width)) rd_st3_55  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[55]), .rdlo_in(a3_wr[119]),  .coef_in(coef[440]), .rdup_out(a4_wr[55]), .rdlo_out(a4_wr[119]));
			radix2 #(.width(width)) rd_st3_56  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[56]), .rdlo_in(a3_wr[120]),  .coef_in(coef[448]), .rdup_out(a4_wr[56]), .rdlo_out(a4_wr[120]));
			radix2 #(.width(width)) rd_st3_57  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[57]), .rdlo_in(a3_wr[121]),  .coef_in(coef[456]), .rdup_out(a4_wr[57]), .rdlo_out(a4_wr[121]));
			radix2 #(.width(width)) rd_st3_58  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[58]), .rdlo_in(a3_wr[122]),  .coef_in(coef[464]), .rdup_out(a4_wr[58]), .rdlo_out(a4_wr[122]));
			radix2 #(.width(width)) rd_st3_59  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[59]), .rdlo_in(a3_wr[123]),  .coef_in(coef[472]), .rdup_out(a4_wr[59]), .rdlo_out(a4_wr[123]));
			radix2 #(.width(width)) rd_st3_60  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[60]), .rdlo_in(a3_wr[124]),  .coef_in(coef[480]), .rdup_out(a4_wr[60]), .rdlo_out(a4_wr[124]));
			radix2 #(.width(width)) rd_st3_61  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[61]), .rdlo_in(a3_wr[125]),  .coef_in(coef[488]), .rdup_out(a4_wr[61]), .rdlo_out(a4_wr[125]));
			radix2 #(.width(width)) rd_st3_62  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[62]), .rdlo_in(a3_wr[126]),  .coef_in(coef[496]), .rdup_out(a4_wr[62]), .rdlo_out(a4_wr[126]));
			radix2 #(.width(width)) rd_st3_63  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[63]), .rdlo_in(a3_wr[127]),  .coef_in(coef[504]), .rdup_out(a4_wr[63]), .rdlo_out(a4_wr[127]));
			radix2 #(.width(width)) rd_st3_128  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[128]), .rdlo_in(a3_wr[192]),  .coef_in(coef[0]), .rdup_out(a4_wr[128]), .rdlo_out(a4_wr[192]));
			radix2 #(.width(width)) rd_st3_129  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[129]), .rdlo_in(a3_wr[193]),  .coef_in(coef[8]), .rdup_out(a4_wr[129]), .rdlo_out(a4_wr[193]));
			radix2 #(.width(width)) rd_st3_130  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[130]), .rdlo_in(a3_wr[194]),  .coef_in(coef[16]), .rdup_out(a4_wr[130]), .rdlo_out(a4_wr[194]));
			radix2 #(.width(width)) rd_st3_131  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[131]), .rdlo_in(a3_wr[195]),  .coef_in(coef[24]), .rdup_out(a4_wr[131]), .rdlo_out(a4_wr[195]));
			radix2 #(.width(width)) rd_st3_132  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[132]), .rdlo_in(a3_wr[196]),  .coef_in(coef[32]), .rdup_out(a4_wr[132]), .rdlo_out(a4_wr[196]));
			radix2 #(.width(width)) rd_st3_133  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[133]), .rdlo_in(a3_wr[197]),  .coef_in(coef[40]), .rdup_out(a4_wr[133]), .rdlo_out(a4_wr[197]));
			radix2 #(.width(width)) rd_st3_134  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[134]), .rdlo_in(a3_wr[198]),  .coef_in(coef[48]), .rdup_out(a4_wr[134]), .rdlo_out(a4_wr[198]));
			radix2 #(.width(width)) rd_st3_135  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[135]), .rdlo_in(a3_wr[199]),  .coef_in(coef[56]), .rdup_out(a4_wr[135]), .rdlo_out(a4_wr[199]));
			radix2 #(.width(width)) rd_st3_136  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[136]), .rdlo_in(a3_wr[200]),  .coef_in(coef[64]), .rdup_out(a4_wr[136]), .rdlo_out(a4_wr[200]));
			radix2 #(.width(width)) rd_st3_137  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[137]), .rdlo_in(a3_wr[201]),  .coef_in(coef[72]), .rdup_out(a4_wr[137]), .rdlo_out(a4_wr[201]));
			radix2 #(.width(width)) rd_st3_138  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[138]), .rdlo_in(a3_wr[202]),  .coef_in(coef[80]), .rdup_out(a4_wr[138]), .rdlo_out(a4_wr[202]));
			radix2 #(.width(width)) rd_st3_139  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[139]), .rdlo_in(a3_wr[203]),  .coef_in(coef[88]), .rdup_out(a4_wr[139]), .rdlo_out(a4_wr[203]));
			radix2 #(.width(width)) rd_st3_140  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[140]), .rdlo_in(a3_wr[204]),  .coef_in(coef[96]), .rdup_out(a4_wr[140]), .rdlo_out(a4_wr[204]));
			radix2 #(.width(width)) rd_st3_141  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[141]), .rdlo_in(a3_wr[205]),  .coef_in(coef[104]), .rdup_out(a4_wr[141]), .rdlo_out(a4_wr[205]));
			radix2 #(.width(width)) rd_st3_142  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[142]), .rdlo_in(a3_wr[206]),  .coef_in(coef[112]), .rdup_out(a4_wr[142]), .rdlo_out(a4_wr[206]));
			radix2 #(.width(width)) rd_st3_143  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[143]), .rdlo_in(a3_wr[207]),  .coef_in(coef[120]), .rdup_out(a4_wr[143]), .rdlo_out(a4_wr[207]));
			radix2 #(.width(width)) rd_st3_144  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[144]), .rdlo_in(a3_wr[208]),  .coef_in(coef[128]), .rdup_out(a4_wr[144]), .rdlo_out(a4_wr[208]));
			radix2 #(.width(width)) rd_st3_145  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[145]), .rdlo_in(a3_wr[209]),  .coef_in(coef[136]), .rdup_out(a4_wr[145]), .rdlo_out(a4_wr[209]));
			radix2 #(.width(width)) rd_st3_146  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[146]), .rdlo_in(a3_wr[210]),  .coef_in(coef[144]), .rdup_out(a4_wr[146]), .rdlo_out(a4_wr[210]));
			radix2 #(.width(width)) rd_st3_147  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[147]), .rdlo_in(a3_wr[211]),  .coef_in(coef[152]), .rdup_out(a4_wr[147]), .rdlo_out(a4_wr[211]));
			radix2 #(.width(width)) rd_st3_148  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[148]), .rdlo_in(a3_wr[212]),  .coef_in(coef[160]), .rdup_out(a4_wr[148]), .rdlo_out(a4_wr[212]));
			radix2 #(.width(width)) rd_st3_149  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[149]), .rdlo_in(a3_wr[213]),  .coef_in(coef[168]), .rdup_out(a4_wr[149]), .rdlo_out(a4_wr[213]));
			radix2 #(.width(width)) rd_st3_150  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[150]), .rdlo_in(a3_wr[214]),  .coef_in(coef[176]), .rdup_out(a4_wr[150]), .rdlo_out(a4_wr[214]));
			radix2 #(.width(width)) rd_st3_151  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[151]), .rdlo_in(a3_wr[215]),  .coef_in(coef[184]), .rdup_out(a4_wr[151]), .rdlo_out(a4_wr[215]));
			radix2 #(.width(width)) rd_st3_152  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[152]), .rdlo_in(a3_wr[216]),  .coef_in(coef[192]), .rdup_out(a4_wr[152]), .rdlo_out(a4_wr[216]));
			radix2 #(.width(width)) rd_st3_153  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[153]), .rdlo_in(a3_wr[217]),  .coef_in(coef[200]), .rdup_out(a4_wr[153]), .rdlo_out(a4_wr[217]));
			radix2 #(.width(width)) rd_st3_154  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[154]), .rdlo_in(a3_wr[218]),  .coef_in(coef[208]), .rdup_out(a4_wr[154]), .rdlo_out(a4_wr[218]));
			radix2 #(.width(width)) rd_st3_155  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[155]), .rdlo_in(a3_wr[219]),  .coef_in(coef[216]), .rdup_out(a4_wr[155]), .rdlo_out(a4_wr[219]));
			radix2 #(.width(width)) rd_st3_156  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[156]), .rdlo_in(a3_wr[220]),  .coef_in(coef[224]), .rdup_out(a4_wr[156]), .rdlo_out(a4_wr[220]));
			radix2 #(.width(width)) rd_st3_157  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[157]), .rdlo_in(a3_wr[221]),  .coef_in(coef[232]), .rdup_out(a4_wr[157]), .rdlo_out(a4_wr[221]));
			radix2 #(.width(width)) rd_st3_158  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[158]), .rdlo_in(a3_wr[222]),  .coef_in(coef[240]), .rdup_out(a4_wr[158]), .rdlo_out(a4_wr[222]));
			radix2 #(.width(width)) rd_st3_159  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[159]), .rdlo_in(a3_wr[223]),  .coef_in(coef[248]), .rdup_out(a4_wr[159]), .rdlo_out(a4_wr[223]));
			radix2 #(.width(width)) rd_st3_160  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[160]), .rdlo_in(a3_wr[224]),  .coef_in(coef[256]), .rdup_out(a4_wr[160]), .rdlo_out(a4_wr[224]));
			radix2 #(.width(width)) rd_st3_161  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[161]), .rdlo_in(a3_wr[225]),  .coef_in(coef[264]), .rdup_out(a4_wr[161]), .rdlo_out(a4_wr[225]));
			radix2 #(.width(width)) rd_st3_162  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[162]), .rdlo_in(a3_wr[226]),  .coef_in(coef[272]), .rdup_out(a4_wr[162]), .rdlo_out(a4_wr[226]));
			radix2 #(.width(width)) rd_st3_163  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[163]), .rdlo_in(a3_wr[227]),  .coef_in(coef[280]), .rdup_out(a4_wr[163]), .rdlo_out(a4_wr[227]));
			radix2 #(.width(width)) rd_st3_164  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[164]), .rdlo_in(a3_wr[228]),  .coef_in(coef[288]), .rdup_out(a4_wr[164]), .rdlo_out(a4_wr[228]));
			radix2 #(.width(width)) rd_st3_165  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[165]), .rdlo_in(a3_wr[229]),  .coef_in(coef[296]), .rdup_out(a4_wr[165]), .rdlo_out(a4_wr[229]));
			radix2 #(.width(width)) rd_st3_166  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[166]), .rdlo_in(a3_wr[230]),  .coef_in(coef[304]), .rdup_out(a4_wr[166]), .rdlo_out(a4_wr[230]));
			radix2 #(.width(width)) rd_st3_167  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[167]), .rdlo_in(a3_wr[231]),  .coef_in(coef[312]), .rdup_out(a4_wr[167]), .rdlo_out(a4_wr[231]));
			radix2 #(.width(width)) rd_st3_168  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[168]), .rdlo_in(a3_wr[232]),  .coef_in(coef[320]), .rdup_out(a4_wr[168]), .rdlo_out(a4_wr[232]));
			radix2 #(.width(width)) rd_st3_169  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[169]), .rdlo_in(a3_wr[233]),  .coef_in(coef[328]), .rdup_out(a4_wr[169]), .rdlo_out(a4_wr[233]));
			radix2 #(.width(width)) rd_st3_170  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[170]), .rdlo_in(a3_wr[234]),  .coef_in(coef[336]), .rdup_out(a4_wr[170]), .rdlo_out(a4_wr[234]));
			radix2 #(.width(width)) rd_st3_171  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[171]), .rdlo_in(a3_wr[235]),  .coef_in(coef[344]), .rdup_out(a4_wr[171]), .rdlo_out(a4_wr[235]));
			radix2 #(.width(width)) rd_st3_172  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[172]), .rdlo_in(a3_wr[236]),  .coef_in(coef[352]), .rdup_out(a4_wr[172]), .rdlo_out(a4_wr[236]));
			radix2 #(.width(width)) rd_st3_173  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[173]), .rdlo_in(a3_wr[237]),  .coef_in(coef[360]), .rdup_out(a4_wr[173]), .rdlo_out(a4_wr[237]));
			radix2 #(.width(width)) rd_st3_174  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[174]), .rdlo_in(a3_wr[238]),  .coef_in(coef[368]), .rdup_out(a4_wr[174]), .rdlo_out(a4_wr[238]));
			radix2 #(.width(width)) rd_st3_175  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[175]), .rdlo_in(a3_wr[239]),  .coef_in(coef[376]), .rdup_out(a4_wr[175]), .rdlo_out(a4_wr[239]));
			radix2 #(.width(width)) rd_st3_176  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[176]), .rdlo_in(a3_wr[240]),  .coef_in(coef[384]), .rdup_out(a4_wr[176]), .rdlo_out(a4_wr[240]));
			radix2 #(.width(width)) rd_st3_177  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[177]), .rdlo_in(a3_wr[241]),  .coef_in(coef[392]), .rdup_out(a4_wr[177]), .rdlo_out(a4_wr[241]));
			radix2 #(.width(width)) rd_st3_178  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[178]), .rdlo_in(a3_wr[242]),  .coef_in(coef[400]), .rdup_out(a4_wr[178]), .rdlo_out(a4_wr[242]));
			radix2 #(.width(width)) rd_st3_179  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[179]), .rdlo_in(a3_wr[243]),  .coef_in(coef[408]), .rdup_out(a4_wr[179]), .rdlo_out(a4_wr[243]));
			radix2 #(.width(width)) rd_st3_180  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[180]), .rdlo_in(a3_wr[244]),  .coef_in(coef[416]), .rdup_out(a4_wr[180]), .rdlo_out(a4_wr[244]));
			radix2 #(.width(width)) rd_st3_181  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[181]), .rdlo_in(a3_wr[245]),  .coef_in(coef[424]), .rdup_out(a4_wr[181]), .rdlo_out(a4_wr[245]));
			radix2 #(.width(width)) rd_st3_182  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[182]), .rdlo_in(a3_wr[246]),  .coef_in(coef[432]), .rdup_out(a4_wr[182]), .rdlo_out(a4_wr[246]));
			radix2 #(.width(width)) rd_st3_183  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[183]), .rdlo_in(a3_wr[247]),  .coef_in(coef[440]), .rdup_out(a4_wr[183]), .rdlo_out(a4_wr[247]));
			radix2 #(.width(width)) rd_st3_184  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[184]), .rdlo_in(a3_wr[248]),  .coef_in(coef[448]), .rdup_out(a4_wr[184]), .rdlo_out(a4_wr[248]));
			radix2 #(.width(width)) rd_st3_185  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[185]), .rdlo_in(a3_wr[249]),  .coef_in(coef[456]), .rdup_out(a4_wr[185]), .rdlo_out(a4_wr[249]));
			radix2 #(.width(width)) rd_st3_186  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[186]), .rdlo_in(a3_wr[250]),  .coef_in(coef[464]), .rdup_out(a4_wr[186]), .rdlo_out(a4_wr[250]));
			radix2 #(.width(width)) rd_st3_187  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[187]), .rdlo_in(a3_wr[251]),  .coef_in(coef[472]), .rdup_out(a4_wr[187]), .rdlo_out(a4_wr[251]));
			radix2 #(.width(width)) rd_st3_188  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[188]), .rdlo_in(a3_wr[252]),  .coef_in(coef[480]), .rdup_out(a4_wr[188]), .rdlo_out(a4_wr[252]));
			radix2 #(.width(width)) rd_st3_189  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[189]), .rdlo_in(a3_wr[253]),  .coef_in(coef[488]), .rdup_out(a4_wr[189]), .rdlo_out(a4_wr[253]));
			radix2 #(.width(width)) rd_st3_190  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[190]), .rdlo_in(a3_wr[254]),  .coef_in(coef[496]), .rdup_out(a4_wr[190]), .rdlo_out(a4_wr[254]));
			radix2 #(.width(width)) rd_st3_191  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[191]), .rdlo_in(a3_wr[255]),  .coef_in(coef[504]), .rdup_out(a4_wr[191]), .rdlo_out(a4_wr[255]));
			radix2 #(.width(width)) rd_st3_256  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[256]), .rdlo_in(a3_wr[320]),  .coef_in(coef[0]), .rdup_out(a4_wr[256]), .rdlo_out(a4_wr[320]));
			radix2 #(.width(width)) rd_st3_257  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[257]), .rdlo_in(a3_wr[321]),  .coef_in(coef[8]), .rdup_out(a4_wr[257]), .rdlo_out(a4_wr[321]));
			radix2 #(.width(width)) rd_st3_258  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[258]), .rdlo_in(a3_wr[322]),  .coef_in(coef[16]), .rdup_out(a4_wr[258]), .rdlo_out(a4_wr[322]));
			radix2 #(.width(width)) rd_st3_259  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[259]), .rdlo_in(a3_wr[323]),  .coef_in(coef[24]), .rdup_out(a4_wr[259]), .rdlo_out(a4_wr[323]));
			radix2 #(.width(width)) rd_st3_260  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[260]), .rdlo_in(a3_wr[324]),  .coef_in(coef[32]), .rdup_out(a4_wr[260]), .rdlo_out(a4_wr[324]));
			radix2 #(.width(width)) rd_st3_261  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[261]), .rdlo_in(a3_wr[325]),  .coef_in(coef[40]), .rdup_out(a4_wr[261]), .rdlo_out(a4_wr[325]));
			radix2 #(.width(width)) rd_st3_262  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[262]), .rdlo_in(a3_wr[326]),  .coef_in(coef[48]), .rdup_out(a4_wr[262]), .rdlo_out(a4_wr[326]));
			radix2 #(.width(width)) rd_st3_263  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[263]), .rdlo_in(a3_wr[327]),  .coef_in(coef[56]), .rdup_out(a4_wr[263]), .rdlo_out(a4_wr[327]));
			radix2 #(.width(width)) rd_st3_264  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[264]), .rdlo_in(a3_wr[328]),  .coef_in(coef[64]), .rdup_out(a4_wr[264]), .rdlo_out(a4_wr[328]));
			radix2 #(.width(width)) rd_st3_265  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[265]), .rdlo_in(a3_wr[329]),  .coef_in(coef[72]), .rdup_out(a4_wr[265]), .rdlo_out(a4_wr[329]));
			radix2 #(.width(width)) rd_st3_266  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[266]), .rdlo_in(a3_wr[330]),  .coef_in(coef[80]), .rdup_out(a4_wr[266]), .rdlo_out(a4_wr[330]));
			radix2 #(.width(width)) rd_st3_267  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[267]), .rdlo_in(a3_wr[331]),  .coef_in(coef[88]), .rdup_out(a4_wr[267]), .rdlo_out(a4_wr[331]));
			radix2 #(.width(width)) rd_st3_268  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[268]), .rdlo_in(a3_wr[332]),  .coef_in(coef[96]), .rdup_out(a4_wr[268]), .rdlo_out(a4_wr[332]));
			radix2 #(.width(width)) rd_st3_269  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[269]), .rdlo_in(a3_wr[333]),  .coef_in(coef[104]), .rdup_out(a4_wr[269]), .rdlo_out(a4_wr[333]));
			radix2 #(.width(width)) rd_st3_270  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[270]), .rdlo_in(a3_wr[334]),  .coef_in(coef[112]), .rdup_out(a4_wr[270]), .rdlo_out(a4_wr[334]));
			radix2 #(.width(width)) rd_st3_271  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[271]), .rdlo_in(a3_wr[335]),  .coef_in(coef[120]), .rdup_out(a4_wr[271]), .rdlo_out(a4_wr[335]));
			radix2 #(.width(width)) rd_st3_272  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[272]), .rdlo_in(a3_wr[336]),  .coef_in(coef[128]), .rdup_out(a4_wr[272]), .rdlo_out(a4_wr[336]));
			radix2 #(.width(width)) rd_st3_273  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[273]), .rdlo_in(a3_wr[337]),  .coef_in(coef[136]), .rdup_out(a4_wr[273]), .rdlo_out(a4_wr[337]));
			radix2 #(.width(width)) rd_st3_274  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[274]), .rdlo_in(a3_wr[338]),  .coef_in(coef[144]), .rdup_out(a4_wr[274]), .rdlo_out(a4_wr[338]));
			radix2 #(.width(width)) rd_st3_275  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[275]), .rdlo_in(a3_wr[339]),  .coef_in(coef[152]), .rdup_out(a4_wr[275]), .rdlo_out(a4_wr[339]));
			radix2 #(.width(width)) rd_st3_276  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[276]), .rdlo_in(a3_wr[340]),  .coef_in(coef[160]), .rdup_out(a4_wr[276]), .rdlo_out(a4_wr[340]));
			radix2 #(.width(width)) rd_st3_277  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[277]), .rdlo_in(a3_wr[341]),  .coef_in(coef[168]), .rdup_out(a4_wr[277]), .rdlo_out(a4_wr[341]));
			radix2 #(.width(width)) rd_st3_278  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[278]), .rdlo_in(a3_wr[342]),  .coef_in(coef[176]), .rdup_out(a4_wr[278]), .rdlo_out(a4_wr[342]));
			radix2 #(.width(width)) rd_st3_279  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[279]), .rdlo_in(a3_wr[343]),  .coef_in(coef[184]), .rdup_out(a4_wr[279]), .rdlo_out(a4_wr[343]));
			radix2 #(.width(width)) rd_st3_280  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[280]), .rdlo_in(a3_wr[344]),  .coef_in(coef[192]), .rdup_out(a4_wr[280]), .rdlo_out(a4_wr[344]));
			radix2 #(.width(width)) rd_st3_281  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[281]), .rdlo_in(a3_wr[345]),  .coef_in(coef[200]), .rdup_out(a4_wr[281]), .rdlo_out(a4_wr[345]));
			radix2 #(.width(width)) rd_st3_282  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[282]), .rdlo_in(a3_wr[346]),  .coef_in(coef[208]), .rdup_out(a4_wr[282]), .rdlo_out(a4_wr[346]));
			radix2 #(.width(width)) rd_st3_283  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[283]), .rdlo_in(a3_wr[347]),  .coef_in(coef[216]), .rdup_out(a4_wr[283]), .rdlo_out(a4_wr[347]));
			radix2 #(.width(width)) rd_st3_284  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[284]), .rdlo_in(a3_wr[348]),  .coef_in(coef[224]), .rdup_out(a4_wr[284]), .rdlo_out(a4_wr[348]));
			radix2 #(.width(width)) rd_st3_285  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[285]), .rdlo_in(a3_wr[349]),  .coef_in(coef[232]), .rdup_out(a4_wr[285]), .rdlo_out(a4_wr[349]));
			radix2 #(.width(width)) rd_st3_286  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[286]), .rdlo_in(a3_wr[350]),  .coef_in(coef[240]), .rdup_out(a4_wr[286]), .rdlo_out(a4_wr[350]));
			radix2 #(.width(width)) rd_st3_287  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[287]), .rdlo_in(a3_wr[351]),  .coef_in(coef[248]), .rdup_out(a4_wr[287]), .rdlo_out(a4_wr[351]));
			radix2 #(.width(width)) rd_st3_288  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[288]), .rdlo_in(a3_wr[352]),  .coef_in(coef[256]), .rdup_out(a4_wr[288]), .rdlo_out(a4_wr[352]));
			radix2 #(.width(width)) rd_st3_289  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[289]), .rdlo_in(a3_wr[353]),  .coef_in(coef[264]), .rdup_out(a4_wr[289]), .rdlo_out(a4_wr[353]));
			radix2 #(.width(width)) rd_st3_290  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[290]), .rdlo_in(a3_wr[354]),  .coef_in(coef[272]), .rdup_out(a4_wr[290]), .rdlo_out(a4_wr[354]));
			radix2 #(.width(width)) rd_st3_291  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[291]), .rdlo_in(a3_wr[355]),  .coef_in(coef[280]), .rdup_out(a4_wr[291]), .rdlo_out(a4_wr[355]));
			radix2 #(.width(width)) rd_st3_292  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[292]), .rdlo_in(a3_wr[356]),  .coef_in(coef[288]), .rdup_out(a4_wr[292]), .rdlo_out(a4_wr[356]));
			radix2 #(.width(width)) rd_st3_293  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[293]), .rdlo_in(a3_wr[357]),  .coef_in(coef[296]), .rdup_out(a4_wr[293]), .rdlo_out(a4_wr[357]));
			radix2 #(.width(width)) rd_st3_294  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[294]), .rdlo_in(a3_wr[358]),  .coef_in(coef[304]), .rdup_out(a4_wr[294]), .rdlo_out(a4_wr[358]));
			radix2 #(.width(width)) rd_st3_295  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[295]), .rdlo_in(a3_wr[359]),  .coef_in(coef[312]), .rdup_out(a4_wr[295]), .rdlo_out(a4_wr[359]));
			radix2 #(.width(width)) rd_st3_296  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[296]), .rdlo_in(a3_wr[360]),  .coef_in(coef[320]), .rdup_out(a4_wr[296]), .rdlo_out(a4_wr[360]));
			radix2 #(.width(width)) rd_st3_297  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[297]), .rdlo_in(a3_wr[361]),  .coef_in(coef[328]), .rdup_out(a4_wr[297]), .rdlo_out(a4_wr[361]));
			radix2 #(.width(width)) rd_st3_298  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[298]), .rdlo_in(a3_wr[362]),  .coef_in(coef[336]), .rdup_out(a4_wr[298]), .rdlo_out(a4_wr[362]));
			radix2 #(.width(width)) rd_st3_299  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[299]), .rdlo_in(a3_wr[363]),  .coef_in(coef[344]), .rdup_out(a4_wr[299]), .rdlo_out(a4_wr[363]));
			radix2 #(.width(width)) rd_st3_300  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[300]), .rdlo_in(a3_wr[364]),  .coef_in(coef[352]), .rdup_out(a4_wr[300]), .rdlo_out(a4_wr[364]));
			radix2 #(.width(width)) rd_st3_301  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[301]), .rdlo_in(a3_wr[365]),  .coef_in(coef[360]), .rdup_out(a4_wr[301]), .rdlo_out(a4_wr[365]));
			radix2 #(.width(width)) rd_st3_302  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[302]), .rdlo_in(a3_wr[366]),  .coef_in(coef[368]), .rdup_out(a4_wr[302]), .rdlo_out(a4_wr[366]));
			radix2 #(.width(width)) rd_st3_303  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[303]), .rdlo_in(a3_wr[367]),  .coef_in(coef[376]), .rdup_out(a4_wr[303]), .rdlo_out(a4_wr[367]));
			radix2 #(.width(width)) rd_st3_304  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[304]), .rdlo_in(a3_wr[368]),  .coef_in(coef[384]), .rdup_out(a4_wr[304]), .rdlo_out(a4_wr[368]));
			radix2 #(.width(width)) rd_st3_305  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[305]), .rdlo_in(a3_wr[369]),  .coef_in(coef[392]), .rdup_out(a4_wr[305]), .rdlo_out(a4_wr[369]));
			radix2 #(.width(width)) rd_st3_306  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[306]), .rdlo_in(a3_wr[370]),  .coef_in(coef[400]), .rdup_out(a4_wr[306]), .rdlo_out(a4_wr[370]));
			radix2 #(.width(width)) rd_st3_307  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[307]), .rdlo_in(a3_wr[371]),  .coef_in(coef[408]), .rdup_out(a4_wr[307]), .rdlo_out(a4_wr[371]));
			radix2 #(.width(width)) rd_st3_308  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[308]), .rdlo_in(a3_wr[372]),  .coef_in(coef[416]), .rdup_out(a4_wr[308]), .rdlo_out(a4_wr[372]));
			radix2 #(.width(width)) rd_st3_309  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[309]), .rdlo_in(a3_wr[373]),  .coef_in(coef[424]), .rdup_out(a4_wr[309]), .rdlo_out(a4_wr[373]));
			radix2 #(.width(width)) rd_st3_310  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[310]), .rdlo_in(a3_wr[374]),  .coef_in(coef[432]), .rdup_out(a4_wr[310]), .rdlo_out(a4_wr[374]));
			radix2 #(.width(width)) rd_st3_311  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[311]), .rdlo_in(a3_wr[375]),  .coef_in(coef[440]), .rdup_out(a4_wr[311]), .rdlo_out(a4_wr[375]));
			radix2 #(.width(width)) rd_st3_312  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[312]), .rdlo_in(a3_wr[376]),  .coef_in(coef[448]), .rdup_out(a4_wr[312]), .rdlo_out(a4_wr[376]));
			radix2 #(.width(width)) rd_st3_313  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[313]), .rdlo_in(a3_wr[377]),  .coef_in(coef[456]), .rdup_out(a4_wr[313]), .rdlo_out(a4_wr[377]));
			radix2 #(.width(width)) rd_st3_314  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[314]), .rdlo_in(a3_wr[378]),  .coef_in(coef[464]), .rdup_out(a4_wr[314]), .rdlo_out(a4_wr[378]));
			radix2 #(.width(width)) rd_st3_315  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[315]), .rdlo_in(a3_wr[379]),  .coef_in(coef[472]), .rdup_out(a4_wr[315]), .rdlo_out(a4_wr[379]));
			radix2 #(.width(width)) rd_st3_316  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[316]), .rdlo_in(a3_wr[380]),  .coef_in(coef[480]), .rdup_out(a4_wr[316]), .rdlo_out(a4_wr[380]));
			radix2 #(.width(width)) rd_st3_317  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[317]), .rdlo_in(a3_wr[381]),  .coef_in(coef[488]), .rdup_out(a4_wr[317]), .rdlo_out(a4_wr[381]));
			radix2 #(.width(width)) rd_st3_318  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[318]), .rdlo_in(a3_wr[382]),  .coef_in(coef[496]), .rdup_out(a4_wr[318]), .rdlo_out(a4_wr[382]));
			radix2 #(.width(width)) rd_st3_319  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[319]), .rdlo_in(a3_wr[383]),  .coef_in(coef[504]), .rdup_out(a4_wr[319]), .rdlo_out(a4_wr[383]));
			radix2 #(.width(width)) rd_st3_384  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[384]), .rdlo_in(a3_wr[448]),  .coef_in(coef[0]), .rdup_out(a4_wr[384]), .rdlo_out(a4_wr[448]));
			radix2 #(.width(width)) rd_st3_385  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[385]), .rdlo_in(a3_wr[449]),  .coef_in(coef[8]), .rdup_out(a4_wr[385]), .rdlo_out(a4_wr[449]));
			radix2 #(.width(width)) rd_st3_386  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[386]), .rdlo_in(a3_wr[450]),  .coef_in(coef[16]), .rdup_out(a4_wr[386]), .rdlo_out(a4_wr[450]));
			radix2 #(.width(width)) rd_st3_387  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[387]), .rdlo_in(a3_wr[451]),  .coef_in(coef[24]), .rdup_out(a4_wr[387]), .rdlo_out(a4_wr[451]));
			radix2 #(.width(width)) rd_st3_388  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[388]), .rdlo_in(a3_wr[452]),  .coef_in(coef[32]), .rdup_out(a4_wr[388]), .rdlo_out(a4_wr[452]));
			radix2 #(.width(width)) rd_st3_389  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[389]), .rdlo_in(a3_wr[453]),  .coef_in(coef[40]), .rdup_out(a4_wr[389]), .rdlo_out(a4_wr[453]));
			radix2 #(.width(width)) rd_st3_390  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[390]), .rdlo_in(a3_wr[454]),  .coef_in(coef[48]), .rdup_out(a4_wr[390]), .rdlo_out(a4_wr[454]));
			radix2 #(.width(width)) rd_st3_391  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[391]), .rdlo_in(a3_wr[455]),  .coef_in(coef[56]), .rdup_out(a4_wr[391]), .rdlo_out(a4_wr[455]));
			radix2 #(.width(width)) rd_st3_392  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[392]), .rdlo_in(a3_wr[456]),  .coef_in(coef[64]), .rdup_out(a4_wr[392]), .rdlo_out(a4_wr[456]));
			radix2 #(.width(width)) rd_st3_393  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[393]), .rdlo_in(a3_wr[457]),  .coef_in(coef[72]), .rdup_out(a4_wr[393]), .rdlo_out(a4_wr[457]));
			radix2 #(.width(width)) rd_st3_394  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[394]), .rdlo_in(a3_wr[458]),  .coef_in(coef[80]), .rdup_out(a4_wr[394]), .rdlo_out(a4_wr[458]));
			radix2 #(.width(width)) rd_st3_395  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[395]), .rdlo_in(a3_wr[459]),  .coef_in(coef[88]), .rdup_out(a4_wr[395]), .rdlo_out(a4_wr[459]));
			radix2 #(.width(width)) rd_st3_396  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[396]), .rdlo_in(a3_wr[460]),  .coef_in(coef[96]), .rdup_out(a4_wr[396]), .rdlo_out(a4_wr[460]));
			radix2 #(.width(width)) rd_st3_397  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[397]), .rdlo_in(a3_wr[461]),  .coef_in(coef[104]), .rdup_out(a4_wr[397]), .rdlo_out(a4_wr[461]));
			radix2 #(.width(width)) rd_st3_398  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[398]), .rdlo_in(a3_wr[462]),  .coef_in(coef[112]), .rdup_out(a4_wr[398]), .rdlo_out(a4_wr[462]));
			radix2 #(.width(width)) rd_st3_399  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[399]), .rdlo_in(a3_wr[463]),  .coef_in(coef[120]), .rdup_out(a4_wr[399]), .rdlo_out(a4_wr[463]));
			radix2 #(.width(width)) rd_st3_400  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[400]), .rdlo_in(a3_wr[464]),  .coef_in(coef[128]), .rdup_out(a4_wr[400]), .rdlo_out(a4_wr[464]));
			radix2 #(.width(width)) rd_st3_401  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[401]), .rdlo_in(a3_wr[465]),  .coef_in(coef[136]), .rdup_out(a4_wr[401]), .rdlo_out(a4_wr[465]));
			radix2 #(.width(width)) rd_st3_402  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[402]), .rdlo_in(a3_wr[466]),  .coef_in(coef[144]), .rdup_out(a4_wr[402]), .rdlo_out(a4_wr[466]));
			radix2 #(.width(width)) rd_st3_403  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[403]), .rdlo_in(a3_wr[467]),  .coef_in(coef[152]), .rdup_out(a4_wr[403]), .rdlo_out(a4_wr[467]));
			radix2 #(.width(width)) rd_st3_404  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[404]), .rdlo_in(a3_wr[468]),  .coef_in(coef[160]), .rdup_out(a4_wr[404]), .rdlo_out(a4_wr[468]));
			radix2 #(.width(width)) rd_st3_405  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[405]), .rdlo_in(a3_wr[469]),  .coef_in(coef[168]), .rdup_out(a4_wr[405]), .rdlo_out(a4_wr[469]));
			radix2 #(.width(width)) rd_st3_406  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[406]), .rdlo_in(a3_wr[470]),  .coef_in(coef[176]), .rdup_out(a4_wr[406]), .rdlo_out(a4_wr[470]));
			radix2 #(.width(width)) rd_st3_407  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[407]), .rdlo_in(a3_wr[471]),  .coef_in(coef[184]), .rdup_out(a4_wr[407]), .rdlo_out(a4_wr[471]));
			radix2 #(.width(width)) rd_st3_408  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[408]), .rdlo_in(a3_wr[472]),  .coef_in(coef[192]), .rdup_out(a4_wr[408]), .rdlo_out(a4_wr[472]));
			radix2 #(.width(width)) rd_st3_409  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[409]), .rdlo_in(a3_wr[473]),  .coef_in(coef[200]), .rdup_out(a4_wr[409]), .rdlo_out(a4_wr[473]));
			radix2 #(.width(width)) rd_st3_410  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[410]), .rdlo_in(a3_wr[474]),  .coef_in(coef[208]), .rdup_out(a4_wr[410]), .rdlo_out(a4_wr[474]));
			radix2 #(.width(width)) rd_st3_411  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[411]), .rdlo_in(a3_wr[475]),  .coef_in(coef[216]), .rdup_out(a4_wr[411]), .rdlo_out(a4_wr[475]));
			radix2 #(.width(width)) rd_st3_412  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[412]), .rdlo_in(a3_wr[476]),  .coef_in(coef[224]), .rdup_out(a4_wr[412]), .rdlo_out(a4_wr[476]));
			radix2 #(.width(width)) rd_st3_413  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[413]), .rdlo_in(a3_wr[477]),  .coef_in(coef[232]), .rdup_out(a4_wr[413]), .rdlo_out(a4_wr[477]));
			radix2 #(.width(width)) rd_st3_414  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[414]), .rdlo_in(a3_wr[478]),  .coef_in(coef[240]), .rdup_out(a4_wr[414]), .rdlo_out(a4_wr[478]));
			radix2 #(.width(width)) rd_st3_415  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[415]), .rdlo_in(a3_wr[479]),  .coef_in(coef[248]), .rdup_out(a4_wr[415]), .rdlo_out(a4_wr[479]));
			radix2 #(.width(width)) rd_st3_416  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[416]), .rdlo_in(a3_wr[480]),  .coef_in(coef[256]), .rdup_out(a4_wr[416]), .rdlo_out(a4_wr[480]));
			radix2 #(.width(width)) rd_st3_417  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[417]), .rdlo_in(a3_wr[481]),  .coef_in(coef[264]), .rdup_out(a4_wr[417]), .rdlo_out(a4_wr[481]));
			radix2 #(.width(width)) rd_st3_418  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[418]), .rdlo_in(a3_wr[482]),  .coef_in(coef[272]), .rdup_out(a4_wr[418]), .rdlo_out(a4_wr[482]));
			radix2 #(.width(width)) rd_st3_419  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[419]), .rdlo_in(a3_wr[483]),  .coef_in(coef[280]), .rdup_out(a4_wr[419]), .rdlo_out(a4_wr[483]));
			radix2 #(.width(width)) rd_st3_420  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[420]), .rdlo_in(a3_wr[484]),  .coef_in(coef[288]), .rdup_out(a4_wr[420]), .rdlo_out(a4_wr[484]));
			radix2 #(.width(width)) rd_st3_421  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[421]), .rdlo_in(a3_wr[485]),  .coef_in(coef[296]), .rdup_out(a4_wr[421]), .rdlo_out(a4_wr[485]));
			radix2 #(.width(width)) rd_st3_422  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[422]), .rdlo_in(a3_wr[486]),  .coef_in(coef[304]), .rdup_out(a4_wr[422]), .rdlo_out(a4_wr[486]));
			radix2 #(.width(width)) rd_st3_423  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[423]), .rdlo_in(a3_wr[487]),  .coef_in(coef[312]), .rdup_out(a4_wr[423]), .rdlo_out(a4_wr[487]));
			radix2 #(.width(width)) rd_st3_424  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[424]), .rdlo_in(a3_wr[488]),  .coef_in(coef[320]), .rdup_out(a4_wr[424]), .rdlo_out(a4_wr[488]));
			radix2 #(.width(width)) rd_st3_425  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[425]), .rdlo_in(a3_wr[489]),  .coef_in(coef[328]), .rdup_out(a4_wr[425]), .rdlo_out(a4_wr[489]));
			radix2 #(.width(width)) rd_st3_426  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[426]), .rdlo_in(a3_wr[490]),  .coef_in(coef[336]), .rdup_out(a4_wr[426]), .rdlo_out(a4_wr[490]));
			radix2 #(.width(width)) rd_st3_427  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[427]), .rdlo_in(a3_wr[491]),  .coef_in(coef[344]), .rdup_out(a4_wr[427]), .rdlo_out(a4_wr[491]));
			radix2 #(.width(width)) rd_st3_428  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[428]), .rdlo_in(a3_wr[492]),  .coef_in(coef[352]), .rdup_out(a4_wr[428]), .rdlo_out(a4_wr[492]));
			radix2 #(.width(width)) rd_st3_429  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[429]), .rdlo_in(a3_wr[493]),  .coef_in(coef[360]), .rdup_out(a4_wr[429]), .rdlo_out(a4_wr[493]));
			radix2 #(.width(width)) rd_st3_430  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[430]), .rdlo_in(a3_wr[494]),  .coef_in(coef[368]), .rdup_out(a4_wr[430]), .rdlo_out(a4_wr[494]));
			radix2 #(.width(width)) rd_st3_431  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[431]), .rdlo_in(a3_wr[495]),  .coef_in(coef[376]), .rdup_out(a4_wr[431]), .rdlo_out(a4_wr[495]));
			radix2 #(.width(width)) rd_st3_432  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[432]), .rdlo_in(a3_wr[496]),  .coef_in(coef[384]), .rdup_out(a4_wr[432]), .rdlo_out(a4_wr[496]));
			radix2 #(.width(width)) rd_st3_433  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[433]), .rdlo_in(a3_wr[497]),  .coef_in(coef[392]), .rdup_out(a4_wr[433]), .rdlo_out(a4_wr[497]));
			radix2 #(.width(width)) rd_st3_434  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[434]), .rdlo_in(a3_wr[498]),  .coef_in(coef[400]), .rdup_out(a4_wr[434]), .rdlo_out(a4_wr[498]));
			radix2 #(.width(width)) rd_st3_435  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[435]), .rdlo_in(a3_wr[499]),  .coef_in(coef[408]), .rdup_out(a4_wr[435]), .rdlo_out(a4_wr[499]));
			radix2 #(.width(width)) rd_st3_436  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[436]), .rdlo_in(a3_wr[500]),  .coef_in(coef[416]), .rdup_out(a4_wr[436]), .rdlo_out(a4_wr[500]));
			radix2 #(.width(width)) rd_st3_437  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[437]), .rdlo_in(a3_wr[501]),  .coef_in(coef[424]), .rdup_out(a4_wr[437]), .rdlo_out(a4_wr[501]));
			radix2 #(.width(width)) rd_st3_438  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[438]), .rdlo_in(a3_wr[502]),  .coef_in(coef[432]), .rdup_out(a4_wr[438]), .rdlo_out(a4_wr[502]));
			radix2 #(.width(width)) rd_st3_439  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[439]), .rdlo_in(a3_wr[503]),  .coef_in(coef[440]), .rdup_out(a4_wr[439]), .rdlo_out(a4_wr[503]));
			radix2 #(.width(width)) rd_st3_440  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[440]), .rdlo_in(a3_wr[504]),  .coef_in(coef[448]), .rdup_out(a4_wr[440]), .rdlo_out(a4_wr[504]));
			radix2 #(.width(width)) rd_st3_441  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[441]), .rdlo_in(a3_wr[505]),  .coef_in(coef[456]), .rdup_out(a4_wr[441]), .rdlo_out(a4_wr[505]));
			radix2 #(.width(width)) rd_st3_442  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[442]), .rdlo_in(a3_wr[506]),  .coef_in(coef[464]), .rdup_out(a4_wr[442]), .rdlo_out(a4_wr[506]));
			radix2 #(.width(width)) rd_st3_443  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[443]), .rdlo_in(a3_wr[507]),  .coef_in(coef[472]), .rdup_out(a4_wr[443]), .rdlo_out(a4_wr[507]));
			radix2 #(.width(width)) rd_st3_444  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[444]), .rdlo_in(a3_wr[508]),  .coef_in(coef[480]), .rdup_out(a4_wr[444]), .rdlo_out(a4_wr[508]));
			radix2 #(.width(width)) rd_st3_445  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[445]), .rdlo_in(a3_wr[509]),  .coef_in(coef[488]), .rdup_out(a4_wr[445]), .rdlo_out(a4_wr[509]));
			radix2 #(.width(width)) rd_st3_446  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[446]), .rdlo_in(a3_wr[510]),  .coef_in(coef[496]), .rdup_out(a4_wr[446]), .rdlo_out(a4_wr[510]));
			radix2 #(.width(width)) rd_st3_447  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[447]), .rdlo_in(a3_wr[511]),  .coef_in(coef[504]), .rdup_out(a4_wr[447]), .rdlo_out(a4_wr[511]));
			radix2 #(.width(width)) rd_st3_512  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[512]), .rdlo_in(a3_wr[576]),  .coef_in(coef[0]), .rdup_out(a4_wr[512]), .rdlo_out(a4_wr[576]));
			radix2 #(.width(width)) rd_st3_513  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[513]), .rdlo_in(a3_wr[577]),  .coef_in(coef[8]), .rdup_out(a4_wr[513]), .rdlo_out(a4_wr[577]));
			radix2 #(.width(width)) rd_st3_514  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[514]), .rdlo_in(a3_wr[578]),  .coef_in(coef[16]), .rdup_out(a4_wr[514]), .rdlo_out(a4_wr[578]));
			radix2 #(.width(width)) rd_st3_515  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[515]), .rdlo_in(a3_wr[579]),  .coef_in(coef[24]), .rdup_out(a4_wr[515]), .rdlo_out(a4_wr[579]));
			radix2 #(.width(width)) rd_st3_516  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[516]), .rdlo_in(a3_wr[580]),  .coef_in(coef[32]), .rdup_out(a4_wr[516]), .rdlo_out(a4_wr[580]));
			radix2 #(.width(width)) rd_st3_517  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[517]), .rdlo_in(a3_wr[581]),  .coef_in(coef[40]), .rdup_out(a4_wr[517]), .rdlo_out(a4_wr[581]));
			radix2 #(.width(width)) rd_st3_518  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[518]), .rdlo_in(a3_wr[582]),  .coef_in(coef[48]), .rdup_out(a4_wr[518]), .rdlo_out(a4_wr[582]));
			radix2 #(.width(width)) rd_st3_519  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[519]), .rdlo_in(a3_wr[583]),  .coef_in(coef[56]), .rdup_out(a4_wr[519]), .rdlo_out(a4_wr[583]));
			radix2 #(.width(width)) rd_st3_520  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[520]), .rdlo_in(a3_wr[584]),  .coef_in(coef[64]), .rdup_out(a4_wr[520]), .rdlo_out(a4_wr[584]));
			radix2 #(.width(width)) rd_st3_521  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[521]), .rdlo_in(a3_wr[585]),  .coef_in(coef[72]), .rdup_out(a4_wr[521]), .rdlo_out(a4_wr[585]));
			radix2 #(.width(width)) rd_st3_522  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[522]), .rdlo_in(a3_wr[586]),  .coef_in(coef[80]), .rdup_out(a4_wr[522]), .rdlo_out(a4_wr[586]));
			radix2 #(.width(width)) rd_st3_523  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[523]), .rdlo_in(a3_wr[587]),  .coef_in(coef[88]), .rdup_out(a4_wr[523]), .rdlo_out(a4_wr[587]));
			radix2 #(.width(width)) rd_st3_524  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[524]), .rdlo_in(a3_wr[588]),  .coef_in(coef[96]), .rdup_out(a4_wr[524]), .rdlo_out(a4_wr[588]));
			radix2 #(.width(width)) rd_st3_525  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[525]), .rdlo_in(a3_wr[589]),  .coef_in(coef[104]), .rdup_out(a4_wr[525]), .rdlo_out(a4_wr[589]));
			radix2 #(.width(width)) rd_st3_526  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[526]), .rdlo_in(a3_wr[590]),  .coef_in(coef[112]), .rdup_out(a4_wr[526]), .rdlo_out(a4_wr[590]));
			radix2 #(.width(width)) rd_st3_527  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[527]), .rdlo_in(a3_wr[591]),  .coef_in(coef[120]), .rdup_out(a4_wr[527]), .rdlo_out(a4_wr[591]));
			radix2 #(.width(width)) rd_st3_528  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[528]), .rdlo_in(a3_wr[592]),  .coef_in(coef[128]), .rdup_out(a4_wr[528]), .rdlo_out(a4_wr[592]));
			radix2 #(.width(width)) rd_st3_529  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[529]), .rdlo_in(a3_wr[593]),  .coef_in(coef[136]), .rdup_out(a4_wr[529]), .rdlo_out(a4_wr[593]));
			radix2 #(.width(width)) rd_st3_530  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[530]), .rdlo_in(a3_wr[594]),  .coef_in(coef[144]), .rdup_out(a4_wr[530]), .rdlo_out(a4_wr[594]));
			radix2 #(.width(width)) rd_st3_531  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[531]), .rdlo_in(a3_wr[595]),  .coef_in(coef[152]), .rdup_out(a4_wr[531]), .rdlo_out(a4_wr[595]));
			radix2 #(.width(width)) rd_st3_532  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[532]), .rdlo_in(a3_wr[596]),  .coef_in(coef[160]), .rdup_out(a4_wr[532]), .rdlo_out(a4_wr[596]));
			radix2 #(.width(width)) rd_st3_533  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[533]), .rdlo_in(a3_wr[597]),  .coef_in(coef[168]), .rdup_out(a4_wr[533]), .rdlo_out(a4_wr[597]));
			radix2 #(.width(width)) rd_st3_534  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[534]), .rdlo_in(a3_wr[598]),  .coef_in(coef[176]), .rdup_out(a4_wr[534]), .rdlo_out(a4_wr[598]));
			radix2 #(.width(width)) rd_st3_535  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[535]), .rdlo_in(a3_wr[599]),  .coef_in(coef[184]), .rdup_out(a4_wr[535]), .rdlo_out(a4_wr[599]));
			radix2 #(.width(width)) rd_st3_536  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[536]), .rdlo_in(a3_wr[600]),  .coef_in(coef[192]), .rdup_out(a4_wr[536]), .rdlo_out(a4_wr[600]));
			radix2 #(.width(width)) rd_st3_537  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[537]), .rdlo_in(a3_wr[601]),  .coef_in(coef[200]), .rdup_out(a4_wr[537]), .rdlo_out(a4_wr[601]));
			radix2 #(.width(width)) rd_st3_538  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[538]), .rdlo_in(a3_wr[602]),  .coef_in(coef[208]), .rdup_out(a4_wr[538]), .rdlo_out(a4_wr[602]));
			radix2 #(.width(width)) rd_st3_539  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[539]), .rdlo_in(a3_wr[603]),  .coef_in(coef[216]), .rdup_out(a4_wr[539]), .rdlo_out(a4_wr[603]));
			radix2 #(.width(width)) rd_st3_540  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[540]), .rdlo_in(a3_wr[604]),  .coef_in(coef[224]), .rdup_out(a4_wr[540]), .rdlo_out(a4_wr[604]));
			radix2 #(.width(width)) rd_st3_541  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[541]), .rdlo_in(a3_wr[605]),  .coef_in(coef[232]), .rdup_out(a4_wr[541]), .rdlo_out(a4_wr[605]));
			radix2 #(.width(width)) rd_st3_542  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[542]), .rdlo_in(a3_wr[606]),  .coef_in(coef[240]), .rdup_out(a4_wr[542]), .rdlo_out(a4_wr[606]));
			radix2 #(.width(width)) rd_st3_543  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[543]), .rdlo_in(a3_wr[607]),  .coef_in(coef[248]), .rdup_out(a4_wr[543]), .rdlo_out(a4_wr[607]));
			radix2 #(.width(width)) rd_st3_544  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[544]), .rdlo_in(a3_wr[608]),  .coef_in(coef[256]), .rdup_out(a4_wr[544]), .rdlo_out(a4_wr[608]));
			radix2 #(.width(width)) rd_st3_545  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[545]), .rdlo_in(a3_wr[609]),  .coef_in(coef[264]), .rdup_out(a4_wr[545]), .rdlo_out(a4_wr[609]));
			radix2 #(.width(width)) rd_st3_546  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[546]), .rdlo_in(a3_wr[610]),  .coef_in(coef[272]), .rdup_out(a4_wr[546]), .rdlo_out(a4_wr[610]));
			radix2 #(.width(width)) rd_st3_547  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[547]), .rdlo_in(a3_wr[611]),  .coef_in(coef[280]), .rdup_out(a4_wr[547]), .rdlo_out(a4_wr[611]));
			radix2 #(.width(width)) rd_st3_548  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[548]), .rdlo_in(a3_wr[612]),  .coef_in(coef[288]), .rdup_out(a4_wr[548]), .rdlo_out(a4_wr[612]));
			radix2 #(.width(width)) rd_st3_549  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[549]), .rdlo_in(a3_wr[613]),  .coef_in(coef[296]), .rdup_out(a4_wr[549]), .rdlo_out(a4_wr[613]));
			radix2 #(.width(width)) rd_st3_550  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[550]), .rdlo_in(a3_wr[614]),  .coef_in(coef[304]), .rdup_out(a4_wr[550]), .rdlo_out(a4_wr[614]));
			radix2 #(.width(width)) rd_st3_551  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[551]), .rdlo_in(a3_wr[615]),  .coef_in(coef[312]), .rdup_out(a4_wr[551]), .rdlo_out(a4_wr[615]));
			radix2 #(.width(width)) rd_st3_552  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[552]), .rdlo_in(a3_wr[616]),  .coef_in(coef[320]), .rdup_out(a4_wr[552]), .rdlo_out(a4_wr[616]));
			radix2 #(.width(width)) rd_st3_553  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[553]), .rdlo_in(a3_wr[617]),  .coef_in(coef[328]), .rdup_out(a4_wr[553]), .rdlo_out(a4_wr[617]));
			radix2 #(.width(width)) rd_st3_554  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[554]), .rdlo_in(a3_wr[618]),  .coef_in(coef[336]), .rdup_out(a4_wr[554]), .rdlo_out(a4_wr[618]));
			radix2 #(.width(width)) rd_st3_555  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[555]), .rdlo_in(a3_wr[619]),  .coef_in(coef[344]), .rdup_out(a4_wr[555]), .rdlo_out(a4_wr[619]));
			radix2 #(.width(width)) rd_st3_556  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[556]), .rdlo_in(a3_wr[620]),  .coef_in(coef[352]), .rdup_out(a4_wr[556]), .rdlo_out(a4_wr[620]));
			radix2 #(.width(width)) rd_st3_557  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[557]), .rdlo_in(a3_wr[621]),  .coef_in(coef[360]), .rdup_out(a4_wr[557]), .rdlo_out(a4_wr[621]));
			radix2 #(.width(width)) rd_st3_558  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[558]), .rdlo_in(a3_wr[622]),  .coef_in(coef[368]), .rdup_out(a4_wr[558]), .rdlo_out(a4_wr[622]));
			radix2 #(.width(width)) rd_st3_559  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[559]), .rdlo_in(a3_wr[623]),  .coef_in(coef[376]), .rdup_out(a4_wr[559]), .rdlo_out(a4_wr[623]));
			radix2 #(.width(width)) rd_st3_560  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[560]), .rdlo_in(a3_wr[624]),  .coef_in(coef[384]), .rdup_out(a4_wr[560]), .rdlo_out(a4_wr[624]));
			radix2 #(.width(width)) rd_st3_561  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[561]), .rdlo_in(a3_wr[625]),  .coef_in(coef[392]), .rdup_out(a4_wr[561]), .rdlo_out(a4_wr[625]));
			radix2 #(.width(width)) rd_st3_562  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[562]), .rdlo_in(a3_wr[626]),  .coef_in(coef[400]), .rdup_out(a4_wr[562]), .rdlo_out(a4_wr[626]));
			radix2 #(.width(width)) rd_st3_563  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[563]), .rdlo_in(a3_wr[627]),  .coef_in(coef[408]), .rdup_out(a4_wr[563]), .rdlo_out(a4_wr[627]));
			radix2 #(.width(width)) rd_st3_564  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[564]), .rdlo_in(a3_wr[628]),  .coef_in(coef[416]), .rdup_out(a4_wr[564]), .rdlo_out(a4_wr[628]));
			radix2 #(.width(width)) rd_st3_565  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[565]), .rdlo_in(a3_wr[629]),  .coef_in(coef[424]), .rdup_out(a4_wr[565]), .rdlo_out(a4_wr[629]));
			radix2 #(.width(width)) rd_st3_566  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[566]), .rdlo_in(a3_wr[630]),  .coef_in(coef[432]), .rdup_out(a4_wr[566]), .rdlo_out(a4_wr[630]));
			radix2 #(.width(width)) rd_st3_567  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[567]), .rdlo_in(a3_wr[631]),  .coef_in(coef[440]), .rdup_out(a4_wr[567]), .rdlo_out(a4_wr[631]));
			radix2 #(.width(width)) rd_st3_568  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[568]), .rdlo_in(a3_wr[632]),  .coef_in(coef[448]), .rdup_out(a4_wr[568]), .rdlo_out(a4_wr[632]));
			radix2 #(.width(width)) rd_st3_569  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[569]), .rdlo_in(a3_wr[633]),  .coef_in(coef[456]), .rdup_out(a4_wr[569]), .rdlo_out(a4_wr[633]));
			radix2 #(.width(width)) rd_st3_570  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[570]), .rdlo_in(a3_wr[634]),  .coef_in(coef[464]), .rdup_out(a4_wr[570]), .rdlo_out(a4_wr[634]));
			radix2 #(.width(width)) rd_st3_571  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[571]), .rdlo_in(a3_wr[635]),  .coef_in(coef[472]), .rdup_out(a4_wr[571]), .rdlo_out(a4_wr[635]));
			radix2 #(.width(width)) rd_st3_572  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[572]), .rdlo_in(a3_wr[636]),  .coef_in(coef[480]), .rdup_out(a4_wr[572]), .rdlo_out(a4_wr[636]));
			radix2 #(.width(width)) rd_st3_573  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[573]), .rdlo_in(a3_wr[637]),  .coef_in(coef[488]), .rdup_out(a4_wr[573]), .rdlo_out(a4_wr[637]));
			radix2 #(.width(width)) rd_st3_574  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[574]), .rdlo_in(a3_wr[638]),  .coef_in(coef[496]), .rdup_out(a4_wr[574]), .rdlo_out(a4_wr[638]));
			radix2 #(.width(width)) rd_st3_575  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[575]), .rdlo_in(a3_wr[639]),  .coef_in(coef[504]), .rdup_out(a4_wr[575]), .rdlo_out(a4_wr[639]));
			radix2 #(.width(width)) rd_st3_640  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[640]), .rdlo_in(a3_wr[704]),  .coef_in(coef[0]), .rdup_out(a4_wr[640]), .rdlo_out(a4_wr[704]));
			radix2 #(.width(width)) rd_st3_641  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[641]), .rdlo_in(a3_wr[705]),  .coef_in(coef[8]), .rdup_out(a4_wr[641]), .rdlo_out(a4_wr[705]));
			radix2 #(.width(width)) rd_st3_642  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[642]), .rdlo_in(a3_wr[706]),  .coef_in(coef[16]), .rdup_out(a4_wr[642]), .rdlo_out(a4_wr[706]));
			radix2 #(.width(width)) rd_st3_643  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[643]), .rdlo_in(a3_wr[707]),  .coef_in(coef[24]), .rdup_out(a4_wr[643]), .rdlo_out(a4_wr[707]));
			radix2 #(.width(width)) rd_st3_644  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[644]), .rdlo_in(a3_wr[708]),  .coef_in(coef[32]), .rdup_out(a4_wr[644]), .rdlo_out(a4_wr[708]));
			radix2 #(.width(width)) rd_st3_645  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[645]), .rdlo_in(a3_wr[709]),  .coef_in(coef[40]), .rdup_out(a4_wr[645]), .rdlo_out(a4_wr[709]));
			radix2 #(.width(width)) rd_st3_646  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[646]), .rdlo_in(a3_wr[710]),  .coef_in(coef[48]), .rdup_out(a4_wr[646]), .rdlo_out(a4_wr[710]));
			radix2 #(.width(width)) rd_st3_647  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[647]), .rdlo_in(a3_wr[711]),  .coef_in(coef[56]), .rdup_out(a4_wr[647]), .rdlo_out(a4_wr[711]));
			radix2 #(.width(width)) rd_st3_648  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[648]), .rdlo_in(a3_wr[712]),  .coef_in(coef[64]), .rdup_out(a4_wr[648]), .rdlo_out(a4_wr[712]));
			radix2 #(.width(width)) rd_st3_649  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[649]), .rdlo_in(a3_wr[713]),  .coef_in(coef[72]), .rdup_out(a4_wr[649]), .rdlo_out(a4_wr[713]));
			radix2 #(.width(width)) rd_st3_650  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[650]), .rdlo_in(a3_wr[714]),  .coef_in(coef[80]), .rdup_out(a4_wr[650]), .rdlo_out(a4_wr[714]));
			radix2 #(.width(width)) rd_st3_651  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[651]), .rdlo_in(a3_wr[715]),  .coef_in(coef[88]), .rdup_out(a4_wr[651]), .rdlo_out(a4_wr[715]));
			radix2 #(.width(width)) rd_st3_652  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[652]), .rdlo_in(a3_wr[716]),  .coef_in(coef[96]), .rdup_out(a4_wr[652]), .rdlo_out(a4_wr[716]));
			radix2 #(.width(width)) rd_st3_653  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[653]), .rdlo_in(a3_wr[717]),  .coef_in(coef[104]), .rdup_out(a4_wr[653]), .rdlo_out(a4_wr[717]));
			radix2 #(.width(width)) rd_st3_654  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[654]), .rdlo_in(a3_wr[718]),  .coef_in(coef[112]), .rdup_out(a4_wr[654]), .rdlo_out(a4_wr[718]));
			radix2 #(.width(width)) rd_st3_655  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[655]), .rdlo_in(a3_wr[719]),  .coef_in(coef[120]), .rdup_out(a4_wr[655]), .rdlo_out(a4_wr[719]));
			radix2 #(.width(width)) rd_st3_656  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[656]), .rdlo_in(a3_wr[720]),  .coef_in(coef[128]), .rdup_out(a4_wr[656]), .rdlo_out(a4_wr[720]));
			radix2 #(.width(width)) rd_st3_657  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[657]), .rdlo_in(a3_wr[721]),  .coef_in(coef[136]), .rdup_out(a4_wr[657]), .rdlo_out(a4_wr[721]));
			radix2 #(.width(width)) rd_st3_658  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[658]), .rdlo_in(a3_wr[722]),  .coef_in(coef[144]), .rdup_out(a4_wr[658]), .rdlo_out(a4_wr[722]));
			radix2 #(.width(width)) rd_st3_659  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[659]), .rdlo_in(a3_wr[723]),  .coef_in(coef[152]), .rdup_out(a4_wr[659]), .rdlo_out(a4_wr[723]));
			radix2 #(.width(width)) rd_st3_660  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[660]), .rdlo_in(a3_wr[724]),  .coef_in(coef[160]), .rdup_out(a4_wr[660]), .rdlo_out(a4_wr[724]));
			radix2 #(.width(width)) rd_st3_661  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[661]), .rdlo_in(a3_wr[725]),  .coef_in(coef[168]), .rdup_out(a4_wr[661]), .rdlo_out(a4_wr[725]));
			radix2 #(.width(width)) rd_st3_662  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[662]), .rdlo_in(a3_wr[726]),  .coef_in(coef[176]), .rdup_out(a4_wr[662]), .rdlo_out(a4_wr[726]));
			radix2 #(.width(width)) rd_st3_663  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[663]), .rdlo_in(a3_wr[727]),  .coef_in(coef[184]), .rdup_out(a4_wr[663]), .rdlo_out(a4_wr[727]));
			radix2 #(.width(width)) rd_st3_664  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[664]), .rdlo_in(a3_wr[728]),  .coef_in(coef[192]), .rdup_out(a4_wr[664]), .rdlo_out(a4_wr[728]));
			radix2 #(.width(width)) rd_st3_665  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[665]), .rdlo_in(a3_wr[729]),  .coef_in(coef[200]), .rdup_out(a4_wr[665]), .rdlo_out(a4_wr[729]));
			radix2 #(.width(width)) rd_st3_666  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[666]), .rdlo_in(a3_wr[730]),  .coef_in(coef[208]), .rdup_out(a4_wr[666]), .rdlo_out(a4_wr[730]));
			radix2 #(.width(width)) rd_st3_667  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[667]), .rdlo_in(a3_wr[731]),  .coef_in(coef[216]), .rdup_out(a4_wr[667]), .rdlo_out(a4_wr[731]));
			radix2 #(.width(width)) rd_st3_668  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[668]), .rdlo_in(a3_wr[732]),  .coef_in(coef[224]), .rdup_out(a4_wr[668]), .rdlo_out(a4_wr[732]));
			radix2 #(.width(width)) rd_st3_669  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[669]), .rdlo_in(a3_wr[733]),  .coef_in(coef[232]), .rdup_out(a4_wr[669]), .rdlo_out(a4_wr[733]));
			radix2 #(.width(width)) rd_st3_670  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[670]), .rdlo_in(a3_wr[734]),  .coef_in(coef[240]), .rdup_out(a4_wr[670]), .rdlo_out(a4_wr[734]));
			radix2 #(.width(width)) rd_st3_671  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[671]), .rdlo_in(a3_wr[735]),  .coef_in(coef[248]), .rdup_out(a4_wr[671]), .rdlo_out(a4_wr[735]));
			radix2 #(.width(width)) rd_st3_672  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[672]), .rdlo_in(a3_wr[736]),  .coef_in(coef[256]), .rdup_out(a4_wr[672]), .rdlo_out(a4_wr[736]));
			radix2 #(.width(width)) rd_st3_673  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[673]), .rdlo_in(a3_wr[737]),  .coef_in(coef[264]), .rdup_out(a4_wr[673]), .rdlo_out(a4_wr[737]));
			radix2 #(.width(width)) rd_st3_674  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[674]), .rdlo_in(a3_wr[738]),  .coef_in(coef[272]), .rdup_out(a4_wr[674]), .rdlo_out(a4_wr[738]));
			radix2 #(.width(width)) rd_st3_675  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[675]), .rdlo_in(a3_wr[739]),  .coef_in(coef[280]), .rdup_out(a4_wr[675]), .rdlo_out(a4_wr[739]));
			radix2 #(.width(width)) rd_st3_676  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[676]), .rdlo_in(a3_wr[740]),  .coef_in(coef[288]), .rdup_out(a4_wr[676]), .rdlo_out(a4_wr[740]));
			radix2 #(.width(width)) rd_st3_677  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[677]), .rdlo_in(a3_wr[741]),  .coef_in(coef[296]), .rdup_out(a4_wr[677]), .rdlo_out(a4_wr[741]));
			radix2 #(.width(width)) rd_st3_678  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[678]), .rdlo_in(a3_wr[742]),  .coef_in(coef[304]), .rdup_out(a4_wr[678]), .rdlo_out(a4_wr[742]));
			radix2 #(.width(width)) rd_st3_679  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[679]), .rdlo_in(a3_wr[743]),  .coef_in(coef[312]), .rdup_out(a4_wr[679]), .rdlo_out(a4_wr[743]));
			radix2 #(.width(width)) rd_st3_680  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[680]), .rdlo_in(a3_wr[744]),  .coef_in(coef[320]), .rdup_out(a4_wr[680]), .rdlo_out(a4_wr[744]));
			radix2 #(.width(width)) rd_st3_681  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[681]), .rdlo_in(a3_wr[745]),  .coef_in(coef[328]), .rdup_out(a4_wr[681]), .rdlo_out(a4_wr[745]));
			radix2 #(.width(width)) rd_st3_682  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[682]), .rdlo_in(a3_wr[746]),  .coef_in(coef[336]), .rdup_out(a4_wr[682]), .rdlo_out(a4_wr[746]));
			radix2 #(.width(width)) rd_st3_683  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[683]), .rdlo_in(a3_wr[747]),  .coef_in(coef[344]), .rdup_out(a4_wr[683]), .rdlo_out(a4_wr[747]));
			radix2 #(.width(width)) rd_st3_684  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[684]), .rdlo_in(a3_wr[748]),  .coef_in(coef[352]), .rdup_out(a4_wr[684]), .rdlo_out(a4_wr[748]));
			radix2 #(.width(width)) rd_st3_685  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[685]), .rdlo_in(a3_wr[749]),  .coef_in(coef[360]), .rdup_out(a4_wr[685]), .rdlo_out(a4_wr[749]));
			radix2 #(.width(width)) rd_st3_686  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[686]), .rdlo_in(a3_wr[750]),  .coef_in(coef[368]), .rdup_out(a4_wr[686]), .rdlo_out(a4_wr[750]));
			radix2 #(.width(width)) rd_st3_687  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[687]), .rdlo_in(a3_wr[751]),  .coef_in(coef[376]), .rdup_out(a4_wr[687]), .rdlo_out(a4_wr[751]));
			radix2 #(.width(width)) rd_st3_688  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[688]), .rdlo_in(a3_wr[752]),  .coef_in(coef[384]), .rdup_out(a4_wr[688]), .rdlo_out(a4_wr[752]));
			radix2 #(.width(width)) rd_st3_689  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[689]), .rdlo_in(a3_wr[753]),  .coef_in(coef[392]), .rdup_out(a4_wr[689]), .rdlo_out(a4_wr[753]));
			radix2 #(.width(width)) rd_st3_690  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[690]), .rdlo_in(a3_wr[754]),  .coef_in(coef[400]), .rdup_out(a4_wr[690]), .rdlo_out(a4_wr[754]));
			radix2 #(.width(width)) rd_st3_691  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[691]), .rdlo_in(a3_wr[755]),  .coef_in(coef[408]), .rdup_out(a4_wr[691]), .rdlo_out(a4_wr[755]));
			radix2 #(.width(width)) rd_st3_692  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[692]), .rdlo_in(a3_wr[756]),  .coef_in(coef[416]), .rdup_out(a4_wr[692]), .rdlo_out(a4_wr[756]));
			radix2 #(.width(width)) rd_st3_693  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[693]), .rdlo_in(a3_wr[757]),  .coef_in(coef[424]), .rdup_out(a4_wr[693]), .rdlo_out(a4_wr[757]));
			radix2 #(.width(width)) rd_st3_694  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[694]), .rdlo_in(a3_wr[758]),  .coef_in(coef[432]), .rdup_out(a4_wr[694]), .rdlo_out(a4_wr[758]));
			radix2 #(.width(width)) rd_st3_695  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[695]), .rdlo_in(a3_wr[759]),  .coef_in(coef[440]), .rdup_out(a4_wr[695]), .rdlo_out(a4_wr[759]));
			radix2 #(.width(width)) rd_st3_696  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[696]), .rdlo_in(a3_wr[760]),  .coef_in(coef[448]), .rdup_out(a4_wr[696]), .rdlo_out(a4_wr[760]));
			radix2 #(.width(width)) rd_st3_697  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[697]), .rdlo_in(a3_wr[761]),  .coef_in(coef[456]), .rdup_out(a4_wr[697]), .rdlo_out(a4_wr[761]));
			radix2 #(.width(width)) rd_st3_698  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[698]), .rdlo_in(a3_wr[762]),  .coef_in(coef[464]), .rdup_out(a4_wr[698]), .rdlo_out(a4_wr[762]));
			radix2 #(.width(width)) rd_st3_699  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[699]), .rdlo_in(a3_wr[763]),  .coef_in(coef[472]), .rdup_out(a4_wr[699]), .rdlo_out(a4_wr[763]));
			radix2 #(.width(width)) rd_st3_700  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[700]), .rdlo_in(a3_wr[764]),  .coef_in(coef[480]), .rdup_out(a4_wr[700]), .rdlo_out(a4_wr[764]));
			radix2 #(.width(width)) rd_st3_701  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[701]), .rdlo_in(a3_wr[765]),  .coef_in(coef[488]), .rdup_out(a4_wr[701]), .rdlo_out(a4_wr[765]));
			radix2 #(.width(width)) rd_st3_702  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[702]), .rdlo_in(a3_wr[766]),  .coef_in(coef[496]), .rdup_out(a4_wr[702]), .rdlo_out(a4_wr[766]));
			radix2 #(.width(width)) rd_st3_703  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[703]), .rdlo_in(a3_wr[767]),  .coef_in(coef[504]), .rdup_out(a4_wr[703]), .rdlo_out(a4_wr[767]));
			radix2 #(.width(width)) rd_st3_768  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[768]), .rdlo_in(a3_wr[832]),  .coef_in(coef[0]), .rdup_out(a4_wr[768]), .rdlo_out(a4_wr[832]));
			radix2 #(.width(width)) rd_st3_769  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[769]), .rdlo_in(a3_wr[833]),  .coef_in(coef[8]), .rdup_out(a4_wr[769]), .rdlo_out(a4_wr[833]));
			radix2 #(.width(width)) rd_st3_770  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[770]), .rdlo_in(a3_wr[834]),  .coef_in(coef[16]), .rdup_out(a4_wr[770]), .rdlo_out(a4_wr[834]));
			radix2 #(.width(width)) rd_st3_771  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[771]), .rdlo_in(a3_wr[835]),  .coef_in(coef[24]), .rdup_out(a4_wr[771]), .rdlo_out(a4_wr[835]));
			radix2 #(.width(width)) rd_st3_772  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[772]), .rdlo_in(a3_wr[836]),  .coef_in(coef[32]), .rdup_out(a4_wr[772]), .rdlo_out(a4_wr[836]));
			radix2 #(.width(width)) rd_st3_773  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[773]), .rdlo_in(a3_wr[837]),  .coef_in(coef[40]), .rdup_out(a4_wr[773]), .rdlo_out(a4_wr[837]));
			radix2 #(.width(width)) rd_st3_774  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[774]), .rdlo_in(a3_wr[838]),  .coef_in(coef[48]), .rdup_out(a4_wr[774]), .rdlo_out(a4_wr[838]));
			radix2 #(.width(width)) rd_st3_775  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[775]), .rdlo_in(a3_wr[839]),  .coef_in(coef[56]), .rdup_out(a4_wr[775]), .rdlo_out(a4_wr[839]));
			radix2 #(.width(width)) rd_st3_776  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[776]), .rdlo_in(a3_wr[840]),  .coef_in(coef[64]), .rdup_out(a4_wr[776]), .rdlo_out(a4_wr[840]));
			radix2 #(.width(width)) rd_st3_777  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[777]), .rdlo_in(a3_wr[841]),  .coef_in(coef[72]), .rdup_out(a4_wr[777]), .rdlo_out(a4_wr[841]));
			radix2 #(.width(width)) rd_st3_778  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[778]), .rdlo_in(a3_wr[842]),  .coef_in(coef[80]), .rdup_out(a4_wr[778]), .rdlo_out(a4_wr[842]));
			radix2 #(.width(width)) rd_st3_779  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[779]), .rdlo_in(a3_wr[843]),  .coef_in(coef[88]), .rdup_out(a4_wr[779]), .rdlo_out(a4_wr[843]));
			radix2 #(.width(width)) rd_st3_780  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[780]), .rdlo_in(a3_wr[844]),  .coef_in(coef[96]), .rdup_out(a4_wr[780]), .rdlo_out(a4_wr[844]));
			radix2 #(.width(width)) rd_st3_781  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[781]), .rdlo_in(a3_wr[845]),  .coef_in(coef[104]), .rdup_out(a4_wr[781]), .rdlo_out(a4_wr[845]));
			radix2 #(.width(width)) rd_st3_782  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[782]), .rdlo_in(a3_wr[846]),  .coef_in(coef[112]), .rdup_out(a4_wr[782]), .rdlo_out(a4_wr[846]));
			radix2 #(.width(width)) rd_st3_783  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[783]), .rdlo_in(a3_wr[847]),  .coef_in(coef[120]), .rdup_out(a4_wr[783]), .rdlo_out(a4_wr[847]));
			radix2 #(.width(width)) rd_st3_784  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[784]), .rdlo_in(a3_wr[848]),  .coef_in(coef[128]), .rdup_out(a4_wr[784]), .rdlo_out(a4_wr[848]));
			radix2 #(.width(width)) rd_st3_785  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[785]), .rdlo_in(a3_wr[849]),  .coef_in(coef[136]), .rdup_out(a4_wr[785]), .rdlo_out(a4_wr[849]));
			radix2 #(.width(width)) rd_st3_786  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[786]), .rdlo_in(a3_wr[850]),  .coef_in(coef[144]), .rdup_out(a4_wr[786]), .rdlo_out(a4_wr[850]));
			radix2 #(.width(width)) rd_st3_787  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[787]), .rdlo_in(a3_wr[851]),  .coef_in(coef[152]), .rdup_out(a4_wr[787]), .rdlo_out(a4_wr[851]));
			radix2 #(.width(width)) rd_st3_788  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[788]), .rdlo_in(a3_wr[852]),  .coef_in(coef[160]), .rdup_out(a4_wr[788]), .rdlo_out(a4_wr[852]));
			radix2 #(.width(width)) rd_st3_789  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[789]), .rdlo_in(a3_wr[853]),  .coef_in(coef[168]), .rdup_out(a4_wr[789]), .rdlo_out(a4_wr[853]));
			radix2 #(.width(width)) rd_st3_790  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[790]), .rdlo_in(a3_wr[854]),  .coef_in(coef[176]), .rdup_out(a4_wr[790]), .rdlo_out(a4_wr[854]));
			radix2 #(.width(width)) rd_st3_791  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[791]), .rdlo_in(a3_wr[855]),  .coef_in(coef[184]), .rdup_out(a4_wr[791]), .rdlo_out(a4_wr[855]));
			radix2 #(.width(width)) rd_st3_792  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[792]), .rdlo_in(a3_wr[856]),  .coef_in(coef[192]), .rdup_out(a4_wr[792]), .rdlo_out(a4_wr[856]));
			radix2 #(.width(width)) rd_st3_793  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[793]), .rdlo_in(a3_wr[857]),  .coef_in(coef[200]), .rdup_out(a4_wr[793]), .rdlo_out(a4_wr[857]));
			radix2 #(.width(width)) rd_st3_794  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[794]), .rdlo_in(a3_wr[858]),  .coef_in(coef[208]), .rdup_out(a4_wr[794]), .rdlo_out(a4_wr[858]));
			radix2 #(.width(width)) rd_st3_795  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[795]), .rdlo_in(a3_wr[859]),  .coef_in(coef[216]), .rdup_out(a4_wr[795]), .rdlo_out(a4_wr[859]));
			radix2 #(.width(width)) rd_st3_796  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[796]), .rdlo_in(a3_wr[860]),  .coef_in(coef[224]), .rdup_out(a4_wr[796]), .rdlo_out(a4_wr[860]));
			radix2 #(.width(width)) rd_st3_797  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[797]), .rdlo_in(a3_wr[861]),  .coef_in(coef[232]), .rdup_out(a4_wr[797]), .rdlo_out(a4_wr[861]));
			radix2 #(.width(width)) rd_st3_798  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[798]), .rdlo_in(a3_wr[862]),  .coef_in(coef[240]), .rdup_out(a4_wr[798]), .rdlo_out(a4_wr[862]));
			radix2 #(.width(width)) rd_st3_799  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[799]), .rdlo_in(a3_wr[863]),  .coef_in(coef[248]), .rdup_out(a4_wr[799]), .rdlo_out(a4_wr[863]));
			radix2 #(.width(width)) rd_st3_800  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[800]), .rdlo_in(a3_wr[864]),  .coef_in(coef[256]), .rdup_out(a4_wr[800]), .rdlo_out(a4_wr[864]));
			radix2 #(.width(width)) rd_st3_801  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[801]), .rdlo_in(a3_wr[865]),  .coef_in(coef[264]), .rdup_out(a4_wr[801]), .rdlo_out(a4_wr[865]));
			radix2 #(.width(width)) rd_st3_802  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[802]), .rdlo_in(a3_wr[866]),  .coef_in(coef[272]), .rdup_out(a4_wr[802]), .rdlo_out(a4_wr[866]));
			radix2 #(.width(width)) rd_st3_803  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[803]), .rdlo_in(a3_wr[867]),  .coef_in(coef[280]), .rdup_out(a4_wr[803]), .rdlo_out(a4_wr[867]));
			radix2 #(.width(width)) rd_st3_804  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[804]), .rdlo_in(a3_wr[868]),  .coef_in(coef[288]), .rdup_out(a4_wr[804]), .rdlo_out(a4_wr[868]));
			radix2 #(.width(width)) rd_st3_805  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[805]), .rdlo_in(a3_wr[869]),  .coef_in(coef[296]), .rdup_out(a4_wr[805]), .rdlo_out(a4_wr[869]));
			radix2 #(.width(width)) rd_st3_806  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[806]), .rdlo_in(a3_wr[870]),  .coef_in(coef[304]), .rdup_out(a4_wr[806]), .rdlo_out(a4_wr[870]));
			radix2 #(.width(width)) rd_st3_807  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[807]), .rdlo_in(a3_wr[871]),  .coef_in(coef[312]), .rdup_out(a4_wr[807]), .rdlo_out(a4_wr[871]));
			radix2 #(.width(width)) rd_st3_808  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[808]), .rdlo_in(a3_wr[872]),  .coef_in(coef[320]), .rdup_out(a4_wr[808]), .rdlo_out(a4_wr[872]));
			radix2 #(.width(width)) rd_st3_809  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[809]), .rdlo_in(a3_wr[873]),  .coef_in(coef[328]), .rdup_out(a4_wr[809]), .rdlo_out(a4_wr[873]));
			radix2 #(.width(width)) rd_st3_810  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[810]), .rdlo_in(a3_wr[874]),  .coef_in(coef[336]), .rdup_out(a4_wr[810]), .rdlo_out(a4_wr[874]));
			radix2 #(.width(width)) rd_st3_811  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[811]), .rdlo_in(a3_wr[875]),  .coef_in(coef[344]), .rdup_out(a4_wr[811]), .rdlo_out(a4_wr[875]));
			radix2 #(.width(width)) rd_st3_812  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[812]), .rdlo_in(a3_wr[876]),  .coef_in(coef[352]), .rdup_out(a4_wr[812]), .rdlo_out(a4_wr[876]));
			radix2 #(.width(width)) rd_st3_813  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[813]), .rdlo_in(a3_wr[877]),  .coef_in(coef[360]), .rdup_out(a4_wr[813]), .rdlo_out(a4_wr[877]));
			radix2 #(.width(width)) rd_st3_814  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[814]), .rdlo_in(a3_wr[878]),  .coef_in(coef[368]), .rdup_out(a4_wr[814]), .rdlo_out(a4_wr[878]));
			radix2 #(.width(width)) rd_st3_815  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[815]), .rdlo_in(a3_wr[879]),  .coef_in(coef[376]), .rdup_out(a4_wr[815]), .rdlo_out(a4_wr[879]));
			radix2 #(.width(width)) rd_st3_816  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[816]), .rdlo_in(a3_wr[880]),  .coef_in(coef[384]), .rdup_out(a4_wr[816]), .rdlo_out(a4_wr[880]));
			radix2 #(.width(width)) rd_st3_817  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[817]), .rdlo_in(a3_wr[881]),  .coef_in(coef[392]), .rdup_out(a4_wr[817]), .rdlo_out(a4_wr[881]));
			radix2 #(.width(width)) rd_st3_818  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[818]), .rdlo_in(a3_wr[882]),  .coef_in(coef[400]), .rdup_out(a4_wr[818]), .rdlo_out(a4_wr[882]));
			radix2 #(.width(width)) rd_st3_819  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[819]), .rdlo_in(a3_wr[883]),  .coef_in(coef[408]), .rdup_out(a4_wr[819]), .rdlo_out(a4_wr[883]));
			radix2 #(.width(width)) rd_st3_820  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[820]), .rdlo_in(a3_wr[884]),  .coef_in(coef[416]), .rdup_out(a4_wr[820]), .rdlo_out(a4_wr[884]));
			radix2 #(.width(width)) rd_st3_821  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[821]), .rdlo_in(a3_wr[885]),  .coef_in(coef[424]), .rdup_out(a4_wr[821]), .rdlo_out(a4_wr[885]));
			radix2 #(.width(width)) rd_st3_822  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[822]), .rdlo_in(a3_wr[886]),  .coef_in(coef[432]), .rdup_out(a4_wr[822]), .rdlo_out(a4_wr[886]));
			radix2 #(.width(width)) rd_st3_823  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[823]), .rdlo_in(a3_wr[887]),  .coef_in(coef[440]), .rdup_out(a4_wr[823]), .rdlo_out(a4_wr[887]));
			radix2 #(.width(width)) rd_st3_824  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[824]), .rdlo_in(a3_wr[888]),  .coef_in(coef[448]), .rdup_out(a4_wr[824]), .rdlo_out(a4_wr[888]));
			radix2 #(.width(width)) rd_st3_825  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[825]), .rdlo_in(a3_wr[889]),  .coef_in(coef[456]), .rdup_out(a4_wr[825]), .rdlo_out(a4_wr[889]));
			radix2 #(.width(width)) rd_st3_826  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[826]), .rdlo_in(a3_wr[890]),  .coef_in(coef[464]), .rdup_out(a4_wr[826]), .rdlo_out(a4_wr[890]));
			radix2 #(.width(width)) rd_st3_827  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[827]), .rdlo_in(a3_wr[891]),  .coef_in(coef[472]), .rdup_out(a4_wr[827]), .rdlo_out(a4_wr[891]));
			radix2 #(.width(width)) rd_st3_828  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[828]), .rdlo_in(a3_wr[892]),  .coef_in(coef[480]), .rdup_out(a4_wr[828]), .rdlo_out(a4_wr[892]));
			radix2 #(.width(width)) rd_st3_829  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[829]), .rdlo_in(a3_wr[893]),  .coef_in(coef[488]), .rdup_out(a4_wr[829]), .rdlo_out(a4_wr[893]));
			radix2 #(.width(width)) rd_st3_830  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[830]), .rdlo_in(a3_wr[894]),  .coef_in(coef[496]), .rdup_out(a4_wr[830]), .rdlo_out(a4_wr[894]));
			radix2 #(.width(width)) rd_st3_831  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[831]), .rdlo_in(a3_wr[895]),  .coef_in(coef[504]), .rdup_out(a4_wr[831]), .rdlo_out(a4_wr[895]));
			radix2 #(.width(width)) rd_st3_896  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[896]), .rdlo_in(a3_wr[960]),  .coef_in(coef[0]), .rdup_out(a4_wr[896]), .rdlo_out(a4_wr[960]));
			radix2 #(.width(width)) rd_st3_897  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[897]), .rdlo_in(a3_wr[961]),  .coef_in(coef[8]), .rdup_out(a4_wr[897]), .rdlo_out(a4_wr[961]));
			radix2 #(.width(width)) rd_st3_898  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[898]), .rdlo_in(a3_wr[962]),  .coef_in(coef[16]), .rdup_out(a4_wr[898]), .rdlo_out(a4_wr[962]));
			radix2 #(.width(width)) rd_st3_899  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[899]), .rdlo_in(a3_wr[963]),  .coef_in(coef[24]), .rdup_out(a4_wr[899]), .rdlo_out(a4_wr[963]));
			radix2 #(.width(width)) rd_st3_900  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[900]), .rdlo_in(a3_wr[964]),  .coef_in(coef[32]), .rdup_out(a4_wr[900]), .rdlo_out(a4_wr[964]));
			radix2 #(.width(width)) rd_st3_901  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[901]), .rdlo_in(a3_wr[965]),  .coef_in(coef[40]), .rdup_out(a4_wr[901]), .rdlo_out(a4_wr[965]));
			radix2 #(.width(width)) rd_st3_902  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[902]), .rdlo_in(a3_wr[966]),  .coef_in(coef[48]), .rdup_out(a4_wr[902]), .rdlo_out(a4_wr[966]));
			radix2 #(.width(width)) rd_st3_903  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[903]), .rdlo_in(a3_wr[967]),  .coef_in(coef[56]), .rdup_out(a4_wr[903]), .rdlo_out(a4_wr[967]));
			radix2 #(.width(width)) rd_st3_904  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[904]), .rdlo_in(a3_wr[968]),  .coef_in(coef[64]), .rdup_out(a4_wr[904]), .rdlo_out(a4_wr[968]));
			radix2 #(.width(width)) rd_st3_905  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[905]), .rdlo_in(a3_wr[969]),  .coef_in(coef[72]), .rdup_out(a4_wr[905]), .rdlo_out(a4_wr[969]));
			radix2 #(.width(width)) rd_st3_906  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[906]), .rdlo_in(a3_wr[970]),  .coef_in(coef[80]), .rdup_out(a4_wr[906]), .rdlo_out(a4_wr[970]));
			radix2 #(.width(width)) rd_st3_907  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[907]), .rdlo_in(a3_wr[971]),  .coef_in(coef[88]), .rdup_out(a4_wr[907]), .rdlo_out(a4_wr[971]));
			radix2 #(.width(width)) rd_st3_908  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[908]), .rdlo_in(a3_wr[972]),  .coef_in(coef[96]), .rdup_out(a4_wr[908]), .rdlo_out(a4_wr[972]));
			radix2 #(.width(width)) rd_st3_909  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[909]), .rdlo_in(a3_wr[973]),  .coef_in(coef[104]), .rdup_out(a4_wr[909]), .rdlo_out(a4_wr[973]));
			radix2 #(.width(width)) rd_st3_910  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[910]), .rdlo_in(a3_wr[974]),  .coef_in(coef[112]), .rdup_out(a4_wr[910]), .rdlo_out(a4_wr[974]));
			radix2 #(.width(width)) rd_st3_911  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[911]), .rdlo_in(a3_wr[975]),  .coef_in(coef[120]), .rdup_out(a4_wr[911]), .rdlo_out(a4_wr[975]));
			radix2 #(.width(width)) rd_st3_912  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[912]), .rdlo_in(a3_wr[976]),  .coef_in(coef[128]), .rdup_out(a4_wr[912]), .rdlo_out(a4_wr[976]));
			radix2 #(.width(width)) rd_st3_913  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[913]), .rdlo_in(a3_wr[977]),  .coef_in(coef[136]), .rdup_out(a4_wr[913]), .rdlo_out(a4_wr[977]));
			radix2 #(.width(width)) rd_st3_914  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[914]), .rdlo_in(a3_wr[978]),  .coef_in(coef[144]), .rdup_out(a4_wr[914]), .rdlo_out(a4_wr[978]));
			radix2 #(.width(width)) rd_st3_915  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[915]), .rdlo_in(a3_wr[979]),  .coef_in(coef[152]), .rdup_out(a4_wr[915]), .rdlo_out(a4_wr[979]));
			radix2 #(.width(width)) rd_st3_916  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[916]), .rdlo_in(a3_wr[980]),  .coef_in(coef[160]), .rdup_out(a4_wr[916]), .rdlo_out(a4_wr[980]));
			radix2 #(.width(width)) rd_st3_917  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[917]), .rdlo_in(a3_wr[981]),  .coef_in(coef[168]), .rdup_out(a4_wr[917]), .rdlo_out(a4_wr[981]));
			radix2 #(.width(width)) rd_st3_918  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[918]), .rdlo_in(a3_wr[982]),  .coef_in(coef[176]), .rdup_out(a4_wr[918]), .rdlo_out(a4_wr[982]));
			radix2 #(.width(width)) rd_st3_919  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[919]), .rdlo_in(a3_wr[983]),  .coef_in(coef[184]), .rdup_out(a4_wr[919]), .rdlo_out(a4_wr[983]));
			radix2 #(.width(width)) rd_st3_920  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[920]), .rdlo_in(a3_wr[984]),  .coef_in(coef[192]), .rdup_out(a4_wr[920]), .rdlo_out(a4_wr[984]));
			radix2 #(.width(width)) rd_st3_921  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[921]), .rdlo_in(a3_wr[985]),  .coef_in(coef[200]), .rdup_out(a4_wr[921]), .rdlo_out(a4_wr[985]));
			radix2 #(.width(width)) rd_st3_922  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[922]), .rdlo_in(a3_wr[986]),  .coef_in(coef[208]), .rdup_out(a4_wr[922]), .rdlo_out(a4_wr[986]));
			radix2 #(.width(width)) rd_st3_923  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[923]), .rdlo_in(a3_wr[987]),  .coef_in(coef[216]), .rdup_out(a4_wr[923]), .rdlo_out(a4_wr[987]));
			radix2 #(.width(width)) rd_st3_924  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[924]), .rdlo_in(a3_wr[988]),  .coef_in(coef[224]), .rdup_out(a4_wr[924]), .rdlo_out(a4_wr[988]));
			radix2 #(.width(width)) rd_st3_925  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[925]), .rdlo_in(a3_wr[989]),  .coef_in(coef[232]), .rdup_out(a4_wr[925]), .rdlo_out(a4_wr[989]));
			radix2 #(.width(width)) rd_st3_926  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[926]), .rdlo_in(a3_wr[990]),  .coef_in(coef[240]), .rdup_out(a4_wr[926]), .rdlo_out(a4_wr[990]));
			radix2 #(.width(width)) rd_st3_927  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[927]), .rdlo_in(a3_wr[991]),  .coef_in(coef[248]), .rdup_out(a4_wr[927]), .rdlo_out(a4_wr[991]));
			radix2 #(.width(width)) rd_st3_928  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[928]), .rdlo_in(a3_wr[992]),  .coef_in(coef[256]), .rdup_out(a4_wr[928]), .rdlo_out(a4_wr[992]));
			radix2 #(.width(width)) rd_st3_929  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[929]), .rdlo_in(a3_wr[993]),  .coef_in(coef[264]), .rdup_out(a4_wr[929]), .rdlo_out(a4_wr[993]));
			radix2 #(.width(width)) rd_st3_930  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[930]), .rdlo_in(a3_wr[994]),  .coef_in(coef[272]), .rdup_out(a4_wr[930]), .rdlo_out(a4_wr[994]));
			radix2 #(.width(width)) rd_st3_931  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[931]), .rdlo_in(a3_wr[995]),  .coef_in(coef[280]), .rdup_out(a4_wr[931]), .rdlo_out(a4_wr[995]));
			radix2 #(.width(width)) rd_st3_932  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[932]), .rdlo_in(a3_wr[996]),  .coef_in(coef[288]), .rdup_out(a4_wr[932]), .rdlo_out(a4_wr[996]));
			radix2 #(.width(width)) rd_st3_933  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[933]), .rdlo_in(a3_wr[997]),  .coef_in(coef[296]), .rdup_out(a4_wr[933]), .rdlo_out(a4_wr[997]));
			radix2 #(.width(width)) rd_st3_934  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[934]), .rdlo_in(a3_wr[998]),  .coef_in(coef[304]), .rdup_out(a4_wr[934]), .rdlo_out(a4_wr[998]));
			radix2 #(.width(width)) rd_st3_935  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[935]), .rdlo_in(a3_wr[999]),  .coef_in(coef[312]), .rdup_out(a4_wr[935]), .rdlo_out(a4_wr[999]));
			radix2 #(.width(width)) rd_st3_936  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[936]), .rdlo_in(a3_wr[1000]),  .coef_in(coef[320]), .rdup_out(a4_wr[936]), .rdlo_out(a4_wr[1000]));
			radix2 #(.width(width)) rd_st3_937  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[937]), .rdlo_in(a3_wr[1001]),  .coef_in(coef[328]), .rdup_out(a4_wr[937]), .rdlo_out(a4_wr[1001]));
			radix2 #(.width(width)) rd_st3_938  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[938]), .rdlo_in(a3_wr[1002]),  .coef_in(coef[336]), .rdup_out(a4_wr[938]), .rdlo_out(a4_wr[1002]));
			radix2 #(.width(width)) rd_st3_939  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[939]), .rdlo_in(a3_wr[1003]),  .coef_in(coef[344]), .rdup_out(a4_wr[939]), .rdlo_out(a4_wr[1003]));
			radix2 #(.width(width)) rd_st3_940  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[940]), .rdlo_in(a3_wr[1004]),  .coef_in(coef[352]), .rdup_out(a4_wr[940]), .rdlo_out(a4_wr[1004]));
			radix2 #(.width(width)) rd_st3_941  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[941]), .rdlo_in(a3_wr[1005]),  .coef_in(coef[360]), .rdup_out(a4_wr[941]), .rdlo_out(a4_wr[1005]));
			radix2 #(.width(width)) rd_st3_942  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[942]), .rdlo_in(a3_wr[1006]),  .coef_in(coef[368]), .rdup_out(a4_wr[942]), .rdlo_out(a4_wr[1006]));
			radix2 #(.width(width)) rd_st3_943  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[943]), .rdlo_in(a3_wr[1007]),  .coef_in(coef[376]), .rdup_out(a4_wr[943]), .rdlo_out(a4_wr[1007]));
			radix2 #(.width(width)) rd_st3_944  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[944]), .rdlo_in(a3_wr[1008]),  .coef_in(coef[384]), .rdup_out(a4_wr[944]), .rdlo_out(a4_wr[1008]));
			radix2 #(.width(width)) rd_st3_945  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[945]), .rdlo_in(a3_wr[1009]),  .coef_in(coef[392]), .rdup_out(a4_wr[945]), .rdlo_out(a4_wr[1009]));
			radix2 #(.width(width)) rd_st3_946  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[946]), .rdlo_in(a3_wr[1010]),  .coef_in(coef[400]), .rdup_out(a4_wr[946]), .rdlo_out(a4_wr[1010]));
			radix2 #(.width(width)) rd_st3_947  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[947]), .rdlo_in(a3_wr[1011]),  .coef_in(coef[408]), .rdup_out(a4_wr[947]), .rdlo_out(a4_wr[1011]));
			radix2 #(.width(width)) rd_st3_948  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[948]), .rdlo_in(a3_wr[1012]),  .coef_in(coef[416]), .rdup_out(a4_wr[948]), .rdlo_out(a4_wr[1012]));
			radix2 #(.width(width)) rd_st3_949  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[949]), .rdlo_in(a3_wr[1013]),  .coef_in(coef[424]), .rdup_out(a4_wr[949]), .rdlo_out(a4_wr[1013]));
			radix2 #(.width(width)) rd_st3_950  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[950]), .rdlo_in(a3_wr[1014]),  .coef_in(coef[432]), .rdup_out(a4_wr[950]), .rdlo_out(a4_wr[1014]));
			radix2 #(.width(width)) rd_st3_951  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[951]), .rdlo_in(a3_wr[1015]),  .coef_in(coef[440]), .rdup_out(a4_wr[951]), .rdlo_out(a4_wr[1015]));
			radix2 #(.width(width)) rd_st3_952  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[952]), .rdlo_in(a3_wr[1016]),  .coef_in(coef[448]), .rdup_out(a4_wr[952]), .rdlo_out(a4_wr[1016]));
			radix2 #(.width(width)) rd_st3_953  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[953]), .rdlo_in(a3_wr[1017]),  .coef_in(coef[456]), .rdup_out(a4_wr[953]), .rdlo_out(a4_wr[1017]));
			radix2 #(.width(width)) rd_st3_954  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[954]), .rdlo_in(a3_wr[1018]),  .coef_in(coef[464]), .rdup_out(a4_wr[954]), .rdlo_out(a4_wr[1018]));
			radix2 #(.width(width)) rd_st3_955  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[955]), .rdlo_in(a3_wr[1019]),  .coef_in(coef[472]), .rdup_out(a4_wr[955]), .rdlo_out(a4_wr[1019]));
			radix2 #(.width(width)) rd_st3_956  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[956]), .rdlo_in(a3_wr[1020]),  .coef_in(coef[480]), .rdup_out(a4_wr[956]), .rdlo_out(a4_wr[1020]));
			radix2 #(.width(width)) rd_st3_957  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[957]), .rdlo_in(a3_wr[1021]),  .coef_in(coef[488]), .rdup_out(a4_wr[957]), .rdlo_out(a4_wr[1021]));
			radix2 #(.width(width)) rd_st3_958  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[958]), .rdlo_in(a3_wr[1022]),  .coef_in(coef[496]), .rdup_out(a4_wr[958]), .rdlo_out(a4_wr[1022]));
			radix2 #(.width(width)) rd_st3_959  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[959]), .rdlo_in(a3_wr[1023]),  .coef_in(coef[504]), .rdup_out(a4_wr[959]), .rdlo_out(a4_wr[1023]));

		//--- radix stage 4
			radix2 #(.width(width)) rd_st4_0   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[0]), .rdlo_in(a4_wr[32]),  .coef_in(coef[0]), .rdup_out(a5_wr[0]), .rdlo_out(a5_wr[32]));
			radix2 #(.width(width)) rd_st4_1   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1]), .rdlo_in(a4_wr[33]),  .coef_in(coef[16]), .rdup_out(a5_wr[1]), .rdlo_out(a5_wr[33]));
			radix2 #(.width(width)) rd_st4_2   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[2]), .rdlo_in(a4_wr[34]),  .coef_in(coef[32]), .rdup_out(a5_wr[2]), .rdlo_out(a5_wr[34]));
			radix2 #(.width(width)) rd_st4_3   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[3]), .rdlo_in(a4_wr[35]),  .coef_in(coef[48]), .rdup_out(a5_wr[3]), .rdlo_out(a5_wr[35]));
			radix2 #(.width(width)) rd_st4_4   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[4]), .rdlo_in(a4_wr[36]),  .coef_in(coef[64]), .rdup_out(a5_wr[4]), .rdlo_out(a5_wr[36]));
			radix2 #(.width(width)) rd_st4_5   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[5]), .rdlo_in(a4_wr[37]),  .coef_in(coef[80]), .rdup_out(a5_wr[5]), .rdlo_out(a5_wr[37]));
			radix2 #(.width(width)) rd_st4_6   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[6]), .rdlo_in(a4_wr[38]),  .coef_in(coef[96]), .rdup_out(a5_wr[6]), .rdlo_out(a5_wr[38]));
			radix2 #(.width(width)) rd_st4_7   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[7]), .rdlo_in(a4_wr[39]),  .coef_in(coef[112]), .rdup_out(a5_wr[7]), .rdlo_out(a5_wr[39]));
			radix2 #(.width(width)) rd_st4_8   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[8]), .rdlo_in(a4_wr[40]),  .coef_in(coef[128]), .rdup_out(a5_wr[8]), .rdlo_out(a5_wr[40]));
			radix2 #(.width(width)) rd_st4_9   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[9]), .rdlo_in(a4_wr[41]),  .coef_in(coef[144]), .rdup_out(a5_wr[9]), .rdlo_out(a5_wr[41]));
			radix2 #(.width(width)) rd_st4_10  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[10]), .rdlo_in(a4_wr[42]),  .coef_in(coef[160]), .rdup_out(a5_wr[10]), .rdlo_out(a5_wr[42]));
			radix2 #(.width(width)) rd_st4_11  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[11]), .rdlo_in(a4_wr[43]),  .coef_in(coef[176]), .rdup_out(a5_wr[11]), .rdlo_out(a5_wr[43]));
			radix2 #(.width(width)) rd_st4_12  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[12]), .rdlo_in(a4_wr[44]),  .coef_in(coef[192]), .rdup_out(a5_wr[12]), .rdlo_out(a5_wr[44]));
			radix2 #(.width(width)) rd_st4_13  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[13]), .rdlo_in(a4_wr[45]),  .coef_in(coef[208]), .rdup_out(a5_wr[13]), .rdlo_out(a5_wr[45]));
			radix2 #(.width(width)) rd_st4_14  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[14]), .rdlo_in(a4_wr[46]),  .coef_in(coef[224]), .rdup_out(a5_wr[14]), .rdlo_out(a5_wr[46]));
			radix2 #(.width(width)) rd_st4_15  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[15]), .rdlo_in(a4_wr[47]),  .coef_in(coef[240]), .rdup_out(a5_wr[15]), .rdlo_out(a5_wr[47]));
			radix2 #(.width(width)) rd_st4_16  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[16]), .rdlo_in(a4_wr[48]),  .coef_in(coef[256]), .rdup_out(a5_wr[16]), .rdlo_out(a5_wr[48]));
			radix2 #(.width(width)) rd_st4_17  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[17]), .rdlo_in(a4_wr[49]),  .coef_in(coef[272]), .rdup_out(a5_wr[17]), .rdlo_out(a5_wr[49]));
			radix2 #(.width(width)) rd_st4_18  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[18]), .rdlo_in(a4_wr[50]),  .coef_in(coef[288]), .rdup_out(a5_wr[18]), .rdlo_out(a5_wr[50]));
			radix2 #(.width(width)) rd_st4_19  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[19]), .rdlo_in(a4_wr[51]),  .coef_in(coef[304]), .rdup_out(a5_wr[19]), .rdlo_out(a5_wr[51]));
			radix2 #(.width(width)) rd_st4_20  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[20]), .rdlo_in(a4_wr[52]),  .coef_in(coef[320]), .rdup_out(a5_wr[20]), .rdlo_out(a5_wr[52]));
			radix2 #(.width(width)) rd_st4_21  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[21]), .rdlo_in(a4_wr[53]),  .coef_in(coef[336]), .rdup_out(a5_wr[21]), .rdlo_out(a5_wr[53]));
			radix2 #(.width(width)) rd_st4_22  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[22]), .rdlo_in(a4_wr[54]),  .coef_in(coef[352]), .rdup_out(a5_wr[22]), .rdlo_out(a5_wr[54]));
			radix2 #(.width(width)) rd_st4_23  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[23]), .rdlo_in(a4_wr[55]),  .coef_in(coef[368]), .rdup_out(a5_wr[23]), .rdlo_out(a5_wr[55]));
			radix2 #(.width(width)) rd_st4_24  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[24]), .rdlo_in(a4_wr[56]),  .coef_in(coef[384]), .rdup_out(a5_wr[24]), .rdlo_out(a5_wr[56]));
			radix2 #(.width(width)) rd_st4_25  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[25]), .rdlo_in(a4_wr[57]),  .coef_in(coef[400]), .rdup_out(a5_wr[25]), .rdlo_out(a5_wr[57]));
			radix2 #(.width(width)) rd_st4_26  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[26]), .rdlo_in(a4_wr[58]),  .coef_in(coef[416]), .rdup_out(a5_wr[26]), .rdlo_out(a5_wr[58]));
			radix2 #(.width(width)) rd_st4_27  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[27]), .rdlo_in(a4_wr[59]),  .coef_in(coef[432]), .rdup_out(a5_wr[27]), .rdlo_out(a5_wr[59]));
			radix2 #(.width(width)) rd_st4_28  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[28]), .rdlo_in(a4_wr[60]),  .coef_in(coef[448]), .rdup_out(a5_wr[28]), .rdlo_out(a5_wr[60]));
			radix2 #(.width(width)) rd_st4_29  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[29]), .rdlo_in(a4_wr[61]),  .coef_in(coef[464]), .rdup_out(a5_wr[29]), .rdlo_out(a5_wr[61]));
			radix2 #(.width(width)) rd_st4_30  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[30]), .rdlo_in(a4_wr[62]),  .coef_in(coef[480]), .rdup_out(a5_wr[30]), .rdlo_out(a5_wr[62]));
			radix2 #(.width(width)) rd_st4_31  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[31]), .rdlo_in(a4_wr[63]),  .coef_in(coef[496]), .rdup_out(a5_wr[31]), .rdlo_out(a5_wr[63]));
			radix2 #(.width(width)) rd_st4_64  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[64]), .rdlo_in(a4_wr[96]),  .coef_in(coef[0]), .rdup_out(a5_wr[64]), .rdlo_out(a5_wr[96]));
			radix2 #(.width(width)) rd_st4_65  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[65]), .rdlo_in(a4_wr[97]),  .coef_in(coef[16]), .rdup_out(a5_wr[65]), .rdlo_out(a5_wr[97]));
			radix2 #(.width(width)) rd_st4_66  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[66]), .rdlo_in(a4_wr[98]),  .coef_in(coef[32]), .rdup_out(a5_wr[66]), .rdlo_out(a5_wr[98]));
			radix2 #(.width(width)) rd_st4_67  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[67]), .rdlo_in(a4_wr[99]),  .coef_in(coef[48]), .rdup_out(a5_wr[67]), .rdlo_out(a5_wr[99]));
			radix2 #(.width(width)) rd_st4_68  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[68]), .rdlo_in(a4_wr[100]),  .coef_in(coef[64]), .rdup_out(a5_wr[68]), .rdlo_out(a5_wr[100]));
			radix2 #(.width(width)) rd_st4_69  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[69]), .rdlo_in(a4_wr[101]),  .coef_in(coef[80]), .rdup_out(a5_wr[69]), .rdlo_out(a5_wr[101]));
			radix2 #(.width(width)) rd_st4_70  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[70]), .rdlo_in(a4_wr[102]),  .coef_in(coef[96]), .rdup_out(a5_wr[70]), .rdlo_out(a5_wr[102]));
			radix2 #(.width(width)) rd_st4_71  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[71]), .rdlo_in(a4_wr[103]),  .coef_in(coef[112]), .rdup_out(a5_wr[71]), .rdlo_out(a5_wr[103]));
			radix2 #(.width(width)) rd_st4_72  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[72]), .rdlo_in(a4_wr[104]),  .coef_in(coef[128]), .rdup_out(a5_wr[72]), .rdlo_out(a5_wr[104]));
			radix2 #(.width(width)) rd_st4_73  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[73]), .rdlo_in(a4_wr[105]),  .coef_in(coef[144]), .rdup_out(a5_wr[73]), .rdlo_out(a5_wr[105]));
			radix2 #(.width(width)) rd_st4_74  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[74]), .rdlo_in(a4_wr[106]),  .coef_in(coef[160]), .rdup_out(a5_wr[74]), .rdlo_out(a5_wr[106]));
			radix2 #(.width(width)) rd_st4_75  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[75]), .rdlo_in(a4_wr[107]),  .coef_in(coef[176]), .rdup_out(a5_wr[75]), .rdlo_out(a5_wr[107]));
			radix2 #(.width(width)) rd_st4_76  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[76]), .rdlo_in(a4_wr[108]),  .coef_in(coef[192]), .rdup_out(a5_wr[76]), .rdlo_out(a5_wr[108]));
			radix2 #(.width(width)) rd_st4_77  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[77]), .rdlo_in(a4_wr[109]),  .coef_in(coef[208]), .rdup_out(a5_wr[77]), .rdlo_out(a5_wr[109]));
			radix2 #(.width(width)) rd_st4_78  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[78]), .rdlo_in(a4_wr[110]),  .coef_in(coef[224]), .rdup_out(a5_wr[78]), .rdlo_out(a5_wr[110]));
			radix2 #(.width(width)) rd_st4_79  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[79]), .rdlo_in(a4_wr[111]),  .coef_in(coef[240]), .rdup_out(a5_wr[79]), .rdlo_out(a5_wr[111]));
			radix2 #(.width(width)) rd_st4_80  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[80]), .rdlo_in(a4_wr[112]),  .coef_in(coef[256]), .rdup_out(a5_wr[80]), .rdlo_out(a5_wr[112]));
			radix2 #(.width(width)) rd_st4_81  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[81]), .rdlo_in(a4_wr[113]),  .coef_in(coef[272]), .rdup_out(a5_wr[81]), .rdlo_out(a5_wr[113]));
			radix2 #(.width(width)) rd_st4_82  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[82]), .rdlo_in(a4_wr[114]),  .coef_in(coef[288]), .rdup_out(a5_wr[82]), .rdlo_out(a5_wr[114]));
			radix2 #(.width(width)) rd_st4_83  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[83]), .rdlo_in(a4_wr[115]),  .coef_in(coef[304]), .rdup_out(a5_wr[83]), .rdlo_out(a5_wr[115]));
			radix2 #(.width(width)) rd_st4_84  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[84]), .rdlo_in(a4_wr[116]),  .coef_in(coef[320]), .rdup_out(a5_wr[84]), .rdlo_out(a5_wr[116]));
			radix2 #(.width(width)) rd_st4_85  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[85]), .rdlo_in(a4_wr[117]),  .coef_in(coef[336]), .rdup_out(a5_wr[85]), .rdlo_out(a5_wr[117]));
			radix2 #(.width(width)) rd_st4_86  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[86]), .rdlo_in(a4_wr[118]),  .coef_in(coef[352]), .rdup_out(a5_wr[86]), .rdlo_out(a5_wr[118]));
			radix2 #(.width(width)) rd_st4_87  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[87]), .rdlo_in(a4_wr[119]),  .coef_in(coef[368]), .rdup_out(a5_wr[87]), .rdlo_out(a5_wr[119]));
			radix2 #(.width(width)) rd_st4_88  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[88]), .rdlo_in(a4_wr[120]),  .coef_in(coef[384]), .rdup_out(a5_wr[88]), .rdlo_out(a5_wr[120]));
			radix2 #(.width(width)) rd_st4_89  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[89]), .rdlo_in(a4_wr[121]),  .coef_in(coef[400]), .rdup_out(a5_wr[89]), .rdlo_out(a5_wr[121]));
			radix2 #(.width(width)) rd_st4_90  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[90]), .rdlo_in(a4_wr[122]),  .coef_in(coef[416]), .rdup_out(a5_wr[90]), .rdlo_out(a5_wr[122]));
			radix2 #(.width(width)) rd_st4_91  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[91]), .rdlo_in(a4_wr[123]),  .coef_in(coef[432]), .rdup_out(a5_wr[91]), .rdlo_out(a5_wr[123]));
			radix2 #(.width(width)) rd_st4_92  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[92]), .rdlo_in(a4_wr[124]),  .coef_in(coef[448]), .rdup_out(a5_wr[92]), .rdlo_out(a5_wr[124]));
			radix2 #(.width(width)) rd_st4_93  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[93]), .rdlo_in(a4_wr[125]),  .coef_in(coef[464]), .rdup_out(a5_wr[93]), .rdlo_out(a5_wr[125]));
			radix2 #(.width(width)) rd_st4_94  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[94]), .rdlo_in(a4_wr[126]),  .coef_in(coef[480]), .rdup_out(a5_wr[94]), .rdlo_out(a5_wr[126]));
			radix2 #(.width(width)) rd_st4_95  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[95]), .rdlo_in(a4_wr[127]),  .coef_in(coef[496]), .rdup_out(a5_wr[95]), .rdlo_out(a5_wr[127]));
			radix2 #(.width(width)) rd_st4_128  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[128]), .rdlo_in(a4_wr[160]),  .coef_in(coef[0]), .rdup_out(a5_wr[128]), .rdlo_out(a5_wr[160]));
			radix2 #(.width(width)) rd_st4_129  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[129]), .rdlo_in(a4_wr[161]),  .coef_in(coef[16]), .rdup_out(a5_wr[129]), .rdlo_out(a5_wr[161]));
			radix2 #(.width(width)) rd_st4_130  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[130]), .rdlo_in(a4_wr[162]),  .coef_in(coef[32]), .rdup_out(a5_wr[130]), .rdlo_out(a5_wr[162]));
			radix2 #(.width(width)) rd_st4_131  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[131]), .rdlo_in(a4_wr[163]),  .coef_in(coef[48]), .rdup_out(a5_wr[131]), .rdlo_out(a5_wr[163]));
			radix2 #(.width(width)) rd_st4_132  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[132]), .rdlo_in(a4_wr[164]),  .coef_in(coef[64]), .rdup_out(a5_wr[132]), .rdlo_out(a5_wr[164]));
			radix2 #(.width(width)) rd_st4_133  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[133]), .rdlo_in(a4_wr[165]),  .coef_in(coef[80]), .rdup_out(a5_wr[133]), .rdlo_out(a5_wr[165]));
			radix2 #(.width(width)) rd_st4_134  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[134]), .rdlo_in(a4_wr[166]),  .coef_in(coef[96]), .rdup_out(a5_wr[134]), .rdlo_out(a5_wr[166]));
			radix2 #(.width(width)) rd_st4_135  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[135]), .rdlo_in(a4_wr[167]),  .coef_in(coef[112]), .rdup_out(a5_wr[135]), .rdlo_out(a5_wr[167]));
			radix2 #(.width(width)) rd_st4_136  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[136]), .rdlo_in(a4_wr[168]),  .coef_in(coef[128]), .rdup_out(a5_wr[136]), .rdlo_out(a5_wr[168]));
			radix2 #(.width(width)) rd_st4_137  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[137]), .rdlo_in(a4_wr[169]),  .coef_in(coef[144]), .rdup_out(a5_wr[137]), .rdlo_out(a5_wr[169]));
			radix2 #(.width(width)) rd_st4_138  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[138]), .rdlo_in(a4_wr[170]),  .coef_in(coef[160]), .rdup_out(a5_wr[138]), .rdlo_out(a5_wr[170]));
			radix2 #(.width(width)) rd_st4_139  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[139]), .rdlo_in(a4_wr[171]),  .coef_in(coef[176]), .rdup_out(a5_wr[139]), .rdlo_out(a5_wr[171]));
			radix2 #(.width(width)) rd_st4_140  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[140]), .rdlo_in(a4_wr[172]),  .coef_in(coef[192]), .rdup_out(a5_wr[140]), .rdlo_out(a5_wr[172]));
			radix2 #(.width(width)) rd_st4_141  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[141]), .rdlo_in(a4_wr[173]),  .coef_in(coef[208]), .rdup_out(a5_wr[141]), .rdlo_out(a5_wr[173]));
			radix2 #(.width(width)) rd_st4_142  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[142]), .rdlo_in(a4_wr[174]),  .coef_in(coef[224]), .rdup_out(a5_wr[142]), .rdlo_out(a5_wr[174]));
			radix2 #(.width(width)) rd_st4_143  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[143]), .rdlo_in(a4_wr[175]),  .coef_in(coef[240]), .rdup_out(a5_wr[143]), .rdlo_out(a5_wr[175]));
			radix2 #(.width(width)) rd_st4_144  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[144]), .rdlo_in(a4_wr[176]),  .coef_in(coef[256]), .rdup_out(a5_wr[144]), .rdlo_out(a5_wr[176]));
			radix2 #(.width(width)) rd_st4_145  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[145]), .rdlo_in(a4_wr[177]),  .coef_in(coef[272]), .rdup_out(a5_wr[145]), .rdlo_out(a5_wr[177]));
			radix2 #(.width(width)) rd_st4_146  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[146]), .rdlo_in(a4_wr[178]),  .coef_in(coef[288]), .rdup_out(a5_wr[146]), .rdlo_out(a5_wr[178]));
			radix2 #(.width(width)) rd_st4_147  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[147]), .rdlo_in(a4_wr[179]),  .coef_in(coef[304]), .rdup_out(a5_wr[147]), .rdlo_out(a5_wr[179]));
			radix2 #(.width(width)) rd_st4_148  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[148]), .rdlo_in(a4_wr[180]),  .coef_in(coef[320]), .rdup_out(a5_wr[148]), .rdlo_out(a5_wr[180]));
			radix2 #(.width(width)) rd_st4_149  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[149]), .rdlo_in(a4_wr[181]),  .coef_in(coef[336]), .rdup_out(a5_wr[149]), .rdlo_out(a5_wr[181]));
			radix2 #(.width(width)) rd_st4_150  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[150]), .rdlo_in(a4_wr[182]),  .coef_in(coef[352]), .rdup_out(a5_wr[150]), .rdlo_out(a5_wr[182]));
			radix2 #(.width(width)) rd_st4_151  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[151]), .rdlo_in(a4_wr[183]),  .coef_in(coef[368]), .rdup_out(a5_wr[151]), .rdlo_out(a5_wr[183]));
			radix2 #(.width(width)) rd_st4_152  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[152]), .rdlo_in(a4_wr[184]),  .coef_in(coef[384]), .rdup_out(a5_wr[152]), .rdlo_out(a5_wr[184]));
			radix2 #(.width(width)) rd_st4_153  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[153]), .rdlo_in(a4_wr[185]),  .coef_in(coef[400]), .rdup_out(a5_wr[153]), .rdlo_out(a5_wr[185]));
			radix2 #(.width(width)) rd_st4_154  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[154]), .rdlo_in(a4_wr[186]),  .coef_in(coef[416]), .rdup_out(a5_wr[154]), .rdlo_out(a5_wr[186]));
			radix2 #(.width(width)) rd_st4_155  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[155]), .rdlo_in(a4_wr[187]),  .coef_in(coef[432]), .rdup_out(a5_wr[155]), .rdlo_out(a5_wr[187]));
			radix2 #(.width(width)) rd_st4_156  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[156]), .rdlo_in(a4_wr[188]),  .coef_in(coef[448]), .rdup_out(a5_wr[156]), .rdlo_out(a5_wr[188]));
			radix2 #(.width(width)) rd_st4_157  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[157]), .rdlo_in(a4_wr[189]),  .coef_in(coef[464]), .rdup_out(a5_wr[157]), .rdlo_out(a5_wr[189]));
			radix2 #(.width(width)) rd_st4_158  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[158]), .rdlo_in(a4_wr[190]),  .coef_in(coef[480]), .rdup_out(a5_wr[158]), .rdlo_out(a5_wr[190]));
			radix2 #(.width(width)) rd_st4_159  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[159]), .rdlo_in(a4_wr[191]),  .coef_in(coef[496]), .rdup_out(a5_wr[159]), .rdlo_out(a5_wr[191]));
			radix2 #(.width(width)) rd_st4_192  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[192]), .rdlo_in(a4_wr[224]),  .coef_in(coef[0]), .rdup_out(a5_wr[192]), .rdlo_out(a5_wr[224]));
			radix2 #(.width(width)) rd_st4_193  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[193]), .rdlo_in(a4_wr[225]),  .coef_in(coef[16]), .rdup_out(a5_wr[193]), .rdlo_out(a5_wr[225]));
			radix2 #(.width(width)) rd_st4_194  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[194]), .rdlo_in(a4_wr[226]),  .coef_in(coef[32]), .rdup_out(a5_wr[194]), .rdlo_out(a5_wr[226]));
			radix2 #(.width(width)) rd_st4_195  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[195]), .rdlo_in(a4_wr[227]),  .coef_in(coef[48]), .rdup_out(a5_wr[195]), .rdlo_out(a5_wr[227]));
			radix2 #(.width(width)) rd_st4_196  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[196]), .rdlo_in(a4_wr[228]),  .coef_in(coef[64]), .rdup_out(a5_wr[196]), .rdlo_out(a5_wr[228]));
			radix2 #(.width(width)) rd_st4_197  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[197]), .rdlo_in(a4_wr[229]),  .coef_in(coef[80]), .rdup_out(a5_wr[197]), .rdlo_out(a5_wr[229]));
			radix2 #(.width(width)) rd_st4_198  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[198]), .rdlo_in(a4_wr[230]),  .coef_in(coef[96]), .rdup_out(a5_wr[198]), .rdlo_out(a5_wr[230]));
			radix2 #(.width(width)) rd_st4_199  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[199]), .rdlo_in(a4_wr[231]),  .coef_in(coef[112]), .rdup_out(a5_wr[199]), .rdlo_out(a5_wr[231]));
			radix2 #(.width(width)) rd_st4_200  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[200]), .rdlo_in(a4_wr[232]),  .coef_in(coef[128]), .rdup_out(a5_wr[200]), .rdlo_out(a5_wr[232]));
			radix2 #(.width(width)) rd_st4_201  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[201]), .rdlo_in(a4_wr[233]),  .coef_in(coef[144]), .rdup_out(a5_wr[201]), .rdlo_out(a5_wr[233]));
			radix2 #(.width(width)) rd_st4_202  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[202]), .rdlo_in(a4_wr[234]),  .coef_in(coef[160]), .rdup_out(a5_wr[202]), .rdlo_out(a5_wr[234]));
			radix2 #(.width(width)) rd_st4_203  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[203]), .rdlo_in(a4_wr[235]),  .coef_in(coef[176]), .rdup_out(a5_wr[203]), .rdlo_out(a5_wr[235]));
			radix2 #(.width(width)) rd_st4_204  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[204]), .rdlo_in(a4_wr[236]),  .coef_in(coef[192]), .rdup_out(a5_wr[204]), .rdlo_out(a5_wr[236]));
			radix2 #(.width(width)) rd_st4_205  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[205]), .rdlo_in(a4_wr[237]),  .coef_in(coef[208]), .rdup_out(a5_wr[205]), .rdlo_out(a5_wr[237]));
			radix2 #(.width(width)) rd_st4_206  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[206]), .rdlo_in(a4_wr[238]),  .coef_in(coef[224]), .rdup_out(a5_wr[206]), .rdlo_out(a5_wr[238]));
			radix2 #(.width(width)) rd_st4_207  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[207]), .rdlo_in(a4_wr[239]),  .coef_in(coef[240]), .rdup_out(a5_wr[207]), .rdlo_out(a5_wr[239]));
			radix2 #(.width(width)) rd_st4_208  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[208]), .rdlo_in(a4_wr[240]),  .coef_in(coef[256]), .rdup_out(a5_wr[208]), .rdlo_out(a5_wr[240]));
			radix2 #(.width(width)) rd_st4_209  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[209]), .rdlo_in(a4_wr[241]),  .coef_in(coef[272]), .rdup_out(a5_wr[209]), .rdlo_out(a5_wr[241]));
			radix2 #(.width(width)) rd_st4_210  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[210]), .rdlo_in(a4_wr[242]),  .coef_in(coef[288]), .rdup_out(a5_wr[210]), .rdlo_out(a5_wr[242]));
			radix2 #(.width(width)) rd_st4_211  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[211]), .rdlo_in(a4_wr[243]),  .coef_in(coef[304]), .rdup_out(a5_wr[211]), .rdlo_out(a5_wr[243]));
			radix2 #(.width(width)) rd_st4_212  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[212]), .rdlo_in(a4_wr[244]),  .coef_in(coef[320]), .rdup_out(a5_wr[212]), .rdlo_out(a5_wr[244]));
			radix2 #(.width(width)) rd_st4_213  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[213]), .rdlo_in(a4_wr[245]),  .coef_in(coef[336]), .rdup_out(a5_wr[213]), .rdlo_out(a5_wr[245]));
			radix2 #(.width(width)) rd_st4_214  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[214]), .rdlo_in(a4_wr[246]),  .coef_in(coef[352]), .rdup_out(a5_wr[214]), .rdlo_out(a5_wr[246]));
			radix2 #(.width(width)) rd_st4_215  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[215]), .rdlo_in(a4_wr[247]),  .coef_in(coef[368]), .rdup_out(a5_wr[215]), .rdlo_out(a5_wr[247]));
			radix2 #(.width(width)) rd_st4_216  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[216]), .rdlo_in(a4_wr[248]),  .coef_in(coef[384]), .rdup_out(a5_wr[216]), .rdlo_out(a5_wr[248]));
			radix2 #(.width(width)) rd_st4_217  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[217]), .rdlo_in(a4_wr[249]),  .coef_in(coef[400]), .rdup_out(a5_wr[217]), .rdlo_out(a5_wr[249]));
			radix2 #(.width(width)) rd_st4_218  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[218]), .rdlo_in(a4_wr[250]),  .coef_in(coef[416]), .rdup_out(a5_wr[218]), .rdlo_out(a5_wr[250]));
			radix2 #(.width(width)) rd_st4_219  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[219]), .rdlo_in(a4_wr[251]),  .coef_in(coef[432]), .rdup_out(a5_wr[219]), .rdlo_out(a5_wr[251]));
			radix2 #(.width(width)) rd_st4_220  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[220]), .rdlo_in(a4_wr[252]),  .coef_in(coef[448]), .rdup_out(a5_wr[220]), .rdlo_out(a5_wr[252]));
			radix2 #(.width(width)) rd_st4_221  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[221]), .rdlo_in(a4_wr[253]),  .coef_in(coef[464]), .rdup_out(a5_wr[221]), .rdlo_out(a5_wr[253]));
			radix2 #(.width(width)) rd_st4_222  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[222]), .rdlo_in(a4_wr[254]),  .coef_in(coef[480]), .rdup_out(a5_wr[222]), .rdlo_out(a5_wr[254]));
			radix2 #(.width(width)) rd_st4_223  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[223]), .rdlo_in(a4_wr[255]),  .coef_in(coef[496]), .rdup_out(a5_wr[223]), .rdlo_out(a5_wr[255]));
			radix2 #(.width(width)) rd_st4_256  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[256]), .rdlo_in(a4_wr[288]),  .coef_in(coef[0]), .rdup_out(a5_wr[256]), .rdlo_out(a5_wr[288]));
			radix2 #(.width(width)) rd_st4_257  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[257]), .rdlo_in(a4_wr[289]),  .coef_in(coef[16]), .rdup_out(a5_wr[257]), .rdlo_out(a5_wr[289]));
			radix2 #(.width(width)) rd_st4_258  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[258]), .rdlo_in(a4_wr[290]),  .coef_in(coef[32]), .rdup_out(a5_wr[258]), .rdlo_out(a5_wr[290]));
			radix2 #(.width(width)) rd_st4_259  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[259]), .rdlo_in(a4_wr[291]),  .coef_in(coef[48]), .rdup_out(a5_wr[259]), .rdlo_out(a5_wr[291]));
			radix2 #(.width(width)) rd_st4_260  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[260]), .rdlo_in(a4_wr[292]),  .coef_in(coef[64]), .rdup_out(a5_wr[260]), .rdlo_out(a5_wr[292]));
			radix2 #(.width(width)) rd_st4_261  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[261]), .rdlo_in(a4_wr[293]),  .coef_in(coef[80]), .rdup_out(a5_wr[261]), .rdlo_out(a5_wr[293]));
			radix2 #(.width(width)) rd_st4_262  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[262]), .rdlo_in(a4_wr[294]),  .coef_in(coef[96]), .rdup_out(a5_wr[262]), .rdlo_out(a5_wr[294]));
			radix2 #(.width(width)) rd_st4_263  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[263]), .rdlo_in(a4_wr[295]),  .coef_in(coef[112]), .rdup_out(a5_wr[263]), .rdlo_out(a5_wr[295]));
			radix2 #(.width(width)) rd_st4_264  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[264]), .rdlo_in(a4_wr[296]),  .coef_in(coef[128]), .rdup_out(a5_wr[264]), .rdlo_out(a5_wr[296]));
			radix2 #(.width(width)) rd_st4_265  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[265]), .rdlo_in(a4_wr[297]),  .coef_in(coef[144]), .rdup_out(a5_wr[265]), .rdlo_out(a5_wr[297]));
			radix2 #(.width(width)) rd_st4_266  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[266]), .rdlo_in(a4_wr[298]),  .coef_in(coef[160]), .rdup_out(a5_wr[266]), .rdlo_out(a5_wr[298]));
			radix2 #(.width(width)) rd_st4_267  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[267]), .rdlo_in(a4_wr[299]),  .coef_in(coef[176]), .rdup_out(a5_wr[267]), .rdlo_out(a5_wr[299]));
			radix2 #(.width(width)) rd_st4_268  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[268]), .rdlo_in(a4_wr[300]),  .coef_in(coef[192]), .rdup_out(a5_wr[268]), .rdlo_out(a5_wr[300]));
			radix2 #(.width(width)) rd_st4_269  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[269]), .rdlo_in(a4_wr[301]),  .coef_in(coef[208]), .rdup_out(a5_wr[269]), .rdlo_out(a5_wr[301]));
			radix2 #(.width(width)) rd_st4_270  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[270]), .rdlo_in(a4_wr[302]),  .coef_in(coef[224]), .rdup_out(a5_wr[270]), .rdlo_out(a5_wr[302]));
			radix2 #(.width(width)) rd_st4_271  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[271]), .rdlo_in(a4_wr[303]),  .coef_in(coef[240]), .rdup_out(a5_wr[271]), .rdlo_out(a5_wr[303]));
			radix2 #(.width(width)) rd_st4_272  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[272]), .rdlo_in(a4_wr[304]),  .coef_in(coef[256]), .rdup_out(a5_wr[272]), .rdlo_out(a5_wr[304]));
			radix2 #(.width(width)) rd_st4_273  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[273]), .rdlo_in(a4_wr[305]),  .coef_in(coef[272]), .rdup_out(a5_wr[273]), .rdlo_out(a5_wr[305]));
			radix2 #(.width(width)) rd_st4_274  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[274]), .rdlo_in(a4_wr[306]),  .coef_in(coef[288]), .rdup_out(a5_wr[274]), .rdlo_out(a5_wr[306]));
			radix2 #(.width(width)) rd_st4_275  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[275]), .rdlo_in(a4_wr[307]),  .coef_in(coef[304]), .rdup_out(a5_wr[275]), .rdlo_out(a5_wr[307]));
			radix2 #(.width(width)) rd_st4_276  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[276]), .rdlo_in(a4_wr[308]),  .coef_in(coef[320]), .rdup_out(a5_wr[276]), .rdlo_out(a5_wr[308]));
			radix2 #(.width(width)) rd_st4_277  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[277]), .rdlo_in(a4_wr[309]),  .coef_in(coef[336]), .rdup_out(a5_wr[277]), .rdlo_out(a5_wr[309]));
			radix2 #(.width(width)) rd_st4_278  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[278]), .rdlo_in(a4_wr[310]),  .coef_in(coef[352]), .rdup_out(a5_wr[278]), .rdlo_out(a5_wr[310]));
			radix2 #(.width(width)) rd_st4_279  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[279]), .rdlo_in(a4_wr[311]),  .coef_in(coef[368]), .rdup_out(a5_wr[279]), .rdlo_out(a5_wr[311]));
			radix2 #(.width(width)) rd_st4_280  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[280]), .rdlo_in(a4_wr[312]),  .coef_in(coef[384]), .rdup_out(a5_wr[280]), .rdlo_out(a5_wr[312]));
			radix2 #(.width(width)) rd_st4_281  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[281]), .rdlo_in(a4_wr[313]),  .coef_in(coef[400]), .rdup_out(a5_wr[281]), .rdlo_out(a5_wr[313]));
			radix2 #(.width(width)) rd_st4_282  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[282]), .rdlo_in(a4_wr[314]),  .coef_in(coef[416]), .rdup_out(a5_wr[282]), .rdlo_out(a5_wr[314]));
			radix2 #(.width(width)) rd_st4_283  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[283]), .rdlo_in(a4_wr[315]),  .coef_in(coef[432]), .rdup_out(a5_wr[283]), .rdlo_out(a5_wr[315]));
			radix2 #(.width(width)) rd_st4_284  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[284]), .rdlo_in(a4_wr[316]),  .coef_in(coef[448]), .rdup_out(a5_wr[284]), .rdlo_out(a5_wr[316]));
			radix2 #(.width(width)) rd_st4_285  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[285]), .rdlo_in(a4_wr[317]),  .coef_in(coef[464]), .rdup_out(a5_wr[285]), .rdlo_out(a5_wr[317]));
			radix2 #(.width(width)) rd_st4_286  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[286]), .rdlo_in(a4_wr[318]),  .coef_in(coef[480]), .rdup_out(a5_wr[286]), .rdlo_out(a5_wr[318]));
			radix2 #(.width(width)) rd_st4_287  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[287]), .rdlo_in(a4_wr[319]),  .coef_in(coef[496]), .rdup_out(a5_wr[287]), .rdlo_out(a5_wr[319]));
			radix2 #(.width(width)) rd_st4_320  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[320]), .rdlo_in(a4_wr[352]),  .coef_in(coef[0]), .rdup_out(a5_wr[320]), .rdlo_out(a5_wr[352]));
			radix2 #(.width(width)) rd_st4_321  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[321]), .rdlo_in(a4_wr[353]),  .coef_in(coef[16]), .rdup_out(a5_wr[321]), .rdlo_out(a5_wr[353]));
			radix2 #(.width(width)) rd_st4_322  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[322]), .rdlo_in(a4_wr[354]),  .coef_in(coef[32]), .rdup_out(a5_wr[322]), .rdlo_out(a5_wr[354]));
			radix2 #(.width(width)) rd_st4_323  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[323]), .rdlo_in(a4_wr[355]),  .coef_in(coef[48]), .rdup_out(a5_wr[323]), .rdlo_out(a5_wr[355]));
			radix2 #(.width(width)) rd_st4_324  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[324]), .rdlo_in(a4_wr[356]),  .coef_in(coef[64]), .rdup_out(a5_wr[324]), .rdlo_out(a5_wr[356]));
			radix2 #(.width(width)) rd_st4_325  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[325]), .rdlo_in(a4_wr[357]),  .coef_in(coef[80]), .rdup_out(a5_wr[325]), .rdlo_out(a5_wr[357]));
			radix2 #(.width(width)) rd_st4_326  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[326]), .rdlo_in(a4_wr[358]),  .coef_in(coef[96]), .rdup_out(a5_wr[326]), .rdlo_out(a5_wr[358]));
			radix2 #(.width(width)) rd_st4_327  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[327]), .rdlo_in(a4_wr[359]),  .coef_in(coef[112]), .rdup_out(a5_wr[327]), .rdlo_out(a5_wr[359]));
			radix2 #(.width(width)) rd_st4_328  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[328]), .rdlo_in(a4_wr[360]),  .coef_in(coef[128]), .rdup_out(a5_wr[328]), .rdlo_out(a5_wr[360]));
			radix2 #(.width(width)) rd_st4_329  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[329]), .rdlo_in(a4_wr[361]),  .coef_in(coef[144]), .rdup_out(a5_wr[329]), .rdlo_out(a5_wr[361]));
			radix2 #(.width(width)) rd_st4_330  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[330]), .rdlo_in(a4_wr[362]),  .coef_in(coef[160]), .rdup_out(a5_wr[330]), .rdlo_out(a5_wr[362]));
			radix2 #(.width(width)) rd_st4_331  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[331]), .rdlo_in(a4_wr[363]),  .coef_in(coef[176]), .rdup_out(a5_wr[331]), .rdlo_out(a5_wr[363]));
			radix2 #(.width(width)) rd_st4_332  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[332]), .rdlo_in(a4_wr[364]),  .coef_in(coef[192]), .rdup_out(a5_wr[332]), .rdlo_out(a5_wr[364]));
			radix2 #(.width(width)) rd_st4_333  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[333]), .rdlo_in(a4_wr[365]),  .coef_in(coef[208]), .rdup_out(a5_wr[333]), .rdlo_out(a5_wr[365]));
			radix2 #(.width(width)) rd_st4_334  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[334]), .rdlo_in(a4_wr[366]),  .coef_in(coef[224]), .rdup_out(a5_wr[334]), .rdlo_out(a5_wr[366]));
			radix2 #(.width(width)) rd_st4_335  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[335]), .rdlo_in(a4_wr[367]),  .coef_in(coef[240]), .rdup_out(a5_wr[335]), .rdlo_out(a5_wr[367]));
			radix2 #(.width(width)) rd_st4_336  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[336]), .rdlo_in(a4_wr[368]),  .coef_in(coef[256]), .rdup_out(a5_wr[336]), .rdlo_out(a5_wr[368]));
			radix2 #(.width(width)) rd_st4_337  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[337]), .rdlo_in(a4_wr[369]),  .coef_in(coef[272]), .rdup_out(a5_wr[337]), .rdlo_out(a5_wr[369]));
			radix2 #(.width(width)) rd_st4_338  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[338]), .rdlo_in(a4_wr[370]),  .coef_in(coef[288]), .rdup_out(a5_wr[338]), .rdlo_out(a5_wr[370]));
			radix2 #(.width(width)) rd_st4_339  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[339]), .rdlo_in(a4_wr[371]),  .coef_in(coef[304]), .rdup_out(a5_wr[339]), .rdlo_out(a5_wr[371]));
			radix2 #(.width(width)) rd_st4_340  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[340]), .rdlo_in(a4_wr[372]),  .coef_in(coef[320]), .rdup_out(a5_wr[340]), .rdlo_out(a5_wr[372]));
			radix2 #(.width(width)) rd_st4_341  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[341]), .rdlo_in(a4_wr[373]),  .coef_in(coef[336]), .rdup_out(a5_wr[341]), .rdlo_out(a5_wr[373]));
			radix2 #(.width(width)) rd_st4_342  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[342]), .rdlo_in(a4_wr[374]),  .coef_in(coef[352]), .rdup_out(a5_wr[342]), .rdlo_out(a5_wr[374]));
			radix2 #(.width(width)) rd_st4_343  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[343]), .rdlo_in(a4_wr[375]),  .coef_in(coef[368]), .rdup_out(a5_wr[343]), .rdlo_out(a5_wr[375]));
			radix2 #(.width(width)) rd_st4_344  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[344]), .rdlo_in(a4_wr[376]),  .coef_in(coef[384]), .rdup_out(a5_wr[344]), .rdlo_out(a5_wr[376]));
			radix2 #(.width(width)) rd_st4_345  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[345]), .rdlo_in(a4_wr[377]),  .coef_in(coef[400]), .rdup_out(a5_wr[345]), .rdlo_out(a5_wr[377]));
			radix2 #(.width(width)) rd_st4_346  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[346]), .rdlo_in(a4_wr[378]),  .coef_in(coef[416]), .rdup_out(a5_wr[346]), .rdlo_out(a5_wr[378]));
			radix2 #(.width(width)) rd_st4_347  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[347]), .rdlo_in(a4_wr[379]),  .coef_in(coef[432]), .rdup_out(a5_wr[347]), .rdlo_out(a5_wr[379]));
			radix2 #(.width(width)) rd_st4_348  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[348]), .rdlo_in(a4_wr[380]),  .coef_in(coef[448]), .rdup_out(a5_wr[348]), .rdlo_out(a5_wr[380]));
			radix2 #(.width(width)) rd_st4_349  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[349]), .rdlo_in(a4_wr[381]),  .coef_in(coef[464]), .rdup_out(a5_wr[349]), .rdlo_out(a5_wr[381]));
			radix2 #(.width(width)) rd_st4_350  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[350]), .rdlo_in(a4_wr[382]),  .coef_in(coef[480]), .rdup_out(a5_wr[350]), .rdlo_out(a5_wr[382]));
			radix2 #(.width(width)) rd_st4_351  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[351]), .rdlo_in(a4_wr[383]),  .coef_in(coef[496]), .rdup_out(a5_wr[351]), .rdlo_out(a5_wr[383]));
			radix2 #(.width(width)) rd_st4_384  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[384]), .rdlo_in(a4_wr[416]),  .coef_in(coef[0]), .rdup_out(a5_wr[384]), .rdlo_out(a5_wr[416]));
			radix2 #(.width(width)) rd_st4_385  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[385]), .rdlo_in(a4_wr[417]),  .coef_in(coef[16]), .rdup_out(a5_wr[385]), .rdlo_out(a5_wr[417]));
			radix2 #(.width(width)) rd_st4_386  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[386]), .rdlo_in(a4_wr[418]),  .coef_in(coef[32]), .rdup_out(a5_wr[386]), .rdlo_out(a5_wr[418]));
			radix2 #(.width(width)) rd_st4_387  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[387]), .rdlo_in(a4_wr[419]),  .coef_in(coef[48]), .rdup_out(a5_wr[387]), .rdlo_out(a5_wr[419]));
			radix2 #(.width(width)) rd_st4_388  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[388]), .rdlo_in(a4_wr[420]),  .coef_in(coef[64]), .rdup_out(a5_wr[388]), .rdlo_out(a5_wr[420]));
			radix2 #(.width(width)) rd_st4_389  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[389]), .rdlo_in(a4_wr[421]),  .coef_in(coef[80]), .rdup_out(a5_wr[389]), .rdlo_out(a5_wr[421]));
			radix2 #(.width(width)) rd_st4_390  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[390]), .rdlo_in(a4_wr[422]),  .coef_in(coef[96]), .rdup_out(a5_wr[390]), .rdlo_out(a5_wr[422]));
			radix2 #(.width(width)) rd_st4_391  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[391]), .rdlo_in(a4_wr[423]),  .coef_in(coef[112]), .rdup_out(a5_wr[391]), .rdlo_out(a5_wr[423]));
			radix2 #(.width(width)) rd_st4_392  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[392]), .rdlo_in(a4_wr[424]),  .coef_in(coef[128]), .rdup_out(a5_wr[392]), .rdlo_out(a5_wr[424]));
			radix2 #(.width(width)) rd_st4_393  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[393]), .rdlo_in(a4_wr[425]),  .coef_in(coef[144]), .rdup_out(a5_wr[393]), .rdlo_out(a5_wr[425]));
			radix2 #(.width(width)) rd_st4_394  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[394]), .rdlo_in(a4_wr[426]),  .coef_in(coef[160]), .rdup_out(a5_wr[394]), .rdlo_out(a5_wr[426]));
			radix2 #(.width(width)) rd_st4_395  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[395]), .rdlo_in(a4_wr[427]),  .coef_in(coef[176]), .rdup_out(a5_wr[395]), .rdlo_out(a5_wr[427]));
			radix2 #(.width(width)) rd_st4_396  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[396]), .rdlo_in(a4_wr[428]),  .coef_in(coef[192]), .rdup_out(a5_wr[396]), .rdlo_out(a5_wr[428]));
			radix2 #(.width(width)) rd_st4_397  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[397]), .rdlo_in(a4_wr[429]),  .coef_in(coef[208]), .rdup_out(a5_wr[397]), .rdlo_out(a5_wr[429]));
			radix2 #(.width(width)) rd_st4_398  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[398]), .rdlo_in(a4_wr[430]),  .coef_in(coef[224]), .rdup_out(a5_wr[398]), .rdlo_out(a5_wr[430]));
			radix2 #(.width(width)) rd_st4_399  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[399]), .rdlo_in(a4_wr[431]),  .coef_in(coef[240]), .rdup_out(a5_wr[399]), .rdlo_out(a5_wr[431]));
			radix2 #(.width(width)) rd_st4_400  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[400]), .rdlo_in(a4_wr[432]),  .coef_in(coef[256]), .rdup_out(a5_wr[400]), .rdlo_out(a5_wr[432]));
			radix2 #(.width(width)) rd_st4_401  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[401]), .rdlo_in(a4_wr[433]),  .coef_in(coef[272]), .rdup_out(a5_wr[401]), .rdlo_out(a5_wr[433]));
			radix2 #(.width(width)) rd_st4_402  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[402]), .rdlo_in(a4_wr[434]),  .coef_in(coef[288]), .rdup_out(a5_wr[402]), .rdlo_out(a5_wr[434]));
			radix2 #(.width(width)) rd_st4_403  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[403]), .rdlo_in(a4_wr[435]),  .coef_in(coef[304]), .rdup_out(a5_wr[403]), .rdlo_out(a5_wr[435]));
			radix2 #(.width(width)) rd_st4_404  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[404]), .rdlo_in(a4_wr[436]),  .coef_in(coef[320]), .rdup_out(a5_wr[404]), .rdlo_out(a5_wr[436]));
			radix2 #(.width(width)) rd_st4_405  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[405]), .rdlo_in(a4_wr[437]),  .coef_in(coef[336]), .rdup_out(a5_wr[405]), .rdlo_out(a5_wr[437]));
			radix2 #(.width(width)) rd_st4_406  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[406]), .rdlo_in(a4_wr[438]),  .coef_in(coef[352]), .rdup_out(a5_wr[406]), .rdlo_out(a5_wr[438]));
			radix2 #(.width(width)) rd_st4_407  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[407]), .rdlo_in(a4_wr[439]),  .coef_in(coef[368]), .rdup_out(a5_wr[407]), .rdlo_out(a5_wr[439]));
			radix2 #(.width(width)) rd_st4_408  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[408]), .rdlo_in(a4_wr[440]),  .coef_in(coef[384]), .rdup_out(a5_wr[408]), .rdlo_out(a5_wr[440]));
			radix2 #(.width(width)) rd_st4_409  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[409]), .rdlo_in(a4_wr[441]),  .coef_in(coef[400]), .rdup_out(a5_wr[409]), .rdlo_out(a5_wr[441]));
			radix2 #(.width(width)) rd_st4_410  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[410]), .rdlo_in(a4_wr[442]),  .coef_in(coef[416]), .rdup_out(a5_wr[410]), .rdlo_out(a5_wr[442]));
			radix2 #(.width(width)) rd_st4_411  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[411]), .rdlo_in(a4_wr[443]),  .coef_in(coef[432]), .rdup_out(a5_wr[411]), .rdlo_out(a5_wr[443]));
			radix2 #(.width(width)) rd_st4_412  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[412]), .rdlo_in(a4_wr[444]),  .coef_in(coef[448]), .rdup_out(a5_wr[412]), .rdlo_out(a5_wr[444]));
			radix2 #(.width(width)) rd_st4_413  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[413]), .rdlo_in(a4_wr[445]),  .coef_in(coef[464]), .rdup_out(a5_wr[413]), .rdlo_out(a5_wr[445]));
			radix2 #(.width(width)) rd_st4_414  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[414]), .rdlo_in(a4_wr[446]),  .coef_in(coef[480]), .rdup_out(a5_wr[414]), .rdlo_out(a5_wr[446]));
			radix2 #(.width(width)) rd_st4_415  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[415]), .rdlo_in(a4_wr[447]),  .coef_in(coef[496]), .rdup_out(a5_wr[415]), .rdlo_out(a5_wr[447]));
			radix2 #(.width(width)) rd_st4_448  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[448]), .rdlo_in(a4_wr[480]),  .coef_in(coef[0]), .rdup_out(a5_wr[448]), .rdlo_out(a5_wr[480]));
			radix2 #(.width(width)) rd_st4_449  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[449]), .rdlo_in(a4_wr[481]),  .coef_in(coef[16]), .rdup_out(a5_wr[449]), .rdlo_out(a5_wr[481]));
			radix2 #(.width(width)) rd_st4_450  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[450]), .rdlo_in(a4_wr[482]),  .coef_in(coef[32]), .rdup_out(a5_wr[450]), .rdlo_out(a5_wr[482]));
			radix2 #(.width(width)) rd_st4_451  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[451]), .rdlo_in(a4_wr[483]),  .coef_in(coef[48]), .rdup_out(a5_wr[451]), .rdlo_out(a5_wr[483]));
			radix2 #(.width(width)) rd_st4_452  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[452]), .rdlo_in(a4_wr[484]),  .coef_in(coef[64]), .rdup_out(a5_wr[452]), .rdlo_out(a5_wr[484]));
			radix2 #(.width(width)) rd_st4_453  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[453]), .rdlo_in(a4_wr[485]),  .coef_in(coef[80]), .rdup_out(a5_wr[453]), .rdlo_out(a5_wr[485]));
			radix2 #(.width(width)) rd_st4_454  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[454]), .rdlo_in(a4_wr[486]),  .coef_in(coef[96]), .rdup_out(a5_wr[454]), .rdlo_out(a5_wr[486]));
			radix2 #(.width(width)) rd_st4_455  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[455]), .rdlo_in(a4_wr[487]),  .coef_in(coef[112]), .rdup_out(a5_wr[455]), .rdlo_out(a5_wr[487]));
			radix2 #(.width(width)) rd_st4_456  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[456]), .rdlo_in(a4_wr[488]),  .coef_in(coef[128]), .rdup_out(a5_wr[456]), .rdlo_out(a5_wr[488]));
			radix2 #(.width(width)) rd_st4_457  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[457]), .rdlo_in(a4_wr[489]),  .coef_in(coef[144]), .rdup_out(a5_wr[457]), .rdlo_out(a5_wr[489]));
			radix2 #(.width(width)) rd_st4_458  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[458]), .rdlo_in(a4_wr[490]),  .coef_in(coef[160]), .rdup_out(a5_wr[458]), .rdlo_out(a5_wr[490]));
			radix2 #(.width(width)) rd_st4_459  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[459]), .rdlo_in(a4_wr[491]),  .coef_in(coef[176]), .rdup_out(a5_wr[459]), .rdlo_out(a5_wr[491]));
			radix2 #(.width(width)) rd_st4_460  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[460]), .rdlo_in(a4_wr[492]),  .coef_in(coef[192]), .rdup_out(a5_wr[460]), .rdlo_out(a5_wr[492]));
			radix2 #(.width(width)) rd_st4_461  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[461]), .rdlo_in(a4_wr[493]),  .coef_in(coef[208]), .rdup_out(a5_wr[461]), .rdlo_out(a5_wr[493]));
			radix2 #(.width(width)) rd_st4_462  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[462]), .rdlo_in(a4_wr[494]),  .coef_in(coef[224]), .rdup_out(a5_wr[462]), .rdlo_out(a5_wr[494]));
			radix2 #(.width(width)) rd_st4_463  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[463]), .rdlo_in(a4_wr[495]),  .coef_in(coef[240]), .rdup_out(a5_wr[463]), .rdlo_out(a5_wr[495]));
			radix2 #(.width(width)) rd_st4_464  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[464]), .rdlo_in(a4_wr[496]),  .coef_in(coef[256]), .rdup_out(a5_wr[464]), .rdlo_out(a5_wr[496]));
			radix2 #(.width(width)) rd_st4_465  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[465]), .rdlo_in(a4_wr[497]),  .coef_in(coef[272]), .rdup_out(a5_wr[465]), .rdlo_out(a5_wr[497]));
			radix2 #(.width(width)) rd_st4_466  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[466]), .rdlo_in(a4_wr[498]),  .coef_in(coef[288]), .rdup_out(a5_wr[466]), .rdlo_out(a5_wr[498]));
			radix2 #(.width(width)) rd_st4_467  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[467]), .rdlo_in(a4_wr[499]),  .coef_in(coef[304]), .rdup_out(a5_wr[467]), .rdlo_out(a5_wr[499]));
			radix2 #(.width(width)) rd_st4_468  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[468]), .rdlo_in(a4_wr[500]),  .coef_in(coef[320]), .rdup_out(a5_wr[468]), .rdlo_out(a5_wr[500]));
			radix2 #(.width(width)) rd_st4_469  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[469]), .rdlo_in(a4_wr[501]),  .coef_in(coef[336]), .rdup_out(a5_wr[469]), .rdlo_out(a5_wr[501]));
			radix2 #(.width(width)) rd_st4_470  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[470]), .rdlo_in(a4_wr[502]),  .coef_in(coef[352]), .rdup_out(a5_wr[470]), .rdlo_out(a5_wr[502]));
			radix2 #(.width(width)) rd_st4_471  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[471]), .rdlo_in(a4_wr[503]),  .coef_in(coef[368]), .rdup_out(a5_wr[471]), .rdlo_out(a5_wr[503]));
			radix2 #(.width(width)) rd_st4_472  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[472]), .rdlo_in(a4_wr[504]),  .coef_in(coef[384]), .rdup_out(a5_wr[472]), .rdlo_out(a5_wr[504]));
			radix2 #(.width(width)) rd_st4_473  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[473]), .rdlo_in(a4_wr[505]),  .coef_in(coef[400]), .rdup_out(a5_wr[473]), .rdlo_out(a5_wr[505]));
			radix2 #(.width(width)) rd_st4_474  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[474]), .rdlo_in(a4_wr[506]),  .coef_in(coef[416]), .rdup_out(a5_wr[474]), .rdlo_out(a5_wr[506]));
			radix2 #(.width(width)) rd_st4_475  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[475]), .rdlo_in(a4_wr[507]),  .coef_in(coef[432]), .rdup_out(a5_wr[475]), .rdlo_out(a5_wr[507]));
			radix2 #(.width(width)) rd_st4_476  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[476]), .rdlo_in(a4_wr[508]),  .coef_in(coef[448]), .rdup_out(a5_wr[476]), .rdlo_out(a5_wr[508]));
			radix2 #(.width(width)) rd_st4_477  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[477]), .rdlo_in(a4_wr[509]),  .coef_in(coef[464]), .rdup_out(a5_wr[477]), .rdlo_out(a5_wr[509]));
			radix2 #(.width(width)) rd_st4_478  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[478]), .rdlo_in(a4_wr[510]),  .coef_in(coef[480]), .rdup_out(a5_wr[478]), .rdlo_out(a5_wr[510]));
			radix2 #(.width(width)) rd_st4_479  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[479]), .rdlo_in(a4_wr[511]),  .coef_in(coef[496]), .rdup_out(a5_wr[479]), .rdlo_out(a5_wr[511]));
			radix2 #(.width(width)) rd_st4_512  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[512]), .rdlo_in(a4_wr[544]),  .coef_in(coef[0]), .rdup_out(a5_wr[512]), .rdlo_out(a5_wr[544]));
			radix2 #(.width(width)) rd_st4_513  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[513]), .rdlo_in(a4_wr[545]),  .coef_in(coef[16]), .rdup_out(a5_wr[513]), .rdlo_out(a5_wr[545]));
			radix2 #(.width(width)) rd_st4_514  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[514]), .rdlo_in(a4_wr[546]),  .coef_in(coef[32]), .rdup_out(a5_wr[514]), .rdlo_out(a5_wr[546]));
			radix2 #(.width(width)) rd_st4_515  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[515]), .rdlo_in(a4_wr[547]),  .coef_in(coef[48]), .rdup_out(a5_wr[515]), .rdlo_out(a5_wr[547]));
			radix2 #(.width(width)) rd_st4_516  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[516]), .rdlo_in(a4_wr[548]),  .coef_in(coef[64]), .rdup_out(a5_wr[516]), .rdlo_out(a5_wr[548]));
			radix2 #(.width(width)) rd_st4_517  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[517]), .rdlo_in(a4_wr[549]),  .coef_in(coef[80]), .rdup_out(a5_wr[517]), .rdlo_out(a5_wr[549]));
			radix2 #(.width(width)) rd_st4_518  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[518]), .rdlo_in(a4_wr[550]),  .coef_in(coef[96]), .rdup_out(a5_wr[518]), .rdlo_out(a5_wr[550]));
			radix2 #(.width(width)) rd_st4_519  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[519]), .rdlo_in(a4_wr[551]),  .coef_in(coef[112]), .rdup_out(a5_wr[519]), .rdlo_out(a5_wr[551]));
			radix2 #(.width(width)) rd_st4_520  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[520]), .rdlo_in(a4_wr[552]),  .coef_in(coef[128]), .rdup_out(a5_wr[520]), .rdlo_out(a5_wr[552]));
			radix2 #(.width(width)) rd_st4_521  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[521]), .rdlo_in(a4_wr[553]),  .coef_in(coef[144]), .rdup_out(a5_wr[521]), .rdlo_out(a5_wr[553]));
			radix2 #(.width(width)) rd_st4_522  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[522]), .rdlo_in(a4_wr[554]),  .coef_in(coef[160]), .rdup_out(a5_wr[522]), .rdlo_out(a5_wr[554]));
			radix2 #(.width(width)) rd_st4_523  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[523]), .rdlo_in(a4_wr[555]),  .coef_in(coef[176]), .rdup_out(a5_wr[523]), .rdlo_out(a5_wr[555]));
			radix2 #(.width(width)) rd_st4_524  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[524]), .rdlo_in(a4_wr[556]),  .coef_in(coef[192]), .rdup_out(a5_wr[524]), .rdlo_out(a5_wr[556]));
			radix2 #(.width(width)) rd_st4_525  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[525]), .rdlo_in(a4_wr[557]),  .coef_in(coef[208]), .rdup_out(a5_wr[525]), .rdlo_out(a5_wr[557]));
			radix2 #(.width(width)) rd_st4_526  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[526]), .rdlo_in(a4_wr[558]),  .coef_in(coef[224]), .rdup_out(a5_wr[526]), .rdlo_out(a5_wr[558]));
			radix2 #(.width(width)) rd_st4_527  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[527]), .rdlo_in(a4_wr[559]),  .coef_in(coef[240]), .rdup_out(a5_wr[527]), .rdlo_out(a5_wr[559]));
			radix2 #(.width(width)) rd_st4_528  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[528]), .rdlo_in(a4_wr[560]),  .coef_in(coef[256]), .rdup_out(a5_wr[528]), .rdlo_out(a5_wr[560]));
			radix2 #(.width(width)) rd_st4_529  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[529]), .rdlo_in(a4_wr[561]),  .coef_in(coef[272]), .rdup_out(a5_wr[529]), .rdlo_out(a5_wr[561]));
			radix2 #(.width(width)) rd_st4_530  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[530]), .rdlo_in(a4_wr[562]),  .coef_in(coef[288]), .rdup_out(a5_wr[530]), .rdlo_out(a5_wr[562]));
			radix2 #(.width(width)) rd_st4_531  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[531]), .rdlo_in(a4_wr[563]),  .coef_in(coef[304]), .rdup_out(a5_wr[531]), .rdlo_out(a5_wr[563]));
			radix2 #(.width(width)) rd_st4_532  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[532]), .rdlo_in(a4_wr[564]),  .coef_in(coef[320]), .rdup_out(a5_wr[532]), .rdlo_out(a5_wr[564]));
			radix2 #(.width(width)) rd_st4_533  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[533]), .rdlo_in(a4_wr[565]),  .coef_in(coef[336]), .rdup_out(a5_wr[533]), .rdlo_out(a5_wr[565]));
			radix2 #(.width(width)) rd_st4_534  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[534]), .rdlo_in(a4_wr[566]),  .coef_in(coef[352]), .rdup_out(a5_wr[534]), .rdlo_out(a5_wr[566]));
			radix2 #(.width(width)) rd_st4_535  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[535]), .rdlo_in(a4_wr[567]),  .coef_in(coef[368]), .rdup_out(a5_wr[535]), .rdlo_out(a5_wr[567]));
			radix2 #(.width(width)) rd_st4_536  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[536]), .rdlo_in(a4_wr[568]),  .coef_in(coef[384]), .rdup_out(a5_wr[536]), .rdlo_out(a5_wr[568]));
			radix2 #(.width(width)) rd_st4_537  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[537]), .rdlo_in(a4_wr[569]),  .coef_in(coef[400]), .rdup_out(a5_wr[537]), .rdlo_out(a5_wr[569]));
			radix2 #(.width(width)) rd_st4_538  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[538]), .rdlo_in(a4_wr[570]),  .coef_in(coef[416]), .rdup_out(a5_wr[538]), .rdlo_out(a5_wr[570]));
			radix2 #(.width(width)) rd_st4_539  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[539]), .rdlo_in(a4_wr[571]),  .coef_in(coef[432]), .rdup_out(a5_wr[539]), .rdlo_out(a5_wr[571]));
			radix2 #(.width(width)) rd_st4_540  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[540]), .rdlo_in(a4_wr[572]),  .coef_in(coef[448]), .rdup_out(a5_wr[540]), .rdlo_out(a5_wr[572]));
			radix2 #(.width(width)) rd_st4_541  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[541]), .rdlo_in(a4_wr[573]),  .coef_in(coef[464]), .rdup_out(a5_wr[541]), .rdlo_out(a5_wr[573]));
			radix2 #(.width(width)) rd_st4_542  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[542]), .rdlo_in(a4_wr[574]),  .coef_in(coef[480]), .rdup_out(a5_wr[542]), .rdlo_out(a5_wr[574]));
			radix2 #(.width(width)) rd_st4_543  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[543]), .rdlo_in(a4_wr[575]),  .coef_in(coef[496]), .rdup_out(a5_wr[543]), .rdlo_out(a5_wr[575]));
			radix2 #(.width(width)) rd_st4_576  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[576]), .rdlo_in(a4_wr[608]),  .coef_in(coef[0]), .rdup_out(a5_wr[576]), .rdlo_out(a5_wr[608]));
			radix2 #(.width(width)) rd_st4_577  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[577]), .rdlo_in(a4_wr[609]),  .coef_in(coef[16]), .rdup_out(a5_wr[577]), .rdlo_out(a5_wr[609]));
			radix2 #(.width(width)) rd_st4_578  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[578]), .rdlo_in(a4_wr[610]),  .coef_in(coef[32]), .rdup_out(a5_wr[578]), .rdlo_out(a5_wr[610]));
			radix2 #(.width(width)) rd_st4_579  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[579]), .rdlo_in(a4_wr[611]),  .coef_in(coef[48]), .rdup_out(a5_wr[579]), .rdlo_out(a5_wr[611]));
			radix2 #(.width(width)) rd_st4_580  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[580]), .rdlo_in(a4_wr[612]),  .coef_in(coef[64]), .rdup_out(a5_wr[580]), .rdlo_out(a5_wr[612]));
			radix2 #(.width(width)) rd_st4_581  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[581]), .rdlo_in(a4_wr[613]),  .coef_in(coef[80]), .rdup_out(a5_wr[581]), .rdlo_out(a5_wr[613]));
			radix2 #(.width(width)) rd_st4_582  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[582]), .rdlo_in(a4_wr[614]),  .coef_in(coef[96]), .rdup_out(a5_wr[582]), .rdlo_out(a5_wr[614]));
			radix2 #(.width(width)) rd_st4_583  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[583]), .rdlo_in(a4_wr[615]),  .coef_in(coef[112]), .rdup_out(a5_wr[583]), .rdlo_out(a5_wr[615]));
			radix2 #(.width(width)) rd_st4_584  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[584]), .rdlo_in(a4_wr[616]),  .coef_in(coef[128]), .rdup_out(a5_wr[584]), .rdlo_out(a5_wr[616]));
			radix2 #(.width(width)) rd_st4_585  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[585]), .rdlo_in(a4_wr[617]),  .coef_in(coef[144]), .rdup_out(a5_wr[585]), .rdlo_out(a5_wr[617]));
			radix2 #(.width(width)) rd_st4_586  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[586]), .rdlo_in(a4_wr[618]),  .coef_in(coef[160]), .rdup_out(a5_wr[586]), .rdlo_out(a5_wr[618]));
			radix2 #(.width(width)) rd_st4_587  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[587]), .rdlo_in(a4_wr[619]),  .coef_in(coef[176]), .rdup_out(a5_wr[587]), .rdlo_out(a5_wr[619]));
			radix2 #(.width(width)) rd_st4_588  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[588]), .rdlo_in(a4_wr[620]),  .coef_in(coef[192]), .rdup_out(a5_wr[588]), .rdlo_out(a5_wr[620]));
			radix2 #(.width(width)) rd_st4_589  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[589]), .rdlo_in(a4_wr[621]),  .coef_in(coef[208]), .rdup_out(a5_wr[589]), .rdlo_out(a5_wr[621]));
			radix2 #(.width(width)) rd_st4_590  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[590]), .rdlo_in(a4_wr[622]),  .coef_in(coef[224]), .rdup_out(a5_wr[590]), .rdlo_out(a5_wr[622]));
			radix2 #(.width(width)) rd_st4_591  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[591]), .rdlo_in(a4_wr[623]),  .coef_in(coef[240]), .rdup_out(a5_wr[591]), .rdlo_out(a5_wr[623]));
			radix2 #(.width(width)) rd_st4_592  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[592]), .rdlo_in(a4_wr[624]),  .coef_in(coef[256]), .rdup_out(a5_wr[592]), .rdlo_out(a5_wr[624]));
			radix2 #(.width(width)) rd_st4_593  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[593]), .rdlo_in(a4_wr[625]),  .coef_in(coef[272]), .rdup_out(a5_wr[593]), .rdlo_out(a5_wr[625]));
			radix2 #(.width(width)) rd_st4_594  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[594]), .rdlo_in(a4_wr[626]),  .coef_in(coef[288]), .rdup_out(a5_wr[594]), .rdlo_out(a5_wr[626]));
			radix2 #(.width(width)) rd_st4_595  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[595]), .rdlo_in(a4_wr[627]),  .coef_in(coef[304]), .rdup_out(a5_wr[595]), .rdlo_out(a5_wr[627]));
			radix2 #(.width(width)) rd_st4_596  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[596]), .rdlo_in(a4_wr[628]),  .coef_in(coef[320]), .rdup_out(a5_wr[596]), .rdlo_out(a5_wr[628]));
			radix2 #(.width(width)) rd_st4_597  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[597]), .rdlo_in(a4_wr[629]),  .coef_in(coef[336]), .rdup_out(a5_wr[597]), .rdlo_out(a5_wr[629]));
			radix2 #(.width(width)) rd_st4_598  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[598]), .rdlo_in(a4_wr[630]),  .coef_in(coef[352]), .rdup_out(a5_wr[598]), .rdlo_out(a5_wr[630]));
			radix2 #(.width(width)) rd_st4_599  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[599]), .rdlo_in(a4_wr[631]),  .coef_in(coef[368]), .rdup_out(a5_wr[599]), .rdlo_out(a5_wr[631]));
			radix2 #(.width(width)) rd_st4_600  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[600]), .rdlo_in(a4_wr[632]),  .coef_in(coef[384]), .rdup_out(a5_wr[600]), .rdlo_out(a5_wr[632]));
			radix2 #(.width(width)) rd_st4_601  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[601]), .rdlo_in(a4_wr[633]),  .coef_in(coef[400]), .rdup_out(a5_wr[601]), .rdlo_out(a5_wr[633]));
			radix2 #(.width(width)) rd_st4_602  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[602]), .rdlo_in(a4_wr[634]),  .coef_in(coef[416]), .rdup_out(a5_wr[602]), .rdlo_out(a5_wr[634]));
			radix2 #(.width(width)) rd_st4_603  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[603]), .rdlo_in(a4_wr[635]),  .coef_in(coef[432]), .rdup_out(a5_wr[603]), .rdlo_out(a5_wr[635]));
			radix2 #(.width(width)) rd_st4_604  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[604]), .rdlo_in(a4_wr[636]),  .coef_in(coef[448]), .rdup_out(a5_wr[604]), .rdlo_out(a5_wr[636]));
			radix2 #(.width(width)) rd_st4_605  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[605]), .rdlo_in(a4_wr[637]),  .coef_in(coef[464]), .rdup_out(a5_wr[605]), .rdlo_out(a5_wr[637]));
			radix2 #(.width(width)) rd_st4_606  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[606]), .rdlo_in(a4_wr[638]),  .coef_in(coef[480]), .rdup_out(a5_wr[606]), .rdlo_out(a5_wr[638]));
			radix2 #(.width(width)) rd_st4_607  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[607]), .rdlo_in(a4_wr[639]),  .coef_in(coef[496]), .rdup_out(a5_wr[607]), .rdlo_out(a5_wr[639]));
			radix2 #(.width(width)) rd_st4_640  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[640]), .rdlo_in(a4_wr[672]),  .coef_in(coef[0]), .rdup_out(a5_wr[640]), .rdlo_out(a5_wr[672]));
			radix2 #(.width(width)) rd_st4_641  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[641]), .rdlo_in(a4_wr[673]),  .coef_in(coef[16]), .rdup_out(a5_wr[641]), .rdlo_out(a5_wr[673]));
			radix2 #(.width(width)) rd_st4_642  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[642]), .rdlo_in(a4_wr[674]),  .coef_in(coef[32]), .rdup_out(a5_wr[642]), .rdlo_out(a5_wr[674]));
			radix2 #(.width(width)) rd_st4_643  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[643]), .rdlo_in(a4_wr[675]),  .coef_in(coef[48]), .rdup_out(a5_wr[643]), .rdlo_out(a5_wr[675]));
			radix2 #(.width(width)) rd_st4_644  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[644]), .rdlo_in(a4_wr[676]),  .coef_in(coef[64]), .rdup_out(a5_wr[644]), .rdlo_out(a5_wr[676]));
			radix2 #(.width(width)) rd_st4_645  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[645]), .rdlo_in(a4_wr[677]),  .coef_in(coef[80]), .rdup_out(a5_wr[645]), .rdlo_out(a5_wr[677]));
			radix2 #(.width(width)) rd_st4_646  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[646]), .rdlo_in(a4_wr[678]),  .coef_in(coef[96]), .rdup_out(a5_wr[646]), .rdlo_out(a5_wr[678]));
			radix2 #(.width(width)) rd_st4_647  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[647]), .rdlo_in(a4_wr[679]),  .coef_in(coef[112]), .rdup_out(a5_wr[647]), .rdlo_out(a5_wr[679]));
			radix2 #(.width(width)) rd_st4_648  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[648]), .rdlo_in(a4_wr[680]),  .coef_in(coef[128]), .rdup_out(a5_wr[648]), .rdlo_out(a5_wr[680]));
			radix2 #(.width(width)) rd_st4_649  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[649]), .rdlo_in(a4_wr[681]),  .coef_in(coef[144]), .rdup_out(a5_wr[649]), .rdlo_out(a5_wr[681]));
			radix2 #(.width(width)) rd_st4_650  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[650]), .rdlo_in(a4_wr[682]),  .coef_in(coef[160]), .rdup_out(a5_wr[650]), .rdlo_out(a5_wr[682]));
			radix2 #(.width(width)) rd_st4_651  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[651]), .rdlo_in(a4_wr[683]),  .coef_in(coef[176]), .rdup_out(a5_wr[651]), .rdlo_out(a5_wr[683]));
			radix2 #(.width(width)) rd_st4_652  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[652]), .rdlo_in(a4_wr[684]),  .coef_in(coef[192]), .rdup_out(a5_wr[652]), .rdlo_out(a5_wr[684]));
			radix2 #(.width(width)) rd_st4_653  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[653]), .rdlo_in(a4_wr[685]),  .coef_in(coef[208]), .rdup_out(a5_wr[653]), .rdlo_out(a5_wr[685]));
			radix2 #(.width(width)) rd_st4_654  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[654]), .rdlo_in(a4_wr[686]),  .coef_in(coef[224]), .rdup_out(a5_wr[654]), .rdlo_out(a5_wr[686]));
			radix2 #(.width(width)) rd_st4_655  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[655]), .rdlo_in(a4_wr[687]),  .coef_in(coef[240]), .rdup_out(a5_wr[655]), .rdlo_out(a5_wr[687]));
			radix2 #(.width(width)) rd_st4_656  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[656]), .rdlo_in(a4_wr[688]),  .coef_in(coef[256]), .rdup_out(a5_wr[656]), .rdlo_out(a5_wr[688]));
			radix2 #(.width(width)) rd_st4_657  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[657]), .rdlo_in(a4_wr[689]),  .coef_in(coef[272]), .rdup_out(a5_wr[657]), .rdlo_out(a5_wr[689]));
			radix2 #(.width(width)) rd_st4_658  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[658]), .rdlo_in(a4_wr[690]),  .coef_in(coef[288]), .rdup_out(a5_wr[658]), .rdlo_out(a5_wr[690]));
			radix2 #(.width(width)) rd_st4_659  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[659]), .rdlo_in(a4_wr[691]),  .coef_in(coef[304]), .rdup_out(a5_wr[659]), .rdlo_out(a5_wr[691]));
			radix2 #(.width(width)) rd_st4_660  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[660]), .rdlo_in(a4_wr[692]),  .coef_in(coef[320]), .rdup_out(a5_wr[660]), .rdlo_out(a5_wr[692]));
			radix2 #(.width(width)) rd_st4_661  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[661]), .rdlo_in(a4_wr[693]),  .coef_in(coef[336]), .rdup_out(a5_wr[661]), .rdlo_out(a5_wr[693]));
			radix2 #(.width(width)) rd_st4_662  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[662]), .rdlo_in(a4_wr[694]),  .coef_in(coef[352]), .rdup_out(a5_wr[662]), .rdlo_out(a5_wr[694]));
			radix2 #(.width(width)) rd_st4_663  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[663]), .rdlo_in(a4_wr[695]),  .coef_in(coef[368]), .rdup_out(a5_wr[663]), .rdlo_out(a5_wr[695]));
			radix2 #(.width(width)) rd_st4_664  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[664]), .rdlo_in(a4_wr[696]),  .coef_in(coef[384]), .rdup_out(a5_wr[664]), .rdlo_out(a5_wr[696]));
			radix2 #(.width(width)) rd_st4_665  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[665]), .rdlo_in(a4_wr[697]),  .coef_in(coef[400]), .rdup_out(a5_wr[665]), .rdlo_out(a5_wr[697]));
			radix2 #(.width(width)) rd_st4_666  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[666]), .rdlo_in(a4_wr[698]),  .coef_in(coef[416]), .rdup_out(a5_wr[666]), .rdlo_out(a5_wr[698]));
			radix2 #(.width(width)) rd_st4_667  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[667]), .rdlo_in(a4_wr[699]),  .coef_in(coef[432]), .rdup_out(a5_wr[667]), .rdlo_out(a5_wr[699]));
			radix2 #(.width(width)) rd_st4_668  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[668]), .rdlo_in(a4_wr[700]),  .coef_in(coef[448]), .rdup_out(a5_wr[668]), .rdlo_out(a5_wr[700]));
			radix2 #(.width(width)) rd_st4_669  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[669]), .rdlo_in(a4_wr[701]),  .coef_in(coef[464]), .rdup_out(a5_wr[669]), .rdlo_out(a5_wr[701]));
			radix2 #(.width(width)) rd_st4_670  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[670]), .rdlo_in(a4_wr[702]),  .coef_in(coef[480]), .rdup_out(a5_wr[670]), .rdlo_out(a5_wr[702]));
			radix2 #(.width(width)) rd_st4_671  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[671]), .rdlo_in(a4_wr[703]),  .coef_in(coef[496]), .rdup_out(a5_wr[671]), .rdlo_out(a5_wr[703]));
			radix2 #(.width(width)) rd_st4_704  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[704]), .rdlo_in(a4_wr[736]),  .coef_in(coef[0]), .rdup_out(a5_wr[704]), .rdlo_out(a5_wr[736]));
			radix2 #(.width(width)) rd_st4_705  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[705]), .rdlo_in(a4_wr[737]),  .coef_in(coef[16]), .rdup_out(a5_wr[705]), .rdlo_out(a5_wr[737]));
			radix2 #(.width(width)) rd_st4_706  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[706]), .rdlo_in(a4_wr[738]),  .coef_in(coef[32]), .rdup_out(a5_wr[706]), .rdlo_out(a5_wr[738]));
			radix2 #(.width(width)) rd_st4_707  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[707]), .rdlo_in(a4_wr[739]),  .coef_in(coef[48]), .rdup_out(a5_wr[707]), .rdlo_out(a5_wr[739]));
			radix2 #(.width(width)) rd_st4_708  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[708]), .rdlo_in(a4_wr[740]),  .coef_in(coef[64]), .rdup_out(a5_wr[708]), .rdlo_out(a5_wr[740]));
			radix2 #(.width(width)) rd_st4_709  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[709]), .rdlo_in(a4_wr[741]),  .coef_in(coef[80]), .rdup_out(a5_wr[709]), .rdlo_out(a5_wr[741]));
			radix2 #(.width(width)) rd_st4_710  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[710]), .rdlo_in(a4_wr[742]),  .coef_in(coef[96]), .rdup_out(a5_wr[710]), .rdlo_out(a5_wr[742]));
			radix2 #(.width(width)) rd_st4_711  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[711]), .rdlo_in(a4_wr[743]),  .coef_in(coef[112]), .rdup_out(a5_wr[711]), .rdlo_out(a5_wr[743]));
			radix2 #(.width(width)) rd_st4_712  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[712]), .rdlo_in(a4_wr[744]),  .coef_in(coef[128]), .rdup_out(a5_wr[712]), .rdlo_out(a5_wr[744]));
			radix2 #(.width(width)) rd_st4_713  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[713]), .rdlo_in(a4_wr[745]),  .coef_in(coef[144]), .rdup_out(a5_wr[713]), .rdlo_out(a5_wr[745]));
			radix2 #(.width(width)) rd_st4_714  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[714]), .rdlo_in(a4_wr[746]),  .coef_in(coef[160]), .rdup_out(a5_wr[714]), .rdlo_out(a5_wr[746]));
			radix2 #(.width(width)) rd_st4_715  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[715]), .rdlo_in(a4_wr[747]),  .coef_in(coef[176]), .rdup_out(a5_wr[715]), .rdlo_out(a5_wr[747]));
			radix2 #(.width(width)) rd_st4_716  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[716]), .rdlo_in(a4_wr[748]),  .coef_in(coef[192]), .rdup_out(a5_wr[716]), .rdlo_out(a5_wr[748]));
			radix2 #(.width(width)) rd_st4_717  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[717]), .rdlo_in(a4_wr[749]),  .coef_in(coef[208]), .rdup_out(a5_wr[717]), .rdlo_out(a5_wr[749]));
			radix2 #(.width(width)) rd_st4_718  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[718]), .rdlo_in(a4_wr[750]),  .coef_in(coef[224]), .rdup_out(a5_wr[718]), .rdlo_out(a5_wr[750]));
			radix2 #(.width(width)) rd_st4_719  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[719]), .rdlo_in(a4_wr[751]),  .coef_in(coef[240]), .rdup_out(a5_wr[719]), .rdlo_out(a5_wr[751]));
			radix2 #(.width(width)) rd_st4_720  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[720]), .rdlo_in(a4_wr[752]),  .coef_in(coef[256]), .rdup_out(a5_wr[720]), .rdlo_out(a5_wr[752]));
			radix2 #(.width(width)) rd_st4_721  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[721]), .rdlo_in(a4_wr[753]),  .coef_in(coef[272]), .rdup_out(a5_wr[721]), .rdlo_out(a5_wr[753]));
			radix2 #(.width(width)) rd_st4_722  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[722]), .rdlo_in(a4_wr[754]),  .coef_in(coef[288]), .rdup_out(a5_wr[722]), .rdlo_out(a5_wr[754]));
			radix2 #(.width(width)) rd_st4_723  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[723]), .rdlo_in(a4_wr[755]),  .coef_in(coef[304]), .rdup_out(a5_wr[723]), .rdlo_out(a5_wr[755]));
			radix2 #(.width(width)) rd_st4_724  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[724]), .rdlo_in(a4_wr[756]),  .coef_in(coef[320]), .rdup_out(a5_wr[724]), .rdlo_out(a5_wr[756]));
			radix2 #(.width(width)) rd_st4_725  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[725]), .rdlo_in(a4_wr[757]),  .coef_in(coef[336]), .rdup_out(a5_wr[725]), .rdlo_out(a5_wr[757]));
			radix2 #(.width(width)) rd_st4_726  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[726]), .rdlo_in(a4_wr[758]),  .coef_in(coef[352]), .rdup_out(a5_wr[726]), .rdlo_out(a5_wr[758]));
			radix2 #(.width(width)) rd_st4_727  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[727]), .rdlo_in(a4_wr[759]),  .coef_in(coef[368]), .rdup_out(a5_wr[727]), .rdlo_out(a5_wr[759]));
			radix2 #(.width(width)) rd_st4_728  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[728]), .rdlo_in(a4_wr[760]),  .coef_in(coef[384]), .rdup_out(a5_wr[728]), .rdlo_out(a5_wr[760]));
			radix2 #(.width(width)) rd_st4_729  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[729]), .rdlo_in(a4_wr[761]),  .coef_in(coef[400]), .rdup_out(a5_wr[729]), .rdlo_out(a5_wr[761]));
			radix2 #(.width(width)) rd_st4_730  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[730]), .rdlo_in(a4_wr[762]),  .coef_in(coef[416]), .rdup_out(a5_wr[730]), .rdlo_out(a5_wr[762]));
			radix2 #(.width(width)) rd_st4_731  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[731]), .rdlo_in(a4_wr[763]),  .coef_in(coef[432]), .rdup_out(a5_wr[731]), .rdlo_out(a5_wr[763]));
			radix2 #(.width(width)) rd_st4_732  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[732]), .rdlo_in(a4_wr[764]),  .coef_in(coef[448]), .rdup_out(a5_wr[732]), .rdlo_out(a5_wr[764]));
			radix2 #(.width(width)) rd_st4_733  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[733]), .rdlo_in(a4_wr[765]),  .coef_in(coef[464]), .rdup_out(a5_wr[733]), .rdlo_out(a5_wr[765]));
			radix2 #(.width(width)) rd_st4_734  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[734]), .rdlo_in(a4_wr[766]),  .coef_in(coef[480]), .rdup_out(a5_wr[734]), .rdlo_out(a5_wr[766]));
			radix2 #(.width(width)) rd_st4_735  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[735]), .rdlo_in(a4_wr[767]),  .coef_in(coef[496]), .rdup_out(a5_wr[735]), .rdlo_out(a5_wr[767]));
			radix2 #(.width(width)) rd_st4_768  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[768]), .rdlo_in(a4_wr[800]),  .coef_in(coef[0]), .rdup_out(a5_wr[768]), .rdlo_out(a5_wr[800]));
			radix2 #(.width(width)) rd_st4_769  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[769]), .rdlo_in(a4_wr[801]),  .coef_in(coef[16]), .rdup_out(a5_wr[769]), .rdlo_out(a5_wr[801]));
			radix2 #(.width(width)) rd_st4_770  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[770]), .rdlo_in(a4_wr[802]),  .coef_in(coef[32]), .rdup_out(a5_wr[770]), .rdlo_out(a5_wr[802]));
			radix2 #(.width(width)) rd_st4_771  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[771]), .rdlo_in(a4_wr[803]),  .coef_in(coef[48]), .rdup_out(a5_wr[771]), .rdlo_out(a5_wr[803]));
			radix2 #(.width(width)) rd_st4_772  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[772]), .rdlo_in(a4_wr[804]),  .coef_in(coef[64]), .rdup_out(a5_wr[772]), .rdlo_out(a5_wr[804]));
			radix2 #(.width(width)) rd_st4_773  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[773]), .rdlo_in(a4_wr[805]),  .coef_in(coef[80]), .rdup_out(a5_wr[773]), .rdlo_out(a5_wr[805]));
			radix2 #(.width(width)) rd_st4_774  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[774]), .rdlo_in(a4_wr[806]),  .coef_in(coef[96]), .rdup_out(a5_wr[774]), .rdlo_out(a5_wr[806]));
			radix2 #(.width(width)) rd_st4_775  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[775]), .rdlo_in(a4_wr[807]),  .coef_in(coef[112]), .rdup_out(a5_wr[775]), .rdlo_out(a5_wr[807]));
			radix2 #(.width(width)) rd_st4_776  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[776]), .rdlo_in(a4_wr[808]),  .coef_in(coef[128]), .rdup_out(a5_wr[776]), .rdlo_out(a5_wr[808]));
			radix2 #(.width(width)) rd_st4_777  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[777]), .rdlo_in(a4_wr[809]),  .coef_in(coef[144]), .rdup_out(a5_wr[777]), .rdlo_out(a5_wr[809]));
			radix2 #(.width(width)) rd_st4_778  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[778]), .rdlo_in(a4_wr[810]),  .coef_in(coef[160]), .rdup_out(a5_wr[778]), .rdlo_out(a5_wr[810]));
			radix2 #(.width(width)) rd_st4_779  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[779]), .rdlo_in(a4_wr[811]),  .coef_in(coef[176]), .rdup_out(a5_wr[779]), .rdlo_out(a5_wr[811]));
			radix2 #(.width(width)) rd_st4_780  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[780]), .rdlo_in(a4_wr[812]),  .coef_in(coef[192]), .rdup_out(a5_wr[780]), .rdlo_out(a5_wr[812]));
			radix2 #(.width(width)) rd_st4_781  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[781]), .rdlo_in(a4_wr[813]),  .coef_in(coef[208]), .rdup_out(a5_wr[781]), .rdlo_out(a5_wr[813]));
			radix2 #(.width(width)) rd_st4_782  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[782]), .rdlo_in(a4_wr[814]),  .coef_in(coef[224]), .rdup_out(a5_wr[782]), .rdlo_out(a5_wr[814]));
			radix2 #(.width(width)) rd_st4_783  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[783]), .rdlo_in(a4_wr[815]),  .coef_in(coef[240]), .rdup_out(a5_wr[783]), .rdlo_out(a5_wr[815]));
			radix2 #(.width(width)) rd_st4_784  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[784]), .rdlo_in(a4_wr[816]),  .coef_in(coef[256]), .rdup_out(a5_wr[784]), .rdlo_out(a5_wr[816]));
			radix2 #(.width(width)) rd_st4_785  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[785]), .rdlo_in(a4_wr[817]),  .coef_in(coef[272]), .rdup_out(a5_wr[785]), .rdlo_out(a5_wr[817]));
			radix2 #(.width(width)) rd_st4_786  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[786]), .rdlo_in(a4_wr[818]),  .coef_in(coef[288]), .rdup_out(a5_wr[786]), .rdlo_out(a5_wr[818]));
			radix2 #(.width(width)) rd_st4_787  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[787]), .rdlo_in(a4_wr[819]),  .coef_in(coef[304]), .rdup_out(a5_wr[787]), .rdlo_out(a5_wr[819]));
			radix2 #(.width(width)) rd_st4_788  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[788]), .rdlo_in(a4_wr[820]),  .coef_in(coef[320]), .rdup_out(a5_wr[788]), .rdlo_out(a5_wr[820]));
			radix2 #(.width(width)) rd_st4_789  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[789]), .rdlo_in(a4_wr[821]),  .coef_in(coef[336]), .rdup_out(a5_wr[789]), .rdlo_out(a5_wr[821]));
			radix2 #(.width(width)) rd_st4_790  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[790]), .rdlo_in(a4_wr[822]),  .coef_in(coef[352]), .rdup_out(a5_wr[790]), .rdlo_out(a5_wr[822]));
			radix2 #(.width(width)) rd_st4_791  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[791]), .rdlo_in(a4_wr[823]),  .coef_in(coef[368]), .rdup_out(a5_wr[791]), .rdlo_out(a5_wr[823]));
			radix2 #(.width(width)) rd_st4_792  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[792]), .rdlo_in(a4_wr[824]),  .coef_in(coef[384]), .rdup_out(a5_wr[792]), .rdlo_out(a5_wr[824]));
			radix2 #(.width(width)) rd_st4_793  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[793]), .rdlo_in(a4_wr[825]),  .coef_in(coef[400]), .rdup_out(a5_wr[793]), .rdlo_out(a5_wr[825]));
			radix2 #(.width(width)) rd_st4_794  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[794]), .rdlo_in(a4_wr[826]),  .coef_in(coef[416]), .rdup_out(a5_wr[794]), .rdlo_out(a5_wr[826]));
			radix2 #(.width(width)) rd_st4_795  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[795]), .rdlo_in(a4_wr[827]),  .coef_in(coef[432]), .rdup_out(a5_wr[795]), .rdlo_out(a5_wr[827]));
			radix2 #(.width(width)) rd_st4_796  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[796]), .rdlo_in(a4_wr[828]),  .coef_in(coef[448]), .rdup_out(a5_wr[796]), .rdlo_out(a5_wr[828]));
			radix2 #(.width(width)) rd_st4_797  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[797]), .rdlo_in(a4_wr[829]),  .coef_in(coef[464]), .rdup_out(a5_wr[797]), .rdlo_out(a5_wr[829]));
			radix2 #(.width(width)) rd_st4_798  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[798]), .rdlo_in(a4_wr[830]),  .coef_in(coef[480]), .rdup_out(a5_wr[798]), .rdlo_out(a5_wr[830]));
			radix2 #(.width(width)) rd_st4_799  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[799]), .rdlo_in(a4_wr[831]),  .coef_in(coef[496]), .rdup_out(a5_wr[799]), .rdlo_out(a5_wr[831]));
			radix2 #(.width(width)) rd_st4_832  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[832]), .rdlo_in(a4_wr[864]),  .coef_in(coef[0]), .rdup_out(a5_wr[832]), .rdlo_out(a5_wr[864]));
			radix2 #(.width(width)) rd_st4_833  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[833]), .rdlo_in(a4_wr[865]),  .coef_in(coef[16]), .rdup_out(a5_wr[833]), .rdlo_out(a5_wr[865]));
			radix2 #(.width(width)) rd_st4_834  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[834]), .rdlo_in(a4_wr[866]),  .coef_in(coef[32]), .rdup_out(a5_wr[834]), .rdlo_out(a5_wr[866]));
			radix2 #(.width(width)) rd_st4_835  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[835]), .rdlo_in(a4_wr[867]),  .coef_in(coef[48]), .rdup_out(a5_wr[835]), .rdlo_out(a5_wr[867]));
			radix2 #(.width(width)) rd_st4_836  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[836]), .rdlo_in(a4_wr[868]),  .coef_in(coef[64]), .rdup_out(a5_wr[836]), .rdlo_out(a5_wr[868]));
			radix2 #(.width(width)) rd_st4_837  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[837]), .rdlo_in(a4_wr[869]),  .coef_in(coef[80]), .rdup_out(a5_wr[837]), .rdlo_out(a5_wr[869]));
			radix2 #(.width(width)) rd_st4_838  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[838]), .rdlo_in(a4_wr[870]),  .coef_in(coef[96]), .rdup_out(a5_wr[838]), .rdlo_out(a5_wr[870]));
			radix2 #(.width(width)) rd_st4_839  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[839]), .rdlo_in(a4_wr[871]),  .coef_in(coef[112]), .rdup_out(a5_wr[839]), .rdlo_out(a5_wr[871]));
			radix2 #(.width(width)) rd_st4_840  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[840]), .rdlo_in(a4_wr[872]),  .coef_in(coef[128]), .rdup_out(a5_wr[840]), .rdlo_out(a5_wr[872]));
			radix2 #(.width(width)) rd_st4_841  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[841]), .rdlo_in(a4_wr[873]),  .coef_in(coef[144]), .rdup_out(a5_wr[841]), .rdlo_out(a5_wr[873]));
			radix2 #(.width(width)) rd_st4_842  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[842]), .rdlo_in(a4_wr[874]),  .coef_in(coef[160]), .rdup_out(a5_wr[842]), .rdlo_out(a5_wr[874]));
			radix2 #(.width(width)) rd_st4_843  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[843]), .rdlo_in(a4_wr[875]),  .coef_in(coef[176]), .rdup_out(a5_wr[843]), .rdlo_out(a5_wr[875]));
			radix2 #(.width(width)) rd_st4_844  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[844]), .rdlo_in(a4_wr[876]),  .coef_in(coef[192]), .rdup_out(a5_wr[844]), .rdlo_out(a5_wr[876]));
			radix2 #(.width(width)) rd_st4_845  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[845]), .rdlo_in(a4_wr[877]),  .coef_in(coef[208]), .rdup_out(a5_wr[845]), .rdlo_out(a5_wr[877]));
			radix2 #(.width(width)) rd_st4_846  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[846]), .rdlo_in(a4_wr[878]),  .coef_in(coef[224]), .rdup_out(a5_wr[846]), .rdlo_out(a5_wr[878]));
			radix2 #(.width(width)) rd_st4_847  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[847]), .rdlo_in(a4_wr[879]),  .coef_in(coef[240]), .rdup_out(a5_wr[847]), .rdlo_out(a5_wr[879]));
			radix2 #(.width(width)) rd_st4_848  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[848]), .rdlo_in(a4_wr[880]),  .coef_in(coef[256]), .rdup_out(a5_wr[848]), .rdlo_out(a5_wr[880]));
			radix2 #(.width(width)) rd_st4_849  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[849]), .rdlo_in(a4_wr[881]),  .coef_in(coef[272]), .rdup_out(a5_wr[849]), .rdlo_out(a5_wr[881]));
			radix2 #(.width(width)) rd_st4_850  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[850]), .rdlo_in(a4_wr[882]),  .coef_in(coef[288]), .rdup_out(a5_wr[850]), .rdlo_out(a5_wr[882]));
			radix2 #(.width(width)) rd_st4_851  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[851]), .rdlo_in(a4_wr[883]),  .coef_in(coef[304]), .rdup_out(a5_wr[851]), .rdlo_out(a5_wr[883]));
			radix2 #(.width(width)) rd_st4_852  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[852]), .rdlo_in(a4_wr[884]),  .coef_in(coef[320]), .rdup_out(a5_wr[852]), .rdlo_out(a5_wr[884]));
			radix2 #(.width(width)) rd_st4_853  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[853]), .rdlo_in(a4_wr[885]),  .coef_in(coef[336]), .rdup_out(a5_wr[853]), .rdlo_out(a5_wr[885]));
			radix2 #(.width(width)) rd_st4_854  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[854]), .rdlo_in(a4_wr[886]),  .coef_in(coef[352]), .rdup_out(a5_wr[854]), .rdlo_out(a5_wr[886]));
			radix2 #(.width(width)) rd_st4_855  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[855]), .rdlo_in(a4_wr[887]),  .coef_in(coef[368]), .rdup_out(a5_wr[855]), .rdlo_out(a5_wr[887]));
			radix2 #(.width(width)) rd_st4_856  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[856]), .rdlo_in(a4_wr[888]),  .coef_in(coef[384]), .rdup_out(a5_wr[856]), .rdlo_out(a5_wr[888]));
			radix2 #(.width(width)) rd_st4_857  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[857]), .rdlo_in(a4_wr[889]),  .coef_in(coef[400]), .rdup_out(a5_wr[857]), .rdlo_out(a5_wr[889]));
			radix2 #(.width(width)) rd_st4_858  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[858]), .rdlo_in(a4_wr[890]),  .coef_in(coef[416]), .rdup_out(a5_wr[858]), .rdlo_out(a5_wr[890]));
			radix2 #(.width(width)) rd_st4_859  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[859]), .rdlo_in(a4_wr[891]),  .coef_in(coef[432]), .rdup_out(a5_wr[859]), .rdlo_out(a5_wr[891]));
			radix2 #(.width(width)) rd_st4_860  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[860]), .rdlo_in(a4_wr[892]),  .coef_in(coef[448]), .rdup_out(a5_wr[860]), .rdlo_out(a5_wr[892]));
			radix2 #(.width(width)) rd_st4_861  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[861]), .rdlo_in(a4_wr[893]),  .coef_in(coef[464]), .rdup_out(a5_wr[861]), .rdlo_out(a5_wr[893]));
			radix2 #(.width(width)) rd_st4_862  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[862]), .rdlo_in(a4_wr[894]),  .coef_in(coef[480]), .rdup_out(a5_wr[862]), .rdlo_out(a5_wr[894]));
			radix2 #(.width(width)) rd_st4_863  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[863]), .rdlo_in(a4_wr[895]),  .coef_in(coef[496]), .rdup_out(a5_wr[863]), .rdlo_out(a5_wr[895]));
			radix2 #(.width(width)) rd_st4_896  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[896]), .rdlo_in(a4_wr[928]),  .coef_in(coef[0]), .rdup_out(a5_wr[896]), .rdlo_out(a5_wr[928]));
			radix2 #(.width(width)) rd_st4_897  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[897]), .rdlo_in(a4_wr[929]),  .coef_in(coef[16]), .rdup_out(a5_wr[897]), .rdlo_out(a5_wr[929]));
			radix2 #(.width(width)) rd_st4_898  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[898]), .rdlo_in(a4_wr[930]),  .coef_in(coef[32]), .rdup_out(a5_wr[898]), .rdlo_out(a5_wr[930]));
			radix2 #(.width(width)) rd_st4_899  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[899]), .rdlo_in(a4_wr[931]),  .coef_in(coef[48]), .rdup_out(a5_wr[899]), .rdlo_out(a5_wr[931]));
			radix2 #(.width(width)) rd_st4_900  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[900]), .rdlo_in(a4_wr[932]),  .coef_in(coef[64]), .rdup_out(a5_wr[900]), .rdlo_out(a5_wr[932]));
			radix2 #(.width(width)) rd_st4_901  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[901]), .rdlo_in(a4_wr[933]),  .coef_in(coef[80]), .rdup_out(a5_wr[901]), .rdlo_out(a5_wr[933]));
			radix2 #(.width(width)) rd_st4_902  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[902]), .rdlo_in(a4_wr[934]),  .coef_in(coef[96]), .rdup_out(a5_wr[902]), .rdlo_out(a5_wr[934]));
			radix2 #(.width(width)) rd_st4_903  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[903]), .rdlo_in(a4_wr[935]),  .coef_in(coef[112]), .rdup_out(a5_wr[903]), .rdlo_out(a5_wr[935]));
			radix2 #(.width(width)) rd_st4_904  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[904]), .rdlo_in(a4_wr[936]),  .coef_in(coef[128]), .rdup_out(a5_wr[904]), .rdlo_out(a5_wr[936]));
			radix2 #(.width(width)) rd_st4_905  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[905]), .rdlo_in(a4_wr[937]),  .coef_in(coef[144]), .rdup_out(a5_wr[905]), .rdlo_out(a5_wr[937]));
			radix2 #(.width(width)) rd_st4_906  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[906]), .rdlo_in(a4_wr[938]),  .coef_in(coef[160]), .rdup_out(a5_wr[906]), .rdlo_out(a5_wr[938]));
			radix2 #(.width(width)) rd_st4_907  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[907]), .rdlo_in(a4_wr[939]),  .coef_in(coef[176]), .rdup_out(a5_wr[907]), .rdlo_out(a5_wr[939]));
			radix2 #(.width(width)) rd_st4_908  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[908]), .rdlo_in(a4_wr[940]),  .coef_in(coef[192]), .rdup_out(a5_wr[908]), .rdlo_out(a5_wr[940]));
			radix2 #(.width(width)) rd_st4_909  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[909]), .rdlo_in(a4_wr[941]),  .coef_in(coef[208]), .rdup_out(a5_wr[909]), .rdlo_out(a5_wr[941]));
			radix2 #(.width(width)) rd_st4_910  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[910]), .rdlo_in(a4_wr[942]),  .coef_in(coef[224]), .rdup_out(a5_wr[910]), .rdlo_out(a5_wr[942]));
			radix2 #(.width(width)) rd_st4_911  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[911]), .rdlo_in(a4_wr[943]),  .coef_in(coef[240]), .rdup_out(a5_wr[911]), .rdlo_out(a5_wr[943]));
			radix2 #(.width(width)) rd_st4_912  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[912]), .rdlo_in(a4_wr[944]),  .coef_in(coef[256]), .rdup_out(a5_wr[912]), .rdlo_out(a5_wr[944]));
			radix2 #(.width(width)) rd_st4_913  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[913]), .rdlo_in(a4_wr[945]),  .coef_in(coef[272]), .rdup_out(a5_wr[913]), .rdlo_out(a5_wr[945]));
			radix2 #(.width(width)) rd_st4_914  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[914]), .rdlo_in(a4_wr[946]),  .coef_in(coef[288]), .rdup_out(a5_wr[914]), .rdlo_out(a5_wr[946]));
			radix2 #(.width(width)) rd_st4_915  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[915]), .rdlo_in(a4_wr[947]),  .coef_in(coef[304]), .rdup_out(a5_wr[915]), .rdlo_out(a5_wr[947]));
			radix2 #(.width(width)) rd_st4_916  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[916]), .rdlo_in(a4_wr[948]),  .coef_in(coef[320]), .rdup_out(a5_wr[916]), .rdlo_out(a5_wr[948]));
			radix2 #(.width(width)) rd_st4_917  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[917]), .rdlo_in(a4_wr[949]),  .coef_in(coef[336]), .rdup_out(a5_wr[917]), .rdlo_out(a5_wr[949]));
			radix2 #(.width(width)) rd_st4_918  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[918]), .rdlo_in(a4_wr[950]),  .coef_in(coef[352]), .rdup_out(a5_wr[918]), .rdlo_out(a5_wr[950]));
			radix2 #(.width(width)) rd_st4_919  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[919]), .rdlo_in(a4_wr[951]),  .coef_in(coef[368]), .rdup_out(a5_wr[919]), .rdlo_out(a5_wr[951]));
			radix2 #(.width(width)) rd_st4_920  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[920]), .rdlo_in(a4_wr[952]),  .coef_in(coef[384]), .rdup_out(a5_wr[920]), .rdlo_out(a5_wr[952]));
			radix2 #(.width(width)) rd_st4_921  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[921]), .rdlo_in(a4_wr[953]),  .coef_in(coef[400]), .rdup_out(a5_wr[921]), .rdlo_out(a5_wr[953]));
			radix2 #(.width(width)) rd_st4_922  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[922]), .rdlo_in(a4_wr[954]),  .coef_in(coef[416]), .rdup_out(a5_wr[922]), .rdlo_out(a5_wr[954]));
			radix2 #(.width(width)) rd_st4_923  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[923]), .rdlo_in(a4_wr[955]),  .coef_in(coef[432]), .rdup_out(a5_wr[923]), .rdlo_out(a5_wr[955]));
			radix2 #(.width(width)) rd_st4_924  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[924]), .rdlo_in(a4_wr[956]),  .coef_in(coef[448]), .rdup_out(a5_wr[924]), .rdlo_out(a5_wr[956]));
			radix2 #(.width(width)) rd_st4_925  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[925]), .rdlo_in(a4_wr[957]),  .coef_in(coef[464]), .rdup_out(a5_wr[925]), .rdlo_out(a5_wr[957]));
			radix2 #(.width(width)) rd_st4_926  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[926]), .rdlo_in(a4_wr[958]),  .coef_in(coef[480]), .rdup_out(a5_wr[926]), .rdlo_out(a5_wr[958]));
			radix2 #(.width(width)) rd_st4_927  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[927]), .rdlo_in(a4_wr[959]),  .coef_in(coef[496]), .rdup_out(a5_wr[927]), .rdlo_out(a5_wr[959]));
			radix2 #(.width(width)) rd_st4_960  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[960]), .rdlo_in(a4_wr[992]),  .coef_in(coef[0]), .rdup_out(a5_wr[960]), .rdlo_out(a5_wr[992]));
			radix2 #(.width(width)) rd_st4_961  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[961]), .rdlo_in(a4_wr[993]),  .coef_in(coef[16]), .rdup_out(a5_wr[961]), .rdlo_out(a5_wr[993]));
			radix2 #(.width(width)) rd_st4_962  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[962]), .rdlo_in(a4_wr[994]),  .coef_in(coef[32]), .rdup_out(a5_wr[962]), .rdlo_out(a5_wr[994]));
			radix2 #(.width(width)) rd_st4_963  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[963]), .rdlo_in(a4_wr[995]),  .coef_in(coef[48]), .rdup_out(a5_wr[963]), .rdlo_out(a5_wr[995]));
			radix2 #(.width(width)) rd_st4_964  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[964]), .rdlo_in(a4_wr[996]),  .coef_in(coef[64]), .rdup_out(a5_wr[964]), .rdlo_out(a5_wr[996]));
			radix2 #(.width(width)) rd_st4_965  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[965]), .rdlo_in(a4_wr[997]),  .coef_in(coef[80]), .rdup_out(a5_wr[965]), .rdlo_out(a5_wr[997]));
			radix2 #(.width(width)) rd_st4_966  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[966]), .rdlo_in(a4_wr[998]),  .coef_in(coef[96]), .rdup_out(a5_wr[966]), .rdlo_out(a5_wr[998]));
			radix2 #(.width(width)) rd_st4_967  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[967]), .rdlo_in(a4_wr[999]),  .coef_in(coef[112]), .rdup_out(a5_wr[967]), .rdlo_out(a5_wr[999]));
			radix2 #(.width(width)) rd_st4_968  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[968]), .rdlo_in(a4_wr[1000]),  .coef_in(coef[128]), .rdup_out(a5_wr[968]), .rdlo_out(a5_wr[1000]));
			radix2 #(.width(width)) rd_st4_969  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[969]), .rdlo_in(a4_wr[1001]),  .coef_in(coef[144]), .rdup_out(a5_wr[969]), .rdlo_out(a5_wr[1001]));
			radix2 #(.width(width)) rd_st4_970  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[970]), .rdlo_in(a4_wr[1002]),  .coef_in(coef[160]), .rdup_out(a5_wr[970]), .rdlo_out(a5_wr[1002]));
			radix2 #(.width(width)) rd_st4_971  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[971]), .rdlo_in(a4_wr[1003]),  .coef_in(coef[176]), .rdup_out(a5_wr[971]), .rdlo_out(a5_wr[1003]));
			radix2 #(.width(width)) rd_st4_972  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[972]), .rdlo_in(a4_wr[1004]),  .coef_in(coef[192]), .rdup_out(a5_wr[972]), .rdlo_out(a5_wr[1004]));
			radix2 #(.width(width)) rd_st4_973  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[973]), .rdlo_in(a4_wr[1005]),  .coef_in(coef[208]), .rdup_out(a5_wr[973]), .rdlo_out(a5_wr[1005]));
			radix2 #(.width(width)) rd_st4_974  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[974]), .rdlo_in(a4_wr[1006]),  .coef_in(coef[224]), .rdup_out(a5_wr[974]), .rdlo_out(a5_wr[1006]));
			radix2 #(.width(width)) rd_st4_975  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[975]), .rdlo_in(a4_wr[1007]),  .coef_in(coef[240]), .rdup_out(a5_wr[975]), .rdlo_out(a5_wr[1007]));
			radix2 #(.width(width)) rd_st4_976  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[976]), .rdlo_in(a4_wr[1008]),  .coef_in(coef[256]), .rdup_out(a5_wr[976]), .rdlo_out(a5_wr[1008]));
			radix2 #(.width(width)) rd_st4_977  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[977]), .rdlo_in(a4_wr[1009]),  .coef_in(coef[272]), .rdup_out(a5_wr[977]), .rdlo_out(a5_wr[1009]));
			radix2 #(.width(width)) rd_st4_978  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[978]), .rdlo_in(a4_wr[1010]),  .coef_in(coef[288]), .rdup_out(a5_wr[978]), .rdlo_out(a5_wr[1010]));
			radix2 #(.width(width)) rd_st4_979  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[979]), .rdlo_in(a4_wr[1011]),  .coef_in(coef[304]), .rdup_out(a5_wr[979]), .rdlo_out(a5_wr[1011]));
			radix2 #(.width(width)) rd_st4_980  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[980]), .rdlo_in(a4_wr[1012]),  .coef_in(coef[320]), .rdup_out(a5_wr[980]), .rdlo_out(a5_wr[1012]));
			radix2 #(.width(width)) rd_st4_981  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[981]), .rdlo_in(a4_wr[1013]),  .coef_in(coef[336]), .rdup_out(a5_wr[981]), .rdlo_out(a5_wr[1013]));
			radix2 #(.width(width)) rd_st4_982  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[982]), .rdlo_in(a4_wr[1014]),  .coef_in(coef[352]), .rdup_out(a5_wr[982]), .rdlo_out(a5_wr[1014]));
			radix2 #(.width(width)) rd_st4_983  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[983]), .rdlo_in(a4_wr[1015]),  .coef_in(coef[368]), .rdup_out(a5_wr[983]), .rdlo_out(a5_wr[1015]));
			radix2 #(.width(width)) rd_st4_984  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[984]), .rdlo_in(a4_wr[1016]),  .coef_in(coef[384]), .rdup_out(a5_wr[984]), .rdlo_out(a5_wr[1016]));
			radix2 #(.width(width)) rd_st4_985  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[985]), .rdlo_in(a4_wr[1017]),  .coef_in(coef[400]), .rdup_out(a5_wr[985]), .rdlo_out(a5_wr[1017]));
			radix2 #(.width(width)) rd_st4_986  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[986]), .rdlo_in(a4_wr[1018]),  .coef_in(coef[416]), .rdup_out(a5_wr[986]), .rdlo_out(a5_wr[1018]));
			radix2 #(.width(width)) rd_st4_987  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[987]), .rdlo_in(a4_wr[1019]),  .coef_in(coef[432]), .rdup_out(a5_wr[987]), .rdlo_out(a5_wr[1019]));
			radix2 #(.width(width)) rd_st4_988  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[988]), .rdlo_in(a4_wr[1020]),  .coef_in(coef[448]), .rdup_out(a5_wr[988]), .rdlo_out(a5_wr[1020]));
			radix2 #(.width(width)) rd_st4_989  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[989]), .rdlo_in(a4_wr[1021]),  .coef_in(coef[464]), .rdup_out(a5_wr[989]), .rdlo_out(a5_wr[1021]));
			radix2 #(.width(width)) rd_st4_990  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[990]), .rdlo_in(a4_wr[1022]),  .coef_in(coef[480]), .rdup_out(a5_wr[990]), .rdlo_out(a5_wr[1022]));
			radix2 #(.width(width)) rd_st4_991  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[991]), .rdlo_in(a4_wr[1023]),  .coef_in(coef[496]), .rdup_out(a5_wr[991]), .rdlo_out(a5_wr[1023]));

		//--- radix stage 5
			radix2 #(.width(width)) rd_st5_0   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[0]), .rdlo_in(a5_wr[16]),  .coef_in(coef[0]), .rdup_out(a6_wr[0]), .rdlo_out(a6_wr[16]));
			radix2 #(.width(width)) rd_st5_1   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1]), .rdlo_in(a5_wr[17]),  .coef_in(coef[32]), .rdup_out(a6_wr[1]), .rdlo_out(a6_wr[17]));
			radix2 #(.width(width)) rd_st5_2   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[2]), .rdlo_in(a5_wr[18]),  .coef_in(coef[64]), .rdup_out(a6_wr[2]), .rdlo_out(a6_wr[18]));
			radix2 #(.width(width)) rd_st5_3   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[3]), .rdlo_in(a5_wr[19]),  .coef_in(coef[96]), .rdup_out(a6_wr[3]), .rdlo_out(a6_wr[19]));
			radix2 #(.width(width)) rd_st5_4   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[4]), .rdlo_in(a5_wr[20]),  .coef_in(coef[128]), .rdup_out(a6_wr[4]), .rdlo_out(a6_wr[20]));
			radix2 #(.width(width)) rd_st5_5   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[5]), .rdlo_in(a5_wr[21]),  .coef_in(coef[160]), .rdup_out(a6_wr[5]), .rdlo_out(a6_wr[21]));
			radix2 #(.width(width)) rd_st5_6   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[6]), .rdlo_in(a5_wr[22]),  .coef_in(coef[192]), .rdup_out(a6_wr[6]), .rdlo_out(a6_wr[22]));
			radix2 #(.width(width)) rd_st5_7   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[7]), .rdlo_in(a5_wr[23]),  .coef_in(coef[224]), .rdup_out(a6_wr[7]), .rdlo_out(a6_wr[23]));
			radix2 #(.width(width)) rd_st5_8   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[8]), .rdlo_in(a5_wr[24]),  .coef_in(coef[256]), .rdup_out(a6_wr[8]), .rdlo_out(a6_wr[24]));
			radix2 #(.width(width)) rd_st5_9   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[9]), .rdlo_in(a5_wr[25]),  .coef_in(coef[288]), .rdup_out(a6_wr[9]), .rdlo_out(a6_wr[25]));
			radix2 #(.width(width)) rd_st5_10  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[10]), .rdlo_in(a5_wr[26]),  .coef_in(coef[320]), .rdup_out(a6_wr[10]), .rdlo_out(a6_wr[26]));
			radix2 #(.width(width)) rd_st5_11  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[11]), .rdlo_in(a5_wr[27]),  .coef_in(coef[352]), .rdup_out(a6_wr[11]), .rdlo_out(a6_wr[27]));
			radix2 #(.width(width)) rd_st5_12  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[12]), .rdlo_in(a5_wr[28]),  .coef_in(coef[384]), .rdup_out(a6_wr[12]), .rdlo_out(a6_wr[28]));
			radix2 #(.width(width)) rd_st5_13  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[13]), .rdlo_in(a5_wr[29]),  .coef_in(coef[416]), .rdup_out(a6_wr[13]), .rdlo_out(a6_wr[29]));
			radix2 #(.width(width)) rd_st5_14  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[14]), .rdlo_in(a5_wr[30]),  .coef_in(coef[448]), .rdup_out(a6_wr[14]), .rdlo_out(a6_wr[30]));
			radix2 #(.width(width)) rd_st5_15  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[15]), .rdlo_in(a5_wr[31]),  .coef_in(coef[480]), .rdup_out(a6_wr[15]), .rdlo_out(a6_wr[31]));
			radix2 #(.width(width)) rd_st5_32  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[32]), .rdlo_in(a5_wr[48]),  .coef_in(coef[0]), .rdup_out(a6_wr[32]), .rdlo_out(a6_wr[48]));
			radix2 #(.width(width)) rd_st5_33  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[33]), .rdlo_in(a5_wr[49]),  .coef_in(coef[32]), .rdup_out(a6_wr[33]), .rdlo_out(a6_wr[49]));
			radix2 #(.width(width)) rd_st5_34  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[34]), .rdlo_in(a5_wr[50]),  .coef_in(coef[64]), .rdup_out(a6_wr[34]), .rdlo_out(a6_wr[50]));
			radix2 #(.width(width)) rd_st5_35  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[35]), .rdlo_in(a5_wr[51]),  .coef_in(coef[96]), .rdup_out(a6_wr[35]), .rdlo_out(a6_wr[51]));
			radix2 #(.width(width)) rd_st5_36  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[36]), .rdlo_in(a5_wr[52]),  .coef_in(coef[128]), .rdup_out(a6_wr[36]), .rdlo_out(a6_wr[52]));
			radix2 #(.width(width)) rd_st5_37  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[37]), .rdlo_in(a5_wr[53]),  .coef_in(coef[160]), .rdup_out(a6_wr[37]), .rdlo_out(a6_wr[53]));
			radix2 #(.width(width)) rd_st5_38  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[38]), .rdlo_in(a5_wr[54]),  .coef_in(coef[192]), .rdup_out(a6_wr[38]), .rdlo_out(a6_wr[54]));
			radix2 #(.width(width)) rd_st5_39  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[39]), .rdlo_in(a5_wr[55]),  .coef_in(coef[224]), .rdup_out(a6_wr[39]), .rdlo_out(a6_wr[55]));
			radix2 #(.width(width)) rd_st5_40  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[40]), .rdlo_in(a5_wr[56]),  .coef_in(coef[256]), .rdup_out(a6_wr[40]), .rdlo_out(a6_wr[56]));
			radix2 #(.width(width)) rd_st5_41  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[41]), .rdlo_in(a5_wr[57]),  .coef_in(coef[288]), .rdup_out(a6_wr[41]), .rdlo_out(a6_wr[57]));
			radix2 #(.width(width)) rd_st5_42  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[42]), .rdlo_in(a5_wr[58]),  .coef_in(coef[320]), .rdup_out(a6_wr[42]), .rdlo_out(a6_wr[58]));
			radix2 #(.width(width)) rd_st5_43  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[43]), .rdlo_in(a5_wr[59]),  .coef_in(coef[352]), .rdup_out(a6_wr[43]), .rdlo_out(a6_wr[59]));
			radix2 #(.width(width)) rd_st5_44  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[44]), .rdlo_in(a5_wr[60]),  .coef_in(coef[384]), .rdup_out(a6_wr[44]), .rdlo_out(a6_wr[60]));
			radix2 #(.width(width)) rd_st5_45  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[45]), .rdlo_in(a5_wr[61]),  .coef_in(coef[416]), .rdup_out(a6_wr[45]), .rdlo_out(a6_wr[61]));
			radix2 #(.width(width)) rd_st5_46  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[46]), .rdlo_in(a5_wr[62]),  .coef_in(coef[448]), .rdup_out(a6_wr[46]), .rdlo_out(a6_wr[62]));
			radix2 #(.width(width)) rd_st5_47  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[47]), .rdlo_in(a5_wr[63]),  .coef_in(coef[480]), .rdup_out(a6_wr[47]), .rdlo_out(a6_wr[63]));
			radix2 #(.width(width)) rd_st5_64  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[64]), .rdlo_in(a5_wr[80]),  .coef_in(coef[0]), .rdup_out(a6_wr[64]), .rdlo_out(a6_wr[80]));
			radix2 #(.width(width)) rd_st5_65  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[65]), .rdlo_in(a5_wr[81]),  .coef_in(coef[32]), .rdup_out(a6_wr[65]), .rdlo_out(a6_wr[81]));
			radix2 #(.width(width)) rd_st5_66  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[66]), .rdlo_in(a5_wr[82]),  .coef_in(coef[64]), .rdup_out(a6_wr[66]), .rdlo_out(a6_wr[82]));
			radix2 #(.width(width)) rd_st5_67  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[67]), .rdlo_in(a5_wr[83]),  .coef_in(coef[96]), .rdup_out(a6_wr[67]), .rdlo_out(a6_wr[83]));
			radix2 #(.width(width)) rd_st5_68  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[68]), .rdlo_in(a5_wr[84]),  .coef_in(coef[128]), .rdup_out(a6_wr[68]), .rdlo_out(a6_wr[84]));
			radix2 #(.width(width)) rd_st5_69  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[69]), .rdlo_in(a5_wr[85]),  .coef_in(coef[160]), .rdup_out(a6_wr[69]), .rdlo_out(a6_wr[85]));
			radix2 #(.width(width)) rd_st5_70  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[70]), .rdlo_in(a5_wr[86]),  .coef_in(coef[192]), .rdup_out(a6_wr[70]), .rdlo_out(a6_wr[86]));
			radix2 #(.width(width)) rd_st5_71  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[71]), .rdlo_in(a5_wr[87]),  .coef_in(coef[224]), .rdup_out(a6_wr[71]), .rdlo_out(a6_wr[87]));
			radix2 #(.width(width)) rd_st5_72  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[72]), .rdlo_in(a5_wr[88]),  .coef_in(coef[256]), .rdup_out(a6_wr[72]), .rdlo_out(a6_wr[88]));
			radix2 #(.width(width)) rd_st5_73  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[73]), .rdlo_in(a5_wr[89]),  .coef_in(coef[288]), .rdup_out(a6_wr[73]), .rdlo_out(a6_wr[89]));
			radix2 #(.width(width)) rd_st5_74  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[74]), .rdlo_in(a5_wr[90]),  .coef_in(coef[320]), .rdup_out(a6_wr[74]), .rdlo_out(a6_wr[90]));
			radix2 #(.width(width)) rd_st5_75  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[75]), .rdlo_in(a5_wr[91]),  .coef_in(coef[352]), .rdup_out(a6_wr[75]), .rdlo_out(a6_wr[91]));
			radix2 #(.width(width)) rd_st5_76  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[76]), .rdlo_in(a5_wr[92]),  .coef_in(coef[384]), .rdup_out(a6_wr[76]), .rdlo_out(a6_wr[92]));
			radix2 #(.width(width)) rd_st5_77  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[77]), .rdlo_in(a5_wr[93]),  .coef_in(coef[416]), .rdup_out(a6_wr[77]), .rdlo_out(a6_wr[93]));
			radix2 #(.width(width)) rd_st5_78  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[78]), .rdlo_in(a5_wr[94]),  .coef_in(coef[448]), .rdup_out(a6_wr[78]), .rdlo_out(a6_wr[94]));
			radix2 #(.width(width)) rd_st5_79  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[79]), .rdlo_in(a5_wr[95]),  .coef_in(coef[480]), .rdup_out(a6_wr[79]), .rdlo_out(a6_wr[95]));
			radix2 #(.width(width)) rd_st5_96  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[96]), .rdlo_in(a5_wr[112]),  .coef_in(coef[0]), .rdup_out(a6_wr[96]), .rdlo_out(a6_wr[112]));
			radix2 #(.width(width)) rd_st5_97  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[97]), .rdlo_in(a5_wr[113]),  .coef_in(coef[32]), .rdup_out(a6_wr[97]), .rdlo_out(a6_wr[113]));
			radix2 #(.width(width)) rd_st5_98  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[98]), .rdlo_in(a5_wr[114]),  .coef_in(coef[64]), .rdup_out(a6_wr[98]), .rdlo_out(a6_wr[114]));
			radix2 #(.width(width)) rd_st5_99  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[99]), .rdlo_in(a5_wr[115]),  .coef_in(coef[96]), .rdup_out(a6_wr[99]), .rdlo_out(a6_wr[115]));
			radix2 #(.width(width)) rd_st5_100  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[100]), .rdlo_in(a5_wr[116]),  .coef_in(coef[128]), .rdup_out(a6_wr[100]), .rdlo_out(a6_wr[116]));
			radix2 #(.width(width)) rd_st5_101  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[101]), .rdlo_in(a5_wr[117]),  .coef_in(coef[160]), .rdup_out(a6_wr[101]), .rdlo_out(a6_wr[117]));
			radix2 #(.width(width)) rd_st5_102  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[102]), .rdlo_in(a5_wr[118]),  .coef_in(coef[192]), .rdup_out(a6_wr[102]), .rdlo_out(a6_wr[118]));
			radix2 #(.width(width)) rd_st5_103  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[103]), .rdlo_in(a5_wr[119]),  .coef_in(coef[224]), .rdup_out(a6_wr[103]), .rdlo_out(a6_wr[119]));
			radix2 #(.width(width)) rd_st5_104  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[104]), .rdlo_in(a5_wr[120]),  .coef_in(coef[256]), .rdup_out(a6_wr[104]), .rdlo_out(a6_wr[120]));
			radix2 #(.width(width)) rd_st5_105  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[105]), .rdlo_in(a5_wr[121]),  .coef_in(coef[288]), .rdup_out(a6_wr[105]), .rdlo_out(a6_wr[121]));
			radix2 #(.width(width)) rd_st5_106  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[106]), .rdlo_in(a5_wr[122]),  .coef_in(coef[320]), .rdup_out(a6_wr[106]), .rdlo_out(a6_wr[122]));
			radix2 #(.width(width)) rd_st5_107  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[107]), .rdlo_in(a5_wr[123]),  .coef_in(coef[352]), .rdup_out(a6_wr[107]), .rdlo_out(a6_wr[123]));
			radix2 #(.width(width)) rd_st5_108  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[108]), .rdlo_in(a5_wr[124]),  .coef_in(coef[384]), .rdup_out(a6_wr[108]), .rdlo_out(a6_wr[124]));
			radix2 #(.width(width)) rd_st5_109  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[109]), .rdlo_in(a5_wr[125]),  .coef_in(coef[416]), .rdup_out(a6_wr[109]), .rdlo_out(a6_wr[125]));
			radix2 #(.width(width)) rd_st5_110  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[110]), .rdlo_in(a5_wr[126]),  .coef_in(coef[448]), .rdup_out(a6_wr[110]), .rdlo_out(a6_wr[126]));
			radix2 #(.width(width)) rd_st5_111  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[111]), .rdlo_in(a5_wr[127]),  .coef_in(coef[480]), .rdup_out(a6_wr[111]), .rdlo_out(a6_wr[127]));
			radix2 #(.width(width)) rd_st5_128  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[128]), .rdlo_in(a5_wr[144]),  .coef_in(coef[0]), .rdup_out(a6_wr[128]), .rdlo_out(a6_wr[144]));
			radix2 #(.width(width)) rd_st5_129  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[129]), .rdlo_in(a5_wr[145]),  .coef_in(coef[32]), .rdup_out(a6_wr[129]), .rdlo_out(a6_wr[145]));
			radix2 #(.width(width)) rd_st5_130  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[130]), .rdlo_in(a5_wr[146]),  .coef_in(coef[64]), .rdup_out(a6_wr[130]), .rdlo_out(a6_wr[146]));
			radix2 #(.width(width)) rd_st5_131  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[131]), .rdlo_in(a5_wr[147]),  .coef_in(coef[96]), .rdup_out(a6_wr[131]), .rdlo_out(a6_wr[147]));
			radix2 #(.width(width)) rd_st5_132  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[132]), .rdlo_in(a5_wr[148]),  .coef_in(coef[128]), .rdup_out(a6_wr[132]), .rdlo_out(a6_wr[148]));
			radix2 #(.width(width)) rd_st5_133  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[133]), .rdlo_in(a5_wr[149]),  .coef_in(coef[160]), .rdup_out(a6_wr[133]), .rdlo_out(a6_wr[149]));
			radix2 #(.width(width)) rd_st5_134  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[134]), .rdlo_in(a5_wr[150]),  .coef_in(coef[192]), .rdup_out(a6_wr[134]), .rdlo_out(a6_wr[150]));
			radix2 #(.width(width)) rd_st5_135  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[135]), .rdlo_in(a5_wr[151]),  .coef_in(coef[224]), .rdup_out(a6_wr[135]), .rdlo_out(a6_wr[151]));
			radix2 #(.width(width)) rd_st5_136  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[136]), .rdlo_in(a5_wr[152]),  .coef_in(coef[256]), .rdup_out(a6_wr[136]), .rdlo_out(a6_wr[152]));
			radix2 #(.width(width)) rd_st5_137  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[137]), .rdlo_in(a5_wr[153]),  .coef_in(coef[288]), .rdup_out(a6_wr[137]), .rdlo_out(a6_wr[153]));
			radix2 #(.width(width)) rd_st5_138  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[138]), .rdlo_in(a5_wr[154]),  .coef_in(coef[320]), .rdup_out(a6_wr[138]), .rdlo_out(a6_wr[154]));
			radix2 #(.width(width)) rd_st5_139  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[139]), .rdlo_in(a5_wr[155]),  .coef_in(coef[352]), .rdup_out(a6_wr[139]), .rdlo_out(a6_wr[155]));
			radix2 #(.width(width)) rd_st5_140  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[140]), .rdlo_in(a5_wr[156]),  .coef_in(coef[384]), .rdup_out(a6_wr[140]), .rdlo_out(a6_wr[156]));
			radix2 #(.width(width)) rd_st5_141  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[141]), .rdlo_in(a5_wr[157]),  .coef_in(coef[416]), .rdup_out(a6_wr[141]), .rdlo_out(a6_wr[157]));
			radix2 #(.width(width)) rd_st5_142  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[142]), .rdlo_in(a5_wr[158]),  .coef_in(coef[448]), .rdup_out(a6_wr[142]), .rdlo_out(a6_wr[158]));
			radix2 #(.width(width)) rd_st5_143  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[143]), .rdlo_in(a5_wr[159]),  .coef_in(coef[480]), .rdup_out(a6_wr[143]), .rdlo_out(a6_wr[159]));
			radix2 #(.width(width)) rd_st5_160  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[160]), .rdlo_in(a5_wr[176]),  .coef_in(coef[0]), .rdup_out(a6_wr[160]), .rdlo_out(a6_wr[176]));
			radix2 #(.width(width)) rd_st5_161  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[161]), .rdlo_in(a5_wr[177]),  .coef_in(coef[32]), .rdup_out(a6_wr[161]), .rdlo_out(a6_wr[177]));
			radix2 #(.width(width)) rd_st5_162  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[162]), .rdlo_in(a5_wr[178]),  .coef_in(coef[64]), .rdup_out(a6_wr[162]), .rdlo_out(a6_wr[178]));
			radix2 #(.width(width)) rd_st5_163  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[163]), .rdlo_in(a5_wr[179]),  .coef_in(coef[96]), .rdup_out(a6_wr[163]), .rdlo_out(a6_wr[179]));
			radix2 #(.width(width)) rd_st5_164  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[164]), .rdlo_in(a5_wr[180]),  .coef_in(coef[128]), .rdup_out(a6_wr[164]), .rdlo_out(a6_wr[180]));
			radix2 #(.width(width)) rd_st5_165  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[165]), .rdlo_in(a5_wr[181]),  .coef_in(coef[160]), .rdup_out(a6_wr[165]), .rdlo_out(a6_wr[181]));
			radix2 #(.width(width)) rd_st5_166  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[166]), .rdlo_in(a5_wr[182]),  .coef_in(coef[192]), .rdup_out(a6_wr[166]), .rdlo_out(a6_wr[182]));
			radix2 #(.width(width)) rd_st5_167  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[167]), .rdlo_in(a5_wr[183]),  .coef_in(coef[224]), .rdup_out(a6_wr[167]), .rdlo_out(a6_wr[183]));
			radix2 #(.width(width)) rd_st5_168  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[168]), .rdlo_in(a5_wr[184]),  .coef_in(coef[256]), .rdup_out(a6_wr[168]), .rdlo_out(a6_wr[184]));
			radix2 #(.width(width)) rd_st5_169  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[169]), .rdlo_in(a5_wr[185]),  .coef_in(coef[288]), .rdup_out(a6_wr[169]), .rdlo_out(a6_wr[185]));
			radix2 #(.width(width)) rd_st5_170  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[170]), .rdlo_in(a5_wr[186]),  .coef_in(coef[320]), .rdup_out(a6_wr[170]), .rdlo_out(a6_wr[186]));
			radix2 #(.width(width)) rd_st5_171  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[171]), .rdlo_in(a5_wr[187]),  .coef_in(coef[352]), .rdup_out(a6_wr[171]), .rdlo_out(a6_wr[187]));
			radix2 #(.width(width)) rd_st5_172  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[172]), .rdlo_in(a5_wr[188]),  .coef_in(coef[384]), .rdup_out(a6_wr[172]), .rdlo_out(a6_wr[188]));
			radix2 #(.width(width)) rd_st5_173  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[173]), .rdlo_in(a5_wr[189]),  .coef_in(coef[416]), .rdup_out(a6_wr[173]), .rdlo_out(a6_wr[189]));
			radix2 #(.width(width)) rd_st5_174  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[174]), .rdlo_in(a5_wr[190]),  .coef_in(coef[448]), .rdup_out(a6_wr[174]), .rdlo_out(a6_wr[190]));
			radix2 #(.width(width)) rd_st5_175  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[175]), .rdlo_in(a5_wr[191]),  .coef_in(coef[480]), .rdup_out(a6_wr[175]), .rdlo_out(a6_wr[191]));
			radix2 #(.width(width)) rd_st5_192  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[192]), .rdlo_in(a5_wr[208]),  .coef_in(coef[0]), .rdup_out(a6_wr[192]), .rdlo_out(a6_wr[208]));
			radix2 #(.width(width)) rd_st5_193  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[193]), .rdlo_in(a5_wr[209]),  .coef_in(coef[32]), .rdup_out(a6_wr[193]), .rdlo_out(a6_wr[209]));
			radix2 #(.width(width)) rd_st5_194  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[194]), .rdlo_in(a5_wr[210]),  .coef_in(coef[64]), .rdup_out(a6_wr[194]), .rdlo_out(a6_wr[210]));
			radix2 #(.width(width)) rd_st5_195  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[195]), .rdlo_in(a5_wr[211]),  .coef_in(coef[96]), .rdup_out(a6_wr[195]), .rdlo_out(a6_wr[211]));
			radix2 #(.width(width)) rd_st5_196  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[196]), .rdlo_in(a5_wr[212]),  .coef_in(coef[128]), .rdup_out(a6_wr[196]), .rdlo_out(a6_wr[212]));
			radix2 #(.width(width)) rd_st5_197  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[197]), .rdlo_in(a5_wr[213]),  .coef_in(coef[160]), .rdup_out(a6_wr[197]), .rdlo_out(a6_wr[213]));
			radix2 #(.width(width)) rd_st5_198  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[198]), .rdlo_in(a5_wr[214]),  .coef_in(coef[192]), .rdup_out(a6_wr[198]), .rdlo_out(a6_wr[214]));
			radix2 #(.width(width)) rd_st5_199  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[199]), .rdlo_in(a5_wr[215]),  .coef_in(coef[224]), .rdup_out(a6_wr[199]), .rdlo_out(a6_wr[215]));
			radix2 #(.width(width)) rd_st5_200  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[200]), .rdlo_in(a5_wr[216]),  .coef_in(coef[256]), .rdup_out(a6_wr[200]), .rdlo_out(a6_wr[216]));
			radix2 #(.width(width)) rd_st5_201  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[201]), .rdlo_in(a5_wr[217]),  .coef_in(coef[288]), .rdup_out(a6_wr[201]), .rdlo_out(a6_wr[217]));
			radix2 #(.width(width)) rd_st5_202  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[202]), .rdlo_in(a5_wr[218]),  .coef_in(coef[320]), .rdup_out(a6_wr[202]), .rdlo_out(a6_wr[218]));
			radix2 #(.width(width)) rd_st5_203  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[203]), .rdlo_in(a5_wr[219]),  .coef_in(coef[352]), .rdup_out(a6_wr[203]), .rdlo_out(a6_wr[219]));
			radix2 #(.width(width)) rd_st5_204  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[204]), .rdlo_in(a5_wr[220]),  .coef_in(coef[384]), .rdup_out(a6_wr[204]), .rdlo_out(a6_wr[220]));
			radix2 #(.width(width)) rd_st5_205  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[205]), .rdlo_in(a5_wr[221]),  .coef_in(coef[416]), .rdup_out(a6_wr[205]), .rdlo_out(a6_wr[221]));
			radix2 #(.width(width)) rd_st5_206  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[206]), .rdlo_in(a5_wr[222]),  .coef_in(coef[448]), .rdup_out(a6_wr[206]), .rdlo_out(a6_wr[222]));
			radix2 #(.width(width)) rd_st5_207  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[207]), .rdlo_in(a5_wr[223]),  .coef_in(coef[480]), .rdup_out(a6_wr[207]), .rdlo_out(a6_wr[223]));
			radix2 #(.width(width)) rd_st5_224  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[224]), .rdlo_in(a5_wr[240]),  .coef_in(coef[0]), .rdup_out(a6_wr[224]), .rdlo_out(a6_wr[240]));
			radix2 #(.width(width)) rd_st5_225  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[225]), .rdlo_in(a5_wr[241]),  .coef_in(coef[32]), .rdup_out(a6_wr[225]), .rdlo_out(a6_wr[241]));
			radix2 #(.width(width)) rd_st5_226  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[226]), .rdlo_in(a5_wr[242]),  .coef_in(coef[64]), .rdup_out(a6_wr[226]), .rdlo_out(a6_wr[242]));
			radix2 #(.width(width)) rd_st5_227  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[227]), .rdlo_in(a5_wr[243]),  .coef_in(coef[96]), .rdup_out(a6_wr[227]), .rdlo_out(a6_wr[243]));
			radix2 #(.width(width)) rd_st5_228  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[228]), .rdlo_in(a5_wr[244]),  .coef_in(coef[128]), .rdup_out(a6_wr[228]), .rdlo_out(a6_wr[244]));
			radix2 #(.width(width)) rd_st5_229  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[229]), .rdlo_in(a5_wr[245]),  .coef_in(coef[160]), .rdup_out(a6_wr[229]), .rdlo_out(a6_wr[245]));
			radix2 #(.width(width)) rd_st5_230  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[230]), .rdlo_in(a5_wr[246]),  .coef_in(coef[192]), .rdup_out(a6_wr[230]), .rdlo_out(a6_wr[246]));
			radix2 #(.width(width)) rd_st5_231  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[231]), .rdlo_in(a5_wr[247]),  .coef_in(coef[224]), .rdup_out(a6_wr[231]), .rdlo_out(a6_wr[247]));
			radix2 #(.width(width)) rd_st5_232  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[232]), .rdlo_in(a5_wr[248]),  .coef_in(coef[256]), .rdup_out(a6_wr[232]), .rdlo_out(a6_wr[248]));
			radix2 #(.width(width)) rd_st5_233  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[233]), .rdlo_in(a5_wr[249]),  .coef_in(coef[288]), .rdup_out(a6_wr[233]), .rdlo_out(a6_wr[249]));
			radix2 #(.width(width)) rd_st5_234  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[234]), .rdlo_in(a5_wr[250]),  .coef_in(coef[320]), .rdup_out(a6_wr[234]), .rdlo_out(a6_wr[250]));
			radix2 #(.width(width)) rd_st5_235  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[235]), .rdlo_in(a5_wr[251]),  .coef_in(coef[352]), .rdup_out(a6_wr[235]), .rdlo_out(a6_wr[251]));
			radix2 #(.width(width)) rd_st5_236  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[236]), .rdlo_in(a5_wr[252]),  .coef_in(coef[384]), .rdup_out(a6_wr[236]), .rdlo_out(a6_wr[252]));
			radix2 #(.width(width)) rd_st5_237  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[237]), .rdlo_in(a5_wr[253]),  .coef_in(coef[416]), .rdup_out(a6_wr[237]), .rdlo_out(a6_wr[253]));
			radix2 #(.width(width)) rd_st5_238  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[238]), .rdlo_in(a5_wr[254]),  .coef_in(coef[448]), .rdup_out(a6_wr[238]), .rdlo_out(a6_wr[254]));
			radix2 #(.width(width)) rd_st5_239  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[239]), .rdlo_in(a5_wr[255]),  .coef_in(coef[480]), .rdup_out(a6_wr[239]), .rdlo_out(a6_wr[255]));
			radix2 #(.width(width)) rd_st5_256  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[256]), .rdlo_in(a5_wr[272]),  .coef_in(coef[0]), .rdup_out(a6_wr[256]), .rdlo_out(a6_wr[272]));
			radix2 #(.width(width)) rd_st5_257  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[257]), .rdlo_in(a5_wr[273]),  .coef_in(coef[32]), .rdup_out(a6_wr[257]), .rdlo_out(a6_wr[273]));
			radix2 #(.width(width)) rd_st5_258  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[258]), .rdlo_in(a5_wr[274]),  .coef_in(coef[64]), .rdup_out(a6_wr[258]), .rdlo_out(a6_wr[274]));
			radix2 #(.width(width)) rd_st5_259  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[259]), .rdlo_in(a5_wr[275]),  .coef_in(coef[96]), .rdup_out(a6_wr[259]), .rdlo_out(a6_wr[275]));
			radix2 #(.width(width)) rd_st5_260  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[260]), .rdlo_in(a5_wr[276]),  .coef_in(coef[128]), .rdup_out(a6_wr[260]), .rdlo_out(a6_wr[276]));
			radix2 #(.width(width)) rd_st5_261  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[261]), .rdlo_in(a5_wr[277]),  .coef_in(coef[160]), .rdup_out(a6_wr[261]), .rdlo_out(a6_wr[277]));
			radix2 #(.width(width)) rd_st5_262  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[262]), .rdlo_in(a5_wr[278]),  .coef_in(coef[192]), .rdup_out(a6_wr[262]), .rdlo_out(a6_wr[278]));
			radix2 #(.width(width)) rd_st5_263  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[263]), .rdlo_in(a5_wr[279]),  .coef_in(coef[224]), .rdup_out(a6_wr[263]), .rdlo_out(a6_wr[279]));
			radix2 #(.width(width)) rd_st5_264  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[264]), .rdlo_in(a5_wr[280]),  .coef_in(coef[256]), .rdup_out(a6_wr[264]), .rdlo_out(a6_wr[280]));
			radix2 #(.width(width)) rd_st5_265  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[265]), .rdlo_in(a5_wr[281]),  .coef_in(coef[288]), .rdup_out(a6_wr[265]), .rdlo_out(a6_wr[281]));
			radix2 #(.width(width)) rd_st5_266  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[266]), .rdlo_in(a5_wr[282]),  .coef_in(coef[320]), .rdup_out(a6_wr[266]), .rdlo_out(a6_wr[282]));
			radix2 #(.width(width)) rd_st5_267  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[267]), .rdlo_in(a5_wr[283]),  .coef_in(coef[352]), .rdup_out(a6_wr[267]), .rdlo_out(a6_wr[283]));
			radix2 #(.width(width)) rd_st5_268  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[268]), .rdlo_in(a5_wr[284]),  .coef_in(coef[384]), .rdup_out(a6_wr[268]), .rdlo_out(a6_wr[284]));
			radix2 #(.width(width)) rd_st5_269  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[269]), .rdlo_in(a5_wr[285]),  .coef_in(coef[416]), .rdup_out(a6_wr[269]), .rdlo_out(a6_wr[285]));
			radix2 #(.width(width)) rd_st5_270  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[270]), .rdlo_in(a5_wr[286]),  .coef_in(coef[448]), .rdup_out(a6_wr[270]), .rdlo_out(a6_wr[286]));
			radix2 #(.width(width)) rd_st5_271  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[271]), .rdlo_in(a5_wr[287]),  .coef_in(coef[480]), .rdup_out(a6_wr[271]), .rdlo_out(a6_wr[287]));
			radix2 #(.width(width)) rd_st5_288  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[288]), .rdlo_in(a5_wr[304]),  .coef_in(coef[0]), .rdup_out(a6_wr[288]), .rdlo_out(a6_wr[304]));
			radix2 #(.width(width)) rd_st5_289  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[289]), .rdlo_in(a5_wr[305]),  .coef_in(coef[32]), .rdup_out(a6_wr[289]), .rdlo_out(a6_wr[305]));
			radix2 #(.width(width)) rd_st5_290  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[290]), .rdlo_in(a5_wr[306]),  .coef_in(coef[64]), .rdup_out(a6_wr[290]), .rdlo_out(a6_wr[306]));
			radix2 #(.width(width)) rd_st5_291  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[291]), .rdlo_in(a5_wr[307]),  .coef_in(coef[96]), .rdup_out(a6_wr[291]), .rdlo_out(a6_wr[307]));
			radix2 #(.width(width)) rd_st5_292  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[292]), .rdlo_in(a5_wr[308]),  .coef_in(coef[128]), .rdup_out(a6_wr[292]), .rdlo_out(a6_wr[308]));
			radix2 #(.width(width)) rd_st5_293  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[293]), .rdlo_in(a5_wr[309]),  .coef_in(coef[160]), .rdup_out(a6_wr[293]), .rdlo_out(a6_wr[309]));
			radix2 #(.width(width)) rd_st5_294  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[294]), .rdlo_in(a5_wr[310]),  .coef_in(coef[192]), .rdup_out(a6_wr[294]), .rdlo_out(a6_wr[310]));
			radix2 #(.width(width)) rd_st5_295  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[295]), .rdlo_in(a5_wr[311]),  .coef_in(coef[224]), .rdup_out(a6_wr[295]), .rdlo_out(a6_wr[311]));
			radix2 #(.width(width)) rd_st5_296  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[296]), .rdlo_in(a5_wr[312]),  .coef_in(coef[256]), .rdup_out(a6_wr[296]), .rdlo_out(a6_wr[312]));
			radix2 #(.width(width)) rd_st5_297  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[297]), .rdlo_in(a5_wr[313]),  .coef_in(coef[288]), .rdup_out(a6_wr[297]), .rdlo_out(a6_wr[313]));
			radix2 #(.width(width)) rd_st5_298  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[298]), .rdlo_in(a5_wr[314]),  .coef_in(coef[320]), .rdup_out(a6_wr[298]), .rdlo_out(a6_wr[314]));
			radix2 #(.width(width)) rd_st5_299  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[299]), .rdlo_in(a5_wr[315]),  .coef_in(coef[352]), .rdup_out(a6_wr[299]), .rdlo_out(a6_wr[315]));
			radix2 #(.width(width)) rd_st5_300  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[300]), .rdlo_in(a5_wr[316]),  .coef_in(coef[384]), .rdup_out(a6_wr[300]), .rdlo_out(a6_wr[316]));
			radix2 #(.width(width)) rd_st5_301  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[301]), .rdlo_in(a5_wr[317]),  .coef_in(coef[416]), .rdup_out(a6_wr[301]), .rdlo_out(a6_wr[317]));
			radix2 #(.width(width)) rd_st5_302  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[302]), .rdlo_in(a5_wr[318]),  .coef_in(coef[448]), .rdup_out(a6_wr[302]), .rdlo_out(a6_wr[318]));
			radix2 #(.width(width)) rd_st5_303  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[303]), .rdlo_in(a5_wr[319]),  .coef_in(coef[480]), .rdup_out(a6_wr[303]), .rdlo_out(a6_wr[319]));
			radix2 #(.width(width)) rd_st5_320  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[320]), .rdlo_in(a5_wr[336]),  .coef_in(coef[0]), .rdup_out(a6_wr[320]), .rdlo_out(a6_wr[336]));
			radix2 #(.width(width)) rd_st5_321  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[321]), .rdlo_in(a5_wr[337]),  .coef_in(coef[32]), .rdup_out(a6_wr[321]), .rdlo_out(a6_wr[337]));
			radix2 #(.width(width)) rd_st5_322  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[322]), .rdlo_in(a5_wr[338]),  .coef_in(coef[64]), .rdup_out(a6_wr[322]), .rdlo_out(a6_wr[338]));
			radix2 #(.width(width)) rd_st5_323  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[323]), .rdlo_in(a5_wr[339]),  .coef_in(coef[96]), .rdup_out(a6_wr[323]), .rdlo_out(a6_wr[339]));
			radix2 #(.width(width)) rd_st5_324  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[324]), .rdlo_in(a5_wr[340]),  .coef_in(coef[128]), .rdup_out(a6_wr[324]), .rdlo_out(a6_wr[340]));
			radix2 #(.width(width)) rd_st5_325  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[325]), .rdlo_in(a5_wr[341]),  .coef_in(coef[160]), .rdup_out(a6_wr[325]), .rdlo_out(a6_wr[341]));
			radix2 #(.width(width)) rd_st5_326  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[326]), .rdlo_in(a5_wr[342]),  .coef_in(coef[192]), .rdup_out(a6_wr[326]), .rdlo_out(a6_wr[342]));
			radix2 #(.width(width)) rd_st5_327  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[327]), .rdlo_in(a5_wr[343]),  .coef_in(coef[224]), .rdup_out(a6_wr[327]), .rdlo_out(a6_wr[343]));
			radix2 #(.width(width)) rd_st5_328  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[328]), .rdlo_in(a5_wr[344]),  .coef_in(coef[256]), .rdup_out(a6_wr[328]), .rdlo_out(a6_wr[344]));
			radix2 #(.width(width)) rd_st5_329  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[329]), .rdlo_in(a5_wr[345]),  .coef_in(coef[288]), .rdup_out(a6_wr[329]), .rdlo_out(a6_wr[345]));
			radix2 #(.width(width)) rd_st5_330  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[330]), .rdlo_in(a5_wr[346]),  .coef_in(coef[320]), .rdup_out(a6_wr[330]), .rdlo_out(a6_wr[346]));
			radix2 #(.width(width)) rd_st5_331  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[331]), .rdlo_in(a5_wr[347]),  .coef_in(coef[352]), .rdup_out(a6_wr[331]), .rdlo_out(a6_wr[347]));
			radix2 #(.width(width)) rd_st5_332  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[332]), .rdlo_in(a5_wr[348]),  .coef_in(coef[384]), .rdup_out(a6_wr[332]), .rdlo_out(a6_wr[348]));
			radix2 #(.width(width)) rd_st5_333  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[333]), .rdlo_in(a5_wr[349]),  .coef_in(coef[416]), .rdup_out(a6_wr[333]), .rdlo_out(a6_wr[349]));
			radix2 #(.width(width)) rd_st5_334  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[334]), .rdlo_in(a5_wr[350]),  .coef_in(coef[448]), .rdup_out(a6_wr[334]), .rdlo_out(a6_wr[350]));
			radix2 #(.width(width)) rd_st5_335  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[335]), .rdlo_in(a5_wr[351]),  .coef_in(coef[480]), .rdup_out(a6_wr[335]), .rdlo_out(a6_wr[351]));
			radix2 #(.width(width)) rd_st5_352  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[352]), .rdlo_in(a5_wr[368]),  .coef_in(coef[0]), .rdup_out(a6_wr[352]), .rdlo_out(a6_wr[368]));
			radix2 #(.width(width)) rd_st5_353  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[353]), .rdlo_in(a5_wr[369]),  .coef_in(coef[32]), .rdup_out(a6_wr[353]), .rdlo_out(a6_wr[369]));
			radix2 #(.width(width)) rd_st5_354  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[354]), .rdlo_in(a5_wr[370]),  .coef_in(coef[64]), .rdup_out(a6_wr[354]), .rdlo_out(a6_wr[370]));
			radix2 #(.width(width)) rd_st5_355  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[355]), .rdlo_in(a5_wr[371]),  .coef_in(coef[96]), .rdup_out(a6_wr[355]), .rdlo_out(a6_wr[371]));
			radix2 #(.width(width)) rd_st5_356  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[356]), .rdlo_in(a5_wr[372]),  .coef_in(coef[128]), .rdup_out(a6_wr[356]), .rdlo_out(a6_wr[372]));
			radix2 #(.width(width)) rd_st5_357  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[357]), .rdlo_in(a5_wr[373]),  .coef_in(coef[160]), .rdup_out(a6_wr[357]), .rdlo_out(a6_wr[373]));
			radix2 #(.width(width)) rd_st5_358  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[358]), .rdlo_in(a5_wr[374]),  .coef_in(coef[192]), .rdup_out(a6_wr[358]), .rdlo_out(a6_wr[374]));
			radix2 #(.width(width)) rd_st5_359  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[359]), .rdlo_in(a5_wr[375]),  .coef_in(coef[224]), .rdup_out(a6_wr[359]), .rdlo_out(a6_wr[375]));
			radix2 #(.width(width)) rd_st5_360  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[360]), .rdlo_in(a5_wr[376]),  .coef_in(coef[256]), .rdup_out(a6_wr[360]), .rdlo_out(a6_wr[376]));
			radix2 #(.width(width)) rd_st5_361  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[361]), .rdlo_in(a5_wr[377]),  .coef_in(coef[288]), .rdup_out(a6_wr[361]), .rdlo_out(a6_wr[377]));
			radix2 #(.width(width)) rd_st5_362  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[362]), .rdlo_in(a5_wr[378]),  .coef_in(coef[320]), .rdup_out(a6_wr[362]), .rdlo_out(a6_wr[378]));
			radix2 #(.width(width)) rd_st5_363  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[363]), .rdlo_in(a5_wr[379]),  .coef_in(coef[352]), .rdup_out(a6_wr[363]), .rdlo_out(a6_wr[379]));
			radix2 #(.width(width)) rd_st5_364  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[364]), .rdlo_in(a5_wr[380]),  .coef_in(coef[384]), .rdup_out(a6_wr[364]), .rdlo_out(a6_wr[380]));
			radix2 #(.width(width)) rd_st5_365  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[365]), .rdlo_in(a5_wr[381]),  .coef_in(coef[416]), .rdup_out(a6_wr[365]), .rdlo_out(a6_wr[381]));
			radix2 #(.width(width)) rd_st5_366  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[366]), .rdlo_in(a5_wr[382]),  .coef_in(coef[448]), .rdup_out(a6_wr[366]), .rdlo_out(a6_wr[382]));
			radix2 #(.width(width)) rd_st5_367  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[367]), .rdlo_in(a5_wr[383]),  .coef_in(coef[480]), .rdup_out(a6_wr[367]), .rdlo_out(a6_wr[383]));
			radix2 #(.width(width)) rd_st5_384  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[384]), .rdlo_in(a5_wr[400]),  .coef_in(coef[0]), .rdup_out(a6_wr[384]), .rdlo_out(a6_wr[400]));
			radix2 #(.width(width)) rd_st5_385  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[385]), .rdlo_in(a5_wr[401]),  .coef_in(coef[32]), .rdup_out(a6_wr[385]), .rdlo_out(a6_wr[401]));
			radix2 #(.width(width)) rd_st5_386  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[386]), .rdlo_in(a5_wr[402]),  .coef_in(coef[64]), .rdup_out(a6_wr[386]), .rdlo_out(a6_wr[402]));
			radix2 #(.width(width)) rd_st5_387  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[387]), .rdlo_in(a5_wr[403]),  .coef_in(coef[96]), .rdup_out(a6_wr[387]), .rdlo_out(a6_wr[403]));
			radix2 #(.width(width)) rd_st5_388  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[388]), .rdlo_in(a5_wr[404]),  .coef_in(coef[128]), .rdup_out(a6_wr[388]), .rdlo_out(a6_wr[404]));
			radix2 #(.width(width)) rd_st5_389  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[389]), .rdlo_in(a5_wr[405]),  .coef_in(coef[160]), .rdup_out(a6_wr[389]), .rdlo_out(a6_wr[405]));
			radix2 #(.width(width)) rd_st5_390  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[390]), .rdlo_in(a5_wr[406]),  .coef_in(coef[192]), .rdup_out(a6_wr[390]), .rdlo_out(a6_wr[406]));
			radix2 #(.width(width)) rd_st5_391  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[391]), .rdlo_in(a5_wr[407]),  .coef_in(coef[224]), .rdup_out(a6_wr[391]), .rdlo_out(a6_wr[407]));
			radix2 #(.width(width)) rd_st5_392  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[392]), .rdlo_in(a5_wr[408]),  .coef_in(coef[256]), .rdup_out(a6_wr[392]), .rdlo_out(a6_wr[408]));
			radix2 #(.width(width)) rd_st5_393  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[393]), .rdlo_in(a5_wr[409]),  .coef_in(coef[288]), .rdup_out(a6_wr[393]), .rdlo_out(a6_wr[409]));
			radix2 #(.width(width)) rd_st5_394  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[394]), .rdlo_in(a5_wr[410]),  .coef_in(coef[320]), .rdup_out(a6_wr[394]), .rdlo_out(a6_wr[410]));
			radix2 #(.width(width)) rd_st5_395  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[395]), .rdlo_in(a5_wr[411]),  .coef_in(coef[352]), .rdup_out(a6_wr[395]), .rdlo_out(a6_wr[411]));
			radix2 #(.width(width)) rd_st5_396  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[396]), .rdlo_in(a5_wr[412]),  .coef_in(coef[384]), .rdup_out(a6_wr[396]), .rdlo_out(a6_wr[412]));
			radix2 #(.width(width)) rd_st5_397  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[397]), .rdlo_in(a5_wr[413]),  .coef_in(coef[416]), .rdup_out(a6_wr[397]), .rdlo_out(a6_wr[413]));
			radix2 #(.width(width)) rd_st5_398  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[398]), .rdlo_in(a5_wr[414]),  .coef_in(coef[448]), .rdup_out(a6_wr[398]), .rdlo_out(a6_wr[414]));
			radix2 #(.width(width)) rd_st5_399  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[399]), .rdlo_in(a5_wr[415]),  .coef_in(coef[480]), .rdup_out(a6_wr[399]), .rdlo_out(a6_wr[415]));
			radix2 #(.width(width)) rd_st5_416  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[416]), .rdlo_in(a5_wr[432]),  .coef_in(coef[0]), .rdup_out(a6_wr[416]), .rdlo_out(a6_wr[432]));
			radix2 #(.width(width)) rd_st5_417  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[417]), .rdlo_in(a5_wr[433]),  .coef_in(coef[32]), .rdup_out(a6_wr[417]), .rdlo_out(a6_wr[433]));
			radix2 #(.width(width)) rd_st5_418  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[418]), .rdlo_in(a5_wr[434]),  .coef_in(coef[64]), .rdup_out(a6_wr[418]), .rdlo_out(a6_wr[434]));
			radix2 #(.width(width)) rd_st5_419  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[419]), .rdlo_in(a5_wr[435]),  .coef_in(coef[96]), .rdup_out(a6_wr[419]), .rdlo_out(a6_wr[435]));
			radix2 #(.width(width)) rd_st5_420  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[420]), .rdlo_in(a5_wr[436]),  .coef_in(coef[128]), .rdup_out(a6_wr[420]), .rdlo_out(a6_wr[436]));
			radix2 #(.width(width)) rd_st5_421  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[421]), .rdlo_in(a5_wr[437]),  .coef_in(coef[160]), .rdup_out(a6_wr[421]), .rdlo_out(a6_wr[437]));
			radix2 #(.width(width)) rd_st5_422  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[422]), .rdlo_in(a5_wr[438]),  .coef_in(coef[192]), .rdup_out(a6_wr[422]), .rdlo_out(a6_wr[438]));
			radix2 #(.width(width)) rd_st5_423  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[423]), .rdlo_in(a5_wr[439]),  .coef_in(coef[224]), .rdup_out(a6_wr[423]), .rdlo_out(a6_wr[439]));
			radix2 #(.width(width)) rd_st5_424  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[424]), .rdlo_in(a5_wr[440]),  .coef_in(coef[256]), .rdup_out(a6_wr[424]), .rdlo_out(a6_wr[440]));
			radix2 #(.width(width)) rd_st5_425  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[425]), .rdlo_in(a5_wr[441]),  .coef_in(coef[288]), .rdup_out(a6_wr[425]), .rdlo_out(a6_wr[441]));
			radix2 #(.width(width)) rd_st5_426  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[426]), .rdlo_in(a5_wr[442]),  .coef_in(coef[320]), .rdup_out(a6_wr[426]), .rdlo_out(a6_wr[442]));
			radix2 #(.width(width)) rd_st5_427  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[427]), .rdlo_in(a5_wr[443]),  .coef_in(coef[352]), .rdup_out(a6_wr[427]), .rdlo_out(a6_wr[443]));
			radix2 #(.width(width)) rd_st5_428  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[428]), .rdlo_in(a5_wr[444]),  .coef_in(coef[384]), .rdup_out(a6_wr[428]), .rdlo_out(a6_wr[444]));
			radix2 #(.width(width)) rd_st5_429  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[429]), .rdlo_in(a5_wr[445]),  .coef_in(coef[416]), .rdup_out(a6_wr[429]), .rdlo_out(a6_wr[445]));
			radix2 #(.width(width)) rd_st5_430  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[430]), .rdlo_in(a5_wr[446]),  .coef_in(coef[448]), .rdup_out(a6_wr[430]), .rdlo_out(a6_wr[446]));
			radix2 #(.width(width)) rd_st5_431  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[431]), .rdlo_in(a5_wr[447]),  .coef_in(coef[480]), .rdup_out(a6_wr[431]), .rdlo_out(a6_wr[447]));
			radix2 #(.width(width)) rd_st5_448  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[448]), .rdlo_in(a5_wr[464]),  .coef_in(coef[0]), .rdup_out(a6_wr[448]), .rdlo_out(a6_wr[464]));
			radix2 #(.width(width)) rd_st5_449  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[449]), .rdlo_in(a5_wr[465]),  .coef_in(coef[32]), .rdup_out(a6_wr[449]), .rdlo_out(a6_wr[465]));
			radix2 #(.width(width)) rd_st5_450  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[450]), .rdlo_in(a5_wr[466]),  .coef_in(coef[64]), .rdup_out(a6_wr[450]), .rdlo_out(a6_wr[466]));
			radix2 #(.width(width)) rd_st5_451  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[451]), .rdlo_in(a5_wr[467]),  .coef_in(coef[96]), .rdup_out(a6_wr[451]), .rdlo_out(a6_wr[467]));
			radix2 #(.width(width)) rd_st5_452  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[452]), .rdlo_in(a5_wr[468]),  .coef_in(coef[128]), .rdup_out(a6_wr[452]), .rdlo_out(a6_wr[468]));
			radix2 #(.width(width)) rd_st5_453  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[453]), .rdlo_in(a5_wr[469]),  .coef_in(coef[160]), .rdup_out(a6_wr[453]), .rdlo_out(a6_wr[469]));
			radix2 #(.width(width)) rd_st5_454  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[454]), .rdlo_in(a5_wr[470]),  .coef_in(coef[192]), .rdup_out(a6_wr[454]), .rdlo_out(a6_wr[470]));
			radix2 #(.width(width)) rd_st5_455  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[455]), .rdlo_in(a5_wr[471]),  .coef_in(coef[224]), .rdup_out(a6_wr[455]), .rdlo_out(a6_wr[471]));
			radix2 #(.width(width)) rd_st5_456  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[456]), .rdlo_in(a5_wr[472]),  .coef_in(coef[256]), .rdup_out(a6_wr[456]), .rdlo_out(a6_wr[472]));
			radix2 #(.width(width)) rd_st5_457  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[457]), .rdlo_in(a5_wr[473]),  .coef_in(coef[288]), .rdup_out(a6_wr[457]), .rdlo_out(a6_wr[473]));
			radix2 #(.width(width)) rd_st5_458  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[458]), .rdlo_in(a5_wr[474]),  .coef_in(coef[320]), .rdup_out(a6_wr[458]), .rdlo_out(a6_wr[474]));
			radix2 #(.width(width)) rd_st5_459  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[459]), .rdlo_in(a5_wr[475]),  .coef_in(coef[352]), .rdup_out(a6_wr[459]), .rdlo_out(a6_wr[475]));
			radix2 #(.width(width)) rd_st5_460  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[460]), .rdlo_in(a5_wr[476]),  .coef_in(coef[384]), .rdup_out(a6_wr[460]), .rdlo_out(a6_wr[476]));
			radix2 #(.width(width)) rd_st5_461  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[461]), .rdlo_in(a5_wr[477]),  .coef_in(coef[416]), .rdup_out(a6_wr[461]), .rdlo_out(a6_wr[477]));
			radix2 #(.width(width)) rd_st5_462  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[462]), .rdlo_in(a5_wr[478]),  .coef_in(coef[448]), .rdup_out(a6_wr[462]), .rdlo_out(a6_wr[478]));
			radix2 #(.width(width)) rd_st5_463  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[463]), .rdlo_in(a5_wr[479]),  .coef_in(coef[480]), .rdup_out(a6_wr[463]), .rdlo_out(a6_wr[479]));
			radix2 #(.width(width)) rd_st5_480  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[480]), .rdlo_in(a5_wr[496]),  .coef_in(coef[0]), .rdup_out(a6_wr[480]), .rdlo_out(a6_wr[496]));
			radix2 #(.width(width)) rd_st5_481  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[481]), .rdlo_in(a5_wr[497]),  .coef_in(coef[32]), .rdup_out(a6_wr[481]), .rdlo_out(a6_wr[497]));
			radix2 #(.width(width)) rd_st5_482  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[482]), .rdlo_in(a5_wr[498]),  .coef_in(coef[64]), .rdup_out(a6_wr[482]), .rdlo_out(a6_wr[498]));
			radix2 #(.width(width)) rd_st5_483  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[483]), .rdlo_in(a5_wr[499]),  .coef_in(coef[96]), .rdup_out(a6_wr[483]), .rdlo_out(a6_wr[499]));
			radix2 #(.width(width)) rd_st5_484  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[484]), .rdlo_in(a5_wr[500]),  .coef_in(coef[128]), .rdup_out(a6_wr[484]), .rdlo_out(a6_wr[500]));
			radix2 #(.width(width)) rd_st5_485  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[485]), .rdlo_in(a5_wr[501]),  .coef_in(coef[160]), .rdup_out(a6_wr[485]), .rdlo_out(a6_wr[501]));
			radix2 #(.width(width)) rd_st5_486  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[486]), .rdlo_in(a5_wr[502]),  .coef_in(coef[192]), .rdup_out(a6_wr[486]), .rdlo_out(a6_wr[502]));
			radix2 #(.width(width)) rd_st5_487  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[487]), .rdlo_in(a5_wr[503]),  .coef_in(coef[224]), .rdup_out(a6_wr[487]), .rdlo_out(a6_wr[503]));
			radix2 #(.width(width)) rd_st5_488  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[488]), .rdlo_in(a5_wr[504]),  .coef_in(coef[256]), .rdup_out(a6_wr[488]), .rdlo_out(a6_wr[504]));
			radix2 #(.width(width)) rd_st5_489  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[489]), .rdlo_in(a5_wr[505]),  .coef_in(coef[288]), .rdup_out(a6_wr[489]), .rdlo_out(a6_wr[505]));
			radix2 #(.width(width)) rd_st5_490  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[490]), .rdlo_in(a5_wr[506]),  .coef_in(coef[320]), .rdup_out(a6_wr[490]), .rdlo_out(a6_wr[506]));
			radix2 #(.width(width)) rd_st5_491  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[491]), .rdlo_in(a5_wr[507]),  .coef_in(coef[352]), .rdup_out(a6_wr[491]), .rdlo_out(a6_wr[507]));
			radix2 #(.width(width)) rd_st5_492  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[492]), .rdlo_in(a5_wr[508]),  .coef_in(coef[384]), .rdup_out(a6_wr[492]), .rdlo_out(a6_wr[508]));
			radix2 #(.width(width)) rd_st5_493  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[493]), .rdlo_in(a5_wr[509]),  .coef_in(coef[416]), .rdup_out(a6_wr[493]), .rdlo_out(a6_wr[509]));
			radix2 #(.width(width)) rd_st5_494  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[494]), .rdlo_in(a5_wr[510]),  .coef_in(coef[448]), .rdup_out(a6_wr[494]), .rdlo_out(a6_wr[510]));
			radix2 #(.width(width)) rd_st5_495  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[495]), .rdlo_in(a5_wr[511]),  .coef_in(coef[480]), .rdup_out(a6_wr[495]), .rdlo_out(a6_wr[511]));
			radix2 #(.width(width)) rd_st5_512  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[512]), .rdlo_in(a5_wr[528]),  .coef_in(coef[0]), .rdup_out(a6_wr[512]), .rdlo_out(a6_wr[528]));
			radix2 #(.width(width)) rd_st5_513  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[513]), .rdlo_in(a5_wr[529]),  .coef_in(coef[32]), .rdup_out(a6_wr[513]), .rdlo_out(a6_wr[529]));
			radix2 #(.width(width)) rd_st5_514  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[514]), .rdlo_in(a5_wr[530]),  .coef_in(coef[64]), .rdup_out(a6_wr[514]), .rdlo_out(a6_wr[530]));
			radix2 #(.width(width)) rd_st5_515  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[515]), .rdlo_in(a5_wr[531]),  .coef_in(coef[96]), .rdup_out(a6_wr[515]), .rdlo_out(a6_wr[531]));
			radix2 #(.width(width)) rd_st5_516  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[516]), .rdlo_in(a5_wr[532]),  .coef_in(coef[128]), .rdup_out(a6_wr[516]), .rdlo_out(a6_wr[532]));
			radix2 #(.width(width)) rd_st5_517  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[517]), .rdlo_in(a5_wr[533]),  .coef_in(coef[160]), .rdup_out(a6_wr[517]), .rdlo_out(a6_wr[533]));
			radix2 #(.width(width)) rd_st5_518  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[518]), .rdlo_in(a5_wr[534]),  .coef_in(coef[192]), .rdup_out(a6_wr[518]), .rdlo_out(a6_wr[534]));
			radix2 #(.width(width)) rd_st5_519  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[519]), .rdlo_in(a5_wr[535]),  .coef_in(coef[224]), .rdup_out(a6_wr[519]), .rdlo_out(a6_wr[535]));
			radix2 #(.width(width)) rd_st5_520  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[520]), .rdlo_in(a5_wr[536]),  .coef_in(coef[256]), .rdup_out(a6_wr[520]), .rdlo_out(a6_wr[536]));
			radix2 #(.width(width)) rd_st5_521  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[521]), .rdlo_in(a5_wr[537]),  .coef_in(coef[288]), .rdup_out(a6_wr[521]), .rdlo_out(a6_wr[537]));
			radix2 #(.width(width)) rd_st5_522  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[522]), .rdlo_in(a5_wr[538]),  .coef_in(coef[320]), .rdup_out(a6_wr[522]), .rdlo_out(a6_wr[538]));
			radix2 #(.width(width)) rd_st5_523  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[523]), .rdlo_in(a5_wr[539]),  .coef_in(coef[352]), .rdup_out(a6_wr[523]), .rdlo_out(a6_wr[539]));
			radix2 #(.width(width)) rd_st5_524  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[524]), .rdlo_in(a5_wr[540]),  .coef_in(coef[384]), .rdup_out(a6_wr[524]), .rdlo_out(a6_wr[540]));
			radix2 #(.width(width)) rd_st5_525  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[525]), .rdlo_in(a5_wr[541]),  .coef_in(coef[416]), .rdup_out(a6_wr[525]), .rdlo_out(a6_wr[541]));
			radix2 #(.width(width)) rd_st5_526  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[526]), .rdlo_in(a5_wr[542]),  .coef_in(coef[448]), .rdup_out(a6_wr[526]), .rdlo_out(a6_wr[542]));
			radix2 #(.width(width)) rd_st5_527  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[527]), .rdlo_in(a5_wr[543]),  .coef_in(coef[480]), .rdup_out(a6_wr[527]), .rdlo_out(a6_wr[543]));
			radix2 #(.width(width)) rd_st5_544  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[544]), .rdlo_in(a5_wr[560]),  .coef_in(coef[0]), .rdup_out(a6_wr[544]), .rdlo_out(a6_wr[560]));
			radix2 #(.width(width)) rd_st5_545  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[545]), .rdlo_in(a5_wr[561]),  .coef_in(coef[32]), .rdup_out(a6_wr[545]), .rdlo_out(a6_wr[561]));
			radix2 #(.width(width)) rd_st5_546  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[546]), .rdlo_in(a5_wr[562]),  .coef_in(coef[64]), .rdup_out(a6_wr[546]), .rdlo_out(a6_wr[562]));
			radix2 #(.width(width)) rd_st5_547  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[547]), .rdlo_in(a5_wr[563]),  .coef_in(coef[96]), .rdup_out(a6_wr[547]), .rdlo_out(a6_wr[563]));
			radix2 #(.width(width)) rd_st5_548  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[548]), .rdlo_in(a5_wr[564]),  .coef_in(coef[128]), .rdup_out(a6_wr[548]), .rdlo_out(a6_wr[564]));
			radix2 #(.width(width)) rd_st5_549  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[549]), .rdlo_in(a5_wr[565]),  .coef_in(coef[160]), .rdup_out(a6_wr[549]), .rdlo_out(a6_wr[565]));
			radix2 #(.width(width)) rd_st5_550  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[550]), .rdlo_in(a5_wr[566]),  .coef_in(coef[192]), .rdup_out(a6_wr[550]), .rdlo_out(a6_wr[566]));
			radix2 #(.width(width)) rd_st5_551  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[551]), .rdlo_in(a5_wr[567]),  .coef_in(coef[224]), .rdup_out(a6_wr[551]), .rdlo_out(a6_wr[567]));
			radix2 #(.width(width)) rd_st5_552  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[552]), .rdlo_in(a5_wr[568]),  .coef_in(coef[256]), .rdup_out(a6_wr[552]), .rdlo_out(a6_wr[568]));
			radix2 #(.width(width)) rd_st5_553  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[553]), .rdlo_in(a5_wr[569]),  .coef_in(coef[288]), .rdup_out(a6_wr[553]), .rdlo_out(a6_wr[569]));
			radix2 #(.width(width)) rd_st5_554  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[554]), .rdlo_in(a5_wr[570]),  .coef_in(coef[320]), .rdup_out(a6_wr[554]), .rdlo_out(a6_wr[570]));
			radix2 #(.width(width)) rd_st5_555  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[555]), .rdlo_in(a5_wr[571]),  .coef_in(coef[352]), .rdup_out(a6_wr[555]), .rdlo_out(a6_wr[571]));
			radix2 #(.width(width)) rd_st5_556  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[556]), .rdlo_in(a5_wr[572]),  .coef_in(coef[384]), .rdup_out(a6_wr[556]), .rdlo_out(a6_wr[572]));
			radix2 #(.width(width)) rd_st5_557  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[557]), .rdlo_in(a5_wr[573]),  .coef_in(coef[416]), .rdup_out(a6_wr[557]), .rdlo_out(a6_wr[573]));
			radix2 #(.width(width)) rd_st5_558  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[558]), .rdlo_in(a5_wr[574]),  .coef_in(coef[448]), .rdup_out(a6_wr[558]), .rdlo_out(a6_wr[574]));
			radix2 #(.width(width)) rd_st5_559  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[559]), .rdlo_in(a5_wr[575]),  .coef_in(coef[480]), .rdup_out(a6_wr[559]), .rdlo_out(a6_wr[575]));
			radix2 #(.width(width)) rd_st5_576  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[576]), .rdlo_in(a5_wr[592]),  .coef_in(coef[0]), .rdup_out(a6_wr[576]), .rdlo_out(a6_wr[592]));
			radix2 #(.width(width)) rd_st5_577  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[577]), .rdlo_in(a5_wr[593]),  .coef_in(coef[32]), .rdup_out(a6_wr[577]), .rdlo_out(a6_wr[593]));
			radix2 #(.width(width)) rd_st5_578  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[578]), .rdlo_in(a5_wr[594]),  .coef_in(coef[64]), .rdup_out(a6_wr[578]), .rdlo_out(a6_wr[594]));
			radix2 #(.width(width)) rd_st5_579  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[579]), .rdlo_in(a5_wr[595]),  .coef_in(coef[96]), .rdup_out(a6_wr[579]), .rdlo_out(a6_wr[595]));
			radix2 #(.width(width)) rd_st5_580  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[580]), .rdlo_in(a5_wr[596]),  .coef_in(coef[128]), .rdup_out(a6_wr[580]), .rdlo_out(a6_wr[596]));
			radix2 #(.width(width)) rd_st5_581  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[581]), .rdlo_in(a5_wr[597]),  .coef_in(coef[160]), .rdup_out(a6_wr[581]), .rdlo_out(a6_wr[597]));
			radix2 #(.width(width)) rd_st5_582  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[582]), .rdlo_in(a5_wr[598]),  .coef_in(coef[192]), .rdup_out(a6_wr[582]), .rdlo_out(a6_wr[598]));
			radix2 #(.width(width)) rd_st5_583  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[583]), .rdlo_in(a5_wr[599]),  .coef_in(coef[224]), .rdup_out(a6_wr[583]), .rdlo_out(a6_wr[599]));
			radix2 #(.width(width)) rd_st5_584  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[584]), .rdlo_in(a5_wr[600]),  .coef_in(coef[256]), .rdup_out(a6_wr[584]), .rdlo_out(a6_wr[600]));
			radix2 #(.width(width)) rd_st5_585  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[585]), .rdlo_in(a5_wr[601]),  .coef_in(coef[288]), .rdup_out(a6_wr[585]), .rdlo_out(a6_wr[601]));
			radix2 #(.width(width)) rd_st5_586  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[586]), .rdlo_in(a5_wr[602]),  .coef_in(coef[320]), .rdup_out(a6_wr[586]), .rdlo_out(a6_wr[602]));
			radix2 #(.width(width)) rd_st5_587  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[587]), .rdlo_in(a5_wr[603]),  .coef_in(coef[352]), .rdup_out(a6_wr[587]), .rdlo_out(a6_wr[603]));
			radix2 #(.width(width)) rd_st5_588  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[588]), .rdlo_in(a5_wr[604]),  .coef_in(coef[384]), .rdup_out(a6_wr[588]), .rdlo_out(a6_wr[604]));
			radix2 #(.width(width)) rd_st5_589  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[589]), .rdlo_in(a5_wr[605]),  .coef_in(coef[416]), .rdup_out(a6_wr[589]), .rdlo_out(a6_wr[605]));
			radix2 #(.width(width)) rd_st5_590  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[590]), .rdlo_in(a5_wr[606]),  .coef_in(coef[448]), .rdup_out(a6_wr[590]), .rdlo_out(a6_wr[606]));
			radix2 #(.width(width)) rd_st5_591  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[591]), .rdlo_in(a5_wr[607]),  .coef_in(coef[480]), .rdup_out(a6_wr[591]), .rdlo_out(a6_wr[607]));
			radix2 #(.width(width)) rd_st5_608  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[608]), .rdlo_in(a5_wr[624]),  .coef_in(coef[0]), .rdup_out(a6_wr[608]), .rdlo_out(a6_wr[624]));
			radix2 #(.width(width)) rd_st5_609  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[609]), .rdlo_in(a5_wr[625]),  .coef_in(coef[32]), .rdup_out(a6_wr[609]), .rdlo_out(a6_wr[625]));
			radix2 #(.width(width)) rd_st5_610  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[610]), .rdlo_in(a5_wr[626]),  .coef_in(coef[64]), .rdup_out(a6_wr[610]), .rdlo_out(a6_wr[626]));
			radix2 #(.width(width)) rd_st5_611  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[611]), .rdlo_in(a5_wr[627]),  .coef_in(coef[96]), .rdup_out(a6_wr[611]), .rdlo_out(a6_wr[627]));
			radix2 #(.width(width)) rd_st5_612  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[612]), .rdlo_in(a5_wr[628]),  .coef_in(coef[128]), .rdup_out(a6_wr[612]), .rdlo_out(a6_wr[628]));
			radix2 #(.width(width)) rd_st5_613  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[613]), .rdlo_in(a5_wr[629]),  .coef_in(coef[160]), .rdup_out(a6_wr[613]), .rdlo_out(a6_wr[629]));
			radix2 #(.width(width)) rd_st5_614  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[614]), .rdlo_in(a5_wr[630]),  .coef_in(coef[192]), .rdup_out(a6_wr[614]), .rdlo_out(a6_wr[630]));
			radix2 #(.width(width)) rd_st5_615  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[615]), .rdlo_in(a5_wr[631]),  .coef_in(coef[224]), .rdup_out(a6_wr[615]), .rdlo_out(a6_wr[631]));
			radix2 #(.width(width)) rd_st5_616  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[616]), .rdlo_in(a5_wr[632]),  .coef_in(coef[256]), .rdup_out(a6_wr[616]), .rdlo_out(a6_wr[632]));
			radix2 #(.width(width)) rd_st5_617  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[617]), .rdlo_in(a5_wr[633]),  .coef_in(coef[288]), .rdup_out(a6_wr[617]), .rdlo_out(a6_wr[633]));
			radix2 #(.width(width)) rd_st5_618  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[618]), .rdlo_in(a5_wr[634]),  .coef_in(coef[320]), .rdup_out(a6_wr[618]), .rdlo_out(a6_wr[634]));
			radix2 #(.width(width)) rd_st5_619  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[619]), .rdlo_in(a5_wr[635]),  .coef_in(coef[352]), .rdup_out(a6_wr[619]), .rdlo_out(a6_wr[635]));
			radix2 #(.width(width)) rd_st5_620  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[620]), .rdlo_in(a5_wr[636]),  .coef_in(coef[384]), .rdup_out(a6_wr[620]), .rdlo_out(a6_wr[636]));
			radix2 #(.width(width)) rd_st5_621  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[621]), .rdlo_in(a5_wr[637]),  .coef_in(coef[416]), .rdup_out(a6_wr[621]), .rdlo_out(a6_wr[637]));
			radix2 #(.width(width)) rd_st5_622  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[622]), .rdlo_in(a5_wr[638]),  .coef_in(coef[448]), .rdup_out(a6_wr[622]), .rdlo_out(a6_wr[638]));
			radix2 #(.width(width)) rd_st5_623  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[623]), .rdlo_in(a5_wr[639]),  .coef_in(coef[480]), .rdup_out(a6_wr[623]), .rdlo_out(a6_wr[639]));
			radix2 #(.width(width)) rd_st5_640  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[640]), .rdlo_in(a5_wr[656]),  .coef_in(coef[0]), .rdup_out(a6_wr[640]), .rdlo_out(a6_wr[656]));
			radix2 #(.width(width)) rd_st5_641  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[641]), .rdlo_in(a5_wr[657]),  .coef_in(coef[32]), .rdup_out(a6_wr[641]), .rdlo_out(a6_wr[657]));
			radix2 #(.width(width)) rd_st5_642  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[642]), .rdlo_in(a5_wr[658]),  .coef_in(coef[64]), .rdup_out(a6_wr[642]), .rdlo_out(a6_wr[658]));
			radix2 #(.width(width)) rd_st5_643  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[643]), .rdlo_in(a5_wr[659]),  .coef_in(coef[96]), .rdup_out(a6_wr[643]), .rdlo_out(a6_wr[659]));
			radix2 #(.width(width)) rd_st5_644  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[644]), .rdlo_in(a5_wr[660]),  .coef_in(coef[128]), .rdup_out(a6_wr[644]), .rdlo_out(a6_wr[660]));
			radix2 #(.width(width)) rd_st5_645  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[645]), .rdlo_in(a5_wr[661]),  .coef_in(coef[160]), .rdup_out(a6_wr[645]), .rdlo_out(a6_wr[661]));
			radix2 #(.width(width)) rd_st5_646  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[646]), .rdlo_in(a5_wr[662]),  .coef_in(coef[192]), .rdup_out(a6_wr[646]), .rdlo_out(a6_wr[662]));
			radix2 #(.width(width)) rd_st5_647  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[647]), .rdlo_in(a5_wr[663]),  .coef_in(coef[224]), .rdup_out(a6_wr[647]), .rdlo_out(a6_wr[663]));
			radix2 #(.width(width)) rd_st5_648  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[648]), .rdlo_in(a5_wr[664]),  .coef_in(coef[256]), .rdup_out(a6_wr[648]), .rdlo_out(a6_wr[664]));
			radix2 #(.width(width)) rd_st5_649  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[649]), .rdlo_in(a5_wr[665]),  .coef_in(coef[288]), .rdup_out(a6_wr[649]), .rdlo_out(a6_wr[665]));
			radix2 #(.width(width)) rd_st5_650  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[650]), .rdlo_in(a5_wr[666]),  .coef_in(coef[320]), .rdup_out(a6_wr[650]), .rdlo_out(a6_wr[666]));
			radix2 #(.width(width)) rd_st5_651  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[651]), .rdlo_in(a5_wr[667]),  .coef_in(coef[352]), .rdup_out(a6_wr[651]), .rdlo_out(a6_wr[667]));
			radix2 #(.width(width)) rd_st5_652  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[652]), .rdlo_in(a5_wr[668]),  .coef_in(coef[384]), .rdup_out(a6_wr[652]), .rdlo_out(a6_wr[668]));
			radix2 #(.width(width)) rd_st5_653  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[653]), .rdlo_in(a5_wr[669]),  .coef_in(coef[416]), .rdup_out(a6_wr[653]), .rdlo_out(a6_wr[669]));
			radix2 #(.width(width)) rd_st5_654  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[654]), .rdlo_in(a5_wr[670]),  .coef_in(coef[448]), .rdup_out(a6_wr[654]), .rdlo_out(a6_wr[670]));
			radix2 #(.width(width)) rd_st5_655  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[655]), .rdlo_in(a5_wr[671]),  .coef_in(coef[480]), .rdup_out(a6_wr[655]), .rdlo_out(a6_wr[671]));
			radix2 #(.width(width)) rd_st5_672  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[672]), .rdlo_in(a5_wr[688]),  .coef_in(coef[0]), .rdup_out(a6_wr[672]), .rdlo_out(a6_wr[688]));
			radix2 #(.width(width)) rd_st5_673  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[673]), .rdlo_in(a5_wr[689]),  .coef_in(coef[32]), .rdup_out(a6_wr[673]), .rdlo_out(a6_wr[689]));
			radix2 #(.width(width)) rd_st5_674  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[674]), .rdlo_in(a5_wr[690]),  .coef_in(coef[64]), .rdup_out(a6_wr[674]), .rdlo_out(a6_wr[690]));
			radix2 #(.width(width)) rd_st5_675  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[675]), .rdlo_in(a5_wr[691]),  .coef_in(coef[96]), .rdup_out(a6_wr[675]), .rdlo_out(a6_wr[691]));
			radix2 #(.width(width)) rd_st5_676  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[676]), .rdlo_in(a5_wr[692]),  .coef_in(coef[128]), .rdup_out(a6_wr[676]), .rdlo_out(a6_wr[692]));
			radix2 #(.width(width)) rd_st5_677  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[677]), .rdlo_in(a5_wr[693]),  .coef_in(coef[160]), .rdup_out(a6_wr[677]), .rdlo_out(a6_wr[693]));
			radix2 #(.width(width)) rd_st5_678  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[678]), .rdlo_in(a5_wr[694]),  .coef_in(coef[192]), .rdup_out(a6_wr[678]), .rdlo_out(a6_wr[694]));
			radix2 #(.width(width)) rd_st5_679  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[679]), .rdlo_in(a5_wr[695]),  .coef_in(coef[224]), .rdup_out(a6_wr[679]), .rdlo_out(a6_wr[695]));
			radix2 #(.width(width)) rd_st5_680  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[680]), .rdlo_in(a5_wr[696]),  .coef_in(coef[256]), .rdup_out(a6_wr[680]), .rdlo_out(a6_wr[696]));
			radix2 #(.width(width)) rd_st5_681  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[681]), .rdlo_in(a5_wr[697]),  .coef_in(coef[288]), .rdup_out(a6_wr[681]), .rdlo_out(a6_wr[697]));
			radix2 #(.width(width)) rd_st5_682  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[682]), .rdlo_in(a5_wr[698]),  .coef_in(coef[320]), .rdup_out(a6_wr[682]), .rdlo_out(a6_wr[698]));
			radix2 #(.width(width)) rd_st5_683  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[683]), .rdlo_in(a5_wr[699]),  .coef_in(coef[352]), .rdup_out(a6_wr[683]), .rdlo_out(a6_wr[699]));
			radix2 #(.width(width)) rd_st5_684  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[684]), .rdlo_in(a5_wr[700]),  .coef_in(coef[384]), .rdup_out(a6_wr[684]), .rdlo_out(a6_wr[700]));
			radix2 #(.width(width)) rd_st5_685  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[685]), .rdlo_in(a5_wr[701]),  .coef_in(coef[416]), .rdup_out(a6_wr[685]), .rdlo_out(a6_wr[701]));
			radix2 #(.width(width)) rd_st5_686  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[686]), .rdlo_in(a5_wr[702]),  .coef_in(coef[448]), .rdup_out(a6_wr[686]), .rdlo_out(a6_wr[702]));
			radix2 #(.width(width)) rd_st5_687  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[687]), .rdlo_in(a5_wr[703]),  .coef_in(coef[480]), .rdup_out(a6_wr[687]), .rdlo_out(a6_wr[703]));
			radix2 #(.width(width)) rd_st5_704  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[704]), .rdlo_in(a5_wr[720]),  .coef_in(coef[0]), .rdup_out(a6_wr[704]), .rdlo_out(a6_wr[720]));
			radix2 #(.width(width)) rd_st5_705  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[705]), .rdlo_in(a5_wr[721]),  .coef_in(coef[32]), .rdup_out(a6_wr[705]), .rdlo_out(a6_wr[721]));
			radix2 #(.width(width)) rd_st5_706  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[706]), .rdlo_in(a5_wr[722]),  .coef_in(coef[64]), .rdup_out(a6_wr[706]), .rdlo_out(a6_wr[722]));
			radix2 #(.width(width)) rd_st5_707  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[707]), .rdlo_in(a5_wr[723]),  .coef_in(coef[96]), .rdup_out(a6_wr[707]), .rdlo_out(a6_wr[723]));
			radix2 #(.width(width)) rd_st5_708  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[708]), .rdlo_in(a5_wr[724]),  .coef_in(coef[128]), .rdup_out(a6_wr[708]), .rdlo_out(a6_wr[724]));
			radix2 #(.width(width)) rd_st5_709  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[709]), .rdlo_in(a5_wr[725]),  .coef_in(coef[160]), .rdup_out(a6_wr[709]), .rdlo_out(a6_wr[725]));
			radix2 #(.width(width)) rd_st5_710  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[710]), .rdlo_in(a5_wr[726]),  .coef_in(coef[192]), .rdup_out(a6_wr[710]), .rdlo_out(a6_wr[726]));
			radix2 #(.width(width)) rd_st5_711  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[711]), .rdlo_in(a5_wr[727]),  .coef_in(coef[224]), .rdup_out(a6_wr[711]), .rdlo_out(a6_wr[727]));
			radix2 #(.width(width)) rd_st5_712  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[712]), .rdlo_in(a5_wr[728]),  .coef_in(coef[256]), .rdup_out(a6_wr[712]), .rdlo_out(a6_wr[728]));
			radix2 #(.width(width)) rd_st5_713  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[713]), .rdlo_in(a5_wr[729]),  .coef_in(coef[288]), .rdup_out(a6_wr[713]), .rdlo_out(a6_wr[729]));
			radix2 #(.width(width)) rd_st5_714  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[714]), .rdlo_in(a5_wr[730]),  .coef_in(coef[320]), .rdup_out(a6_wr[714]), .rdlo_out(a6_wr[730]));
			radix2 #(.width(width)) rd_st5_715  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[715]), .rdlo_in(a5_wr[731]),  .coef_in(coef[352]), .rdup_out(a6_wr[715]), .rdlo_out(a6_wr[731]));
			radix2 #(.width(width)) rd_st5_716  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[716]), .rdlo_in(a5_wr[732]),  .coef_in(coef[384]), .rdup_out(a6_wr[716]), .rdlo_out(a6_wr[732]));
			radix2 #(.width(width)) rd_st5_717  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[717]), .rdlo_in(a5_wr[733]),  .coef_in(coef[416]), .rdup_out(a6_wr[717]), .rdlo_out(a6_wr[733]));
			radix2 #(.width(width)) rd_st5_718  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[718]), .rdlo_in(a5_wr[734]),  .coef_in(coef[448]), .rdup_out(a6_wr[718]), .rdlo_out(a6_wr[734]));
			radix2 #(.width(width)) rd_st5_719  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[719]), .rdlo_in(a5_wr[735]),  .coef_in(coef[480]), .rdup_out(a6_wr[719]), .rdlo_out(a6_wr[735]));
			radix2 #(.width(width)) rd_st5_736  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[736]), .rdlo_in(a5_wr[752]),  .coef_in(coef[0]), .rdup_out(a6_wr[736]), .rdlo_out(a6_wr[752]));
			radix2 #(.width(width)) rd_st5_737  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[737]), .rdlo_in(a5_wr[753]),  .coef_in(coef[32]), .rdup_out(a6_wr[737]), .rdlo_out(a6_wr[753]));
			radix2 #(.width(width)) rd_st5_738  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[738]), .rdlo_in(a5_wr[754]),  .coef_in(coef[64]), .rdup_out(a6_wr[738]), .rdlo_out(a6_wr[754]));
			radix2 #(.width(width)) rd_st5_739  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[739]), .rdlo_in(a5_wr[755]),  .coef_in(coef[96]), .rdup_out(a6_wr[739]), .rdlo_out(a6_wr[755]));
			radix2 #(.width(width)) rd_st5_740  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[740]), .rdlo_in(a5_wr[756]),  .coef_in(coef[128]), .rdup_out(a6_wr[740]), .rdlo_out(a6_wr[756]));
			radix2 #(.width(width)) rd_st5_741  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[741]), .rdlo_in(a5_wr[757]),  .coef_in(coef[160]), .rdup_out(a6_wr[741]), .rdlo_out(a6_wr[757]));
			radix2 #(.width(width)) rd_st5_742  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[742]), .rdlo_in(a5_wr[758]),  .coef_in(coef[192]), .rdup_out(a6_wr[742]), .rdlo_out(a6_wr[758]));
			radix2 #(.width(width)) rd_st5_743  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[743]), .rdlo_in(a5_wr[759]),  .coef_in(coef[224]), .rdup_out(a6_wr[743]), .rdlo_out(a6_wr[759]));
			radix2 #(.width(width)) rd_st5_744  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[744]), .rdlo_in(a5_wr[760]),  .coef_in(coef[256]), .rdup_out(a6_wr[744]), .rdlo_out(a6_wr[760]));
			radix2 #(.width(width)) rd_st5_745  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[745]), .rdlo_in(a5_wr[761]),  .coef_in(coef[288]), .rdup_out(a6_wr[745]), .rdlo_out(a6_wr[761]));
			radix2 #(.width(width)) rd_st5_746  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[746]), .rdlo_in(a5_wr[762]),  .coef_in(coef[320]), .rdup_out(a6_wr[746]), .rdlo_out(a6_wr[762]));
			radix2 #(.width(width)) rd_st5_747  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[747]), .rdlo_in(a5_wr[763]),  .coef_in(coef[352]), .rdup_out(a6_wr[747]), .rdlo_out(a6_wr[763]));
			radix2 #(.width(width)) rd_st5_748  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[748]), .rdlo_in(a5_wr[764]),  .coef_in(coef[384]), .rdup_out(a6_wr[748]), .rdlo_out(a6_wr[764]));
			radix2 #(.width(width)) rd_st5_749  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[749]), .rdlo_in(a5_wr[765]),  .coef_in(coef[416]), .rdup_out(a6_wr[749]), .rdlo_out(a6_wr[765]));
			radix2 #(.width(width)) rd_st5_750  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[750]), .rdlo_in(a5_wr[766]),  .coef_in(coef[448]), .rdup_out(a6_wr[750]), .rdlo_out(a6_wr[766]));
			radix2 #(.width(width)) rd_st5_751  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[751]), .rdlo_in(a5_wr[767]),  .coef_in(coef[480]), .rdup_out(a6_wr[751]), .rdlo_out(a6_wr[767]));
			radix2 #(.width(width)) rd_st5_768  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[768]), .rdlo_in(a5_wr[784]),  .coef_in(coef[0]), .rdup_out(a6_wr[768]), .rdlo_out(a6_wr[784]));
			radix2 #(.width(width)) rd_st5_769  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[769]), .rdlo_in(a5_wr[785]),  .coef_in(coef[32]), .rdup_out(a6_wr[769]), .rdlo_out(a6_wr[785]));
			radix2 #(.width(width)) rd_st5_770  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[770]), .rdlo_in(a5_wr[786]),  .coef_in(coef[64]), .rdup_out(a6_wr[770]), .rdlo_out(a6_wr[786]));
			radix2 #(.width(width)) rd_st5_771  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[771]), .rdlo_in(a5_wr[787]),  .coef_in(coef[96]), .rdup_out(a6_wr[771]), .rdlo_out(a6_wr[787]));
			radix2 #(.width(width)) rd_st5_772  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[772]), .rdlo_in(a5_wr[788]),  .coef_in(coef[128]), .rdup_out(a6_wr[772]), .rdlo_out(a6_wr[788]));
			radix2 #(.width(width)) rd_st5_773  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[773]), .rdlo_in(a5_wr[789]),  .coef_in(coef[160]), .rdup_out(a6_wr[773]), .rdlo_out(a6_wr[789]));
			radix2 #(.width(width)) rd_st5_774  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[774]), .rdlo_in(a5_wr[790]),  .coef_in(coef[192]), .rdup_out(a6_wr[774]), .rdlo_out(a6_wr[790]));
			radix2 #(.width(width)) rd_st5_775  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[775]), .rdlo_in(a5_wr[791]),  .coef_in(coef[224]), .rdup_out(a6_wr[775]), .rdlo_out(a6_wr[791]));
			radix2 #(.width(width)) rd_st5_776  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[776]), .rdlo_in(a5_wr[792]),  .coef_in(coef[256]), .rdup_out(a6_wr[776]), .rdlo_out(a6_wr[792]));
			radix2 #(.width(width)) rd_st5_777  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[777]), .rdlo_in(a5_wr[793]),  .coef_in(coef[288]), .rdup_out(a6_wr[777]), .rdlo_out(a6_wr[793]));
			radix2 #(.width(width)) rd_st5_778  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[778]), .rdlo_in(a5_wr[794]),  .coef_in(coef[320]), .rdup_out(a6_wr[778]), .rdlo_out(a6_wr[794]));
			radix2 #(.width(width)) rd_st5_779  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[779]), .rdlo_in(a5_wr[795]),  .coef_in(coef[352]), .rdup_out(a6_wr[779]), .rdlo_out(a6_wr[795]));
			radix2 #(.width(width)) rd_st5_780  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[780]), .rdlo_in(a5_wr[796]),  .coef_in(coef[384]), .rdup_out(a6_wr[780]), .rdlo_out(a6_wr[796]));
			radix2 #(.width(width)) rd_st5_781  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[781]), .rdlo_in(a5_wr[797]),  .coef_in(coef[416]), .rdup_out(a6_wr[781]), .rdlo_out(a6_wr[797]));
			radix2 #(.width(width)) rd_st5_782  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[782]), .rdlo_in(a5_wr[798]),  .coef_in(coef[448]), .rdup_out(a6_wr[782]), .rdlo_out(a6_wr[798]));
			radix2 #(.width(width)) rd_st5_783  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[783]), .rdlo_in(a5_wr[799]),  .coef_in(coef[480]), .rdup_out(a6_wr[783]), .rdlo_out(a6_wr[799]));
			radix2 #(.width(width)) rd_st5_800  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[800]), .rdlo_in(a5_wr[816]),  .coef_in(coef[0]), .rdup_out(a6_wr[800]), .rdlo_out(a6_wr[816]));
			radix2 #(.width(width)) rd_st5_801  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[801]), .rdlo_in(a5_wr[817]),  .coef_in(coef[32]), .rdup_out(a6_wr[801]), .rdlo_out(a6_wr[817]));
			radix2 #(.width(width)) rd_st5_802  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[802]), .rdlo_in(a5_wr[818]),  .coef_in(coef[64]), .rdup_out(a6_wr[802]), .rdlo_out(a6_wr[818]));
			radix2 #(.width(width)) rd_st5_803  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[803]), .rdlo_in(a5_wr[819]),  .coef_in(coef[96]), .rdup_out(a6_wr[803]), .rdlo_out(a6_wr[819]));
			radix2 #(.width(width)) rd_st5_804  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[804]), .rdlo_in(a5_wr[820]),  .coef_in(coef[128]), .rdup_out(a6_wr[804]), .rdlo_out(a6_wr[820]));
			radix2 #(.width(width)) rd_st5_805  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[805]), .rdlo_in(a5_wr[821]),  .coef_in(coef[160]), .rdup_out(a6_wr[805]), .rdlo_out(a6_wr[821]));
			radix2 #(.width(width)) rd_st5_806  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[806]), .rdlo_in(a5_wr[822]),  .coef_in(coef[192]), .rdup_out(a6_wr[806]), .rdlo_out(a6_wr[822]));
			radix2 #(.width(width)) rd_st5_807  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[807]), .rdlo_in(a5_wr[823]),  .coef_in(coef[224]), .rdup_out(a6_wr[807]), .rdlo_out(a6_wr[823]));
			radix2 #(.width(width)) rd_st5_808  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[808]), .rdlo_in(a5_wr[824]),  .coef_in(coef[256]), .rdup_out(a6_wr[808]), .rdlo_out(a6_wr[824]));
			radix2 #(.width(width)) rd_st5_809  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[809]), .rdlo_in(a5_wr[825]),  .coef_in(coef[288]), .rdup_out(a6_wr[809]), .rdlo_out(a6_wr[825]));
			radix2 #(.width(width)) rd_st5_810  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[810]), .rdlo_in(a5_wr[826]),  .coef_in(coef[320]), .rdup_out(a6_wr[810]), .rdlo_out(a6_wr[826]));
			radix2 #(.width(width)) rd_st5_811  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[811]), .rdlo_in(a5_wr[827]),  .coef_in(coef[352]), .rdup_out(a6_wr[811]), .rdlo_out(a6_wr[827]));
			radix2 #(.width(width)) rd_st5_812  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[812]), .rdlo_in(a5_wr[828]),  .coef_in(coef[384]), .rdup_out(a6_wr[812]), .rdlo_out(a6_wr[828]));
			radix2 #(.width(width)) rd_st5_813  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[813]), .rdlo_in(a5_wr[829]),  .coef_in(coef[416]), .rdup_out(a6_wr[813]), .rdlo_out(a6_wr[829]));
			radix2 #(.width(width)) rd_st5_814  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[814]), .rdlo_in(a5_wr[830]),  .coef_in(coef[448]), .rdup_out(a6_wr[814]), .rdlo_out(a6_wr[830]));
			radix2 #(.width(width)) rd_st5_815  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[815]), .rdlo_in(a5_wr[831]),  .coef_in(coef[480]), .rdup_out(a6_wr[815]), .rdlo_out(a6_wr[831]));
			radix2 #(.width(width)) rd_st5_832  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[832]), .rdlo_in(a5_wr[848]),  .coef_in(coef[0]), .rdup_out(a6_wr[832]), .rdlo_out(a6_wr[848]));
			radix2 #(.width(width)) rd_st5_833  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[833]), .rdlo_in(a5_wr[849]),  .coef_in(coef[32]), .rdup_out(a6_wr[833]), .rdlo_out(a6_wr[849]));
			radix2 #(.width(width)) rd_st5_834  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[834]), .rdlo_in(a5_wr[850]),  .coef_in(coef[64]), .rdup_out(a6_wr[834]), .rdlo_out(a6_wr[850]));
			radix2 #(.width(width)) rd_st5_835  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[835]), .rdlo_in(a5_wr[851]),  .coef_in(coef[96]), .rdup_out(a6_wr[835]), .rdlo_out(a6_wr[851]));
			radix2 #(.width(width)) rd_st5_836  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[836]), .rdlo_in(a5_wr[852]),  .coef_in(coef[128]), .rdup_out(a6_wr[836]), .rdlo_out(a6_wr[852]));
			radix2 #(.width(width)) rd_st5_837  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[837]), .rdlo_in(a5_wr[853]),  .coef_in(coef[160]), .rdup_out(a6_wr[837]), .rdlo_out(a6_wr[853]));
			radix2 #(.width(width)) rd_st5_838  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[838]), .rdlo_in(a5_wr[854]),  .coef_in(coef[192]), .rdup_out(a6_wr[838]), .rdlo_out(a6_wr[854]));
			radix2 #(.width(width)) rd_st5_839  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[839]), .rdlo_in(a5_wr[855]),  .coef_in(coef[224]), .rdup_out(a6_wr[839]), .rdlo_out(a6_wr[855]));
			radix2 #(.width(width)) rd_st5_840  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[840]), .rdlo_in(a5_wr[856]),  .coef_in(coef[256]), .rdup_out(a6_wr[840]), .rdlo_out(a6_wr[856]));
			radix2 #(.width(width)) rd_st5_841  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[841]), .rdlo_in(a5_wr[857]),  .coef_in(coef[288]), .rdup_out(a6_wr[841]), .rdlo_out(a6_wr[857]));
			radix2 #(.width(width)) rd_st5_842  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[842]), .rdlo_in(a5_wr[858]),  .coef_in(coef[320]), .rdup_out(a6_wr[842]), .rdlo_out(a6_wr[858]));
			radix2 #(.width(width)) rd_st5_843  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[843]), .rdlo_in(a5_wr[859]),  .coef_in(coef[352]), .rdup_out(a6_wr[843]), .rdlo_out(a6_wr[859]));
			radix2 #(.width(width)) rd_st5_844  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[844]), .rdlo_in(a5_wr[860]),  .coef_in(coef[384]), .rdup_out(a6_wr[844]), .rdlo_out(a6_wr[860]));
			radix2 #(.width(width)) rd_st5_845  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[845]), .rdlo_in(a5_wr[861]),  .coef_in(coef[416]), .rdup_out(a6_wr[845]), .rdlo_out(a6_wr[861]));
			radix2 #(.width(width)) rd_st5_846  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[846]), .rdlo_in(a5_wr[862]),  .coef_in(coef[448]), .rdup_out(a6_wr[846]), .rdlo_out(a6_wr[862]));
			radix2 #(.width(width)) rd_st5_847  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[847]), .rdlo_in(a5_wr[863]),  .coef_in(coef[480]), .rdup_out(a6_wr[847]), .rdlo_out(a6_wr[863]));
			radix2 #(.width(width)) rd_st5_864  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[864]), .rdlo_in(a5_wr[880]),  .coef_in(coef[0]), .rdup_out(a6_wr[864]), .rdlo_out(a6_wr[880]));
			radix2 #(.width(width)) rd_st5_865  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[865]), .rdlo_in(a5_wr[881]),  .coef_in(coef[32]), .rdup_out(a6_wr[865]), .rdlo_out(a6_wr[881]));
			radix2 #(.width(width)) rd_st5_866  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[866]), .rdlo_in(a5_wr[882]),  .coef_in(coef[64]), .rdup_out(a6_wr[866]), .rdlo_out(a6_wr[882]));
			radix2 #(.width(width)) rd_st5_867  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[867]), .rdlo_in(a5_wr[883]),  .coef_in(coef[96]), .rdup_out(a6_wr[867]), .rdlo_out(a6_wr[883]));
			radix2 #(.width(width)) rd_st5_868  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[868]), .rdlo_in(a5_wr[884]),  .coef_in(coef[128]), .rdup_out(a6_wr[868]), .rdlo_out(a6_wr[884]));
			radix2 #(.width(width)) rd_st5_869  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[869]), .rdlo_in(a5_wr[885]),  .coef_in(coef[160]), .rdup_out(a6_wr[869]), .rdlo_out(a6_wr[885]));
			radix2 #(.width(width)) rd_st5_870  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[870]), .rdlo_in(a5_wr[886]),  .coef_in(coef[192]), .rdup_out(a6_wr[870]), .rdlo_out(a6_wr[886]));
			radix2 #(.width(width)) rd_st5_871  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[871]), .rdlo_in(a5_wr[887]),  .coef_in(coef[224]), .rdup_out(a6_wr[871]), .rdlo_out(a6_wr[887]));
			radix2 #(.width(width)) rd_st5_872  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[872]), .rdlo_in(a5_wr[888]),  .coef_in(coef[256]), .rdup_out(a6_wr[872]), .rdlo_out(a6_wr[888]));
			radix2 #(.width(width)) rd_st5_873  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[873]), .rdlo_in(a5_wr[889]),  .coef_in(coef[288]), .rdup_out(a6_wr[873]), .rdlo_out(a6_wr[889]));
			radix2 #(.width(width)) rd_st5_874  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[874]), .rdlo_in(a5_wr[890]),  .coef_in(coef[320]), .rdup_out(a6_wr[874]), .rdlo_out(a6_wr[890]));
			radix2 #(.width(width)) rd_st5_875  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[875]), .rdlo_in(a5_wr[891]),  .coef_in(coef[352]), .rdup_out(a6_wr[875]), .rdlo_out(a6_wr[891]));
			radix2 #(.width(width)) rd_st5_876  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[876]), .rdlo_in(a5_wr[892]),  .coef_in(coef[384]), .rdup_out(a6_wr[876]), .rdlo_out(a6_wr[892]));
			radix2 #(.width(width)) rd_st5_877  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[877]), .rdlo_in(a5_wr[893]),  .coef_in(coef[416]), .rdup_out(a6_wr[877]), .rdlo_out(a6_wr[893]));
			radix2 #(.width(width)) rd_st5_878  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[878]), .rdlo_in(a5_wr[894]),  .coef_in(coef[448]), .rdup_out(a6_wr[878]), .rdlo_out(a6_wr[894]));
			radix2 #(.width(width)) rd_st5_879  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[879]), .rdlo_in(a5_wr[895]),  .coef_in(coef[480]), .rdup_out(a6_wr[879]), .rdlo_out(a6_wr[895]));
			radix2 #(.width(width)) rd_st5_896  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[896]), .rdlo_in(a5_wr[912]),  .coef_in(coef[0]), .rdup_out(a6_wr[896]), .rdlo_out(a6_wr[912]));
			radix2 #(.width(width)) rd_st5_897  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[897]), .rdlo_in(a5_wr[913]),  .coef_in(coef[32]), .rdup_out(a6_wr[897]), .rdlo_out(a6_wr[913]));
			radix2 #(.width(width)) rd_st5_898  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[898]), .rdlo_in(a5_wr[914]),  .coef_in(coef[64]), .rdup_out(a6_wr[898]), .rdlo_out(a6_wr[914]));
			radix2 #(.width(width)) rd_st5_899  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[899]), .rdlo_in(a5_wr[915]),  .coef_in(coef[96]), .rdup_out(a6_wr[899]), .rdlo_out(a6_wr[915]));
			radix2 #(.width(width)) rd_st5_900  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[900]), .rdlo_in(a5_wr[916]),  .coef_in(coef[128]), .rdup_out(a6_wr[900]), .rdlo_out(a6_wr[916]));
			radix2 #(.width(width)) rd_st5_901  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[901]), .rdlo_in(a5_wr[917]),  .coef_in(coef[160]), .rdup_out(a6_wr[901]), .rdlo_out(a6_wr[917]));
			radix2 #(.width(width)) rd_st5_902  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[902]), .rdlo_in(a5_wr[918]),  .coef_in(coef[192]), .rdup_out(a6_wr[902]), .rdlo_out(a6_wr[918]));
			radix2 #(.width(width)) rd_st5_903  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[903]), .rdlo_in(a5_wr[919]),  .coef_in(coef[224]), .rdup_out(a6_wr[903]), .rdlo_out(a6_wr[919]));
			radix2 #(.width(width)) rd_st5_904  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[904]), .rdlo_in(a5_wr[920]),  .coef_in(coef[256]), .rdup_out(a6_wr[904]), .rdlo_out(a6_wr[920]));
			radix2 #(.width(width)) rd_st5_905  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[905]), .rdlo_in(a5_wr[921]),  .coef_in(coef[288]), .rdup_out(a6_wr[905]), .rdlo_out(a6_wr[921]));
			radix2 #(.width(width)) rd_st5_906  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[906]), .rdlo_in(a5_wr[922]),  .coef_in(coef[320]), .rdup_out(a6_wr[906]), .rdlo_out(a6_wr[922]));
			radix2 #(.width(width)) rd_st5_907  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[907]), .rdlo_in(a5_wr[923]),  .coef_in(coef[352]), .rdup_out(a6_wr[907]), .rdlo_out(a6_wr[923]));
			radix2 #(.width(width)) rd_st5_908  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[908]), .rdlo_in(a5_wr[924]),  .coef_in(coef[384]), .rdup_out(a6_wr[908]), .rdlo_out(a6_wr[924]));
			radix2 #(.width(width)) rd_st5_909  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[909]), .rdlo_in(a5_wr[925]),  .coef_in(coef[416]), .rdup_out(a6_wr[909]), .rdlo_out(a6_wr[925]));
			radix2 #(.width(width)) rd_st5_910  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[910]), .rdlo_in(a5_wr[926]),  .coef_in(coef[448]), .rdup_out(a6_wr[910]), .rdlo_out(a6_wr[926]));
			radix2 #(.width(width)) rd_st5_911  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[911]), .rdlo_in(a5_wr[927]),  .coef_in(coef[480]), .rdup_out(a6_wr[911]), .rdlo_out(a6_wr[927]));
			radix2 #(.width(width)) rd_st5_928  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[928]), .rdlo_in(a5_wr[944]),  .coef_in(coef[0]), .rdup_out(a6_wr[928]), .rdlo_out(a6_wr[944]));
			radix2 #(.width(width)) rd_st5_929  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[929]), .rdlo_in(a5_wr[945]),  .coef_in(coef[32]), .rdup_out(a6_wr[929]), .rdlo_out(a6_wr[945]));
			radix2 #(.width(width)) rd_st5_930  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[930]), .rdlo_in(a5_wr[946]),  .coef_in(coef[64]), .rdup_out(a6_wr[930]), .rdlo_out(a6_wr[946]));
			radix2 #(.width(width)) rd_st5_931  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[931]), .rdlo_in(a5_wr[947]),  .coef_in(coef[96]), .rdup_out(a6_wr[931]), .rdlo_out(a6_wr[947]));
			radix2 #(.width(width)) rd_st5_932  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[932]), .rdlo_in(a5_wr[948]),  .coef_in(coef[128]), .rdup_out(a6_wr[932]), .rdlo_out(a6_wr[948]));
			radix2 #(.width(width)) rd_st5_933  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[933]), .rdlo_in(a5_wr[949]),  .coef_in(coef[160]), .rdup_out(a6_wr[933]), .rdlo_out(a6_wr[949]));
			radix2 #(.width(width)) rd_st5_934  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[934]), .rdlo_in(a5_wr[950]),  .coef_in(coef[192]), .rdup_out(a6_wr[934]), .rdlo_out(a6_wr[950]));
			radix2 #(.width(width)) rd_st5_935  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[935]), .rdlo_in(a5_wr[951]),  .coef_in(coef[224]), .rdup_out(a6_wr[935]), .rdlo_out(a6_wr[951]));
			radix2 #(.width(width)) rd_st5_936  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[936]), .rdlo_in(a5_wr[952]),  .coef_in(coef[256]), .rdup_out(a6_wr[936]), .rdlo_out(a6_wr[952]));
			radix2 #(.width(width)) rd_st5_937  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[937]), .rdlo_in(a5_wr[953]),  .coef_in(coef[288]), .rdup_out(a6_wr[937]), .rdlo_out(a6_wr[953]));
			radix2 #(.width(width)) rd_st5_938  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[938]), .rdlo_in(a5_wr[954]),  .coef_in(coef[320]), .rdup_out(a6_wr[938]), .rdlo_out(a6_wr[954]));
			radix2 #(.width(width)) rd_st5_939  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[939]), .rdlo_in(a5_wr[955]),  .coef_in(coef[352]), .rdup_out(a6_wr[939]), .rdlo_out(a6_wr[955]));
			radix2 #(.width(width)) rd_st5_940  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[940]), .rdlo_in(a5_wr[956]),  .coef_in(coef[384]), .rdup_out(a6_wr[940]), .rdlo_out(a6_wr[956]));
			radix2 #(.width(width)) rd_st5_941  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[941]), .rdlo_in(a5_wr[957]),  .coef_in(coef[416]), .rdup_out(a6_wr[941]), .rdlo_out(a6_wr[957]));
			radix2 #(.width(width)) rd_st5_942  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[942]), .rdlo_in(a5_wr[958]),  .coef_in(coef[448]), .rdup_out(a6_wr[942]), .rdlo_out(a6_wr[958]));
			radix2 #(.width(width)) rd_st5_943  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[943]), .rdlo_in(a5_wr[959]),  .coef_in(coef[480]), .rdup_out(a6_wr[943]), .rdlo_out(a6_wr[959]));
			radix2 #(.width(width)) rd_st5_960  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[960]), .rdlo_in(a5_wr[976]),  .coef_in(coef[0]), .rdup_out(a6_wr[960]), .rdlo_out(a6_wr[976]));
			radix2 #(.width(width)) rd_st5_961  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[961]), .rdlo_in(a5_wr[977]),  .coef_in(coef[32]), .rdup_out(a6_wr[961]), .rdlo_out(a6_wr[977]));
			radix2 #(.width(width)) rd_st5_962  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[962]), .rdlo_in(a5_wr[978]),  .coef_in(coef[64]), .rdup_out(a6_wr[962]), .rdlo_out(a6_wr[978]));
			radix2 #(.width(width)) rd_st5_963  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[963]), .rdlo_in(a5_wr[979]),  .coef_in(coef[96]), .rdup_out(a6_wr[963]), .rdlo_out(a6_wr[979]));
			radix2 #(.width(width)) rd_st5_964  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[964]), .rdlo_in(a5_wr[980]),  .coef_in(coef[128]), .rdup_out(a6_wr[964]), .rdlo_out(a6_wr[980]));
			radix2 #(.width(width)) rd_st5_965  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[965]), .rdlo_in(a5_wr[981]),  .coef_in(coef[160]), .rdup_out(a6_wr[965]), .rdlo_out(a6_wr[981]));
			radix2 #(.width(width)) rd_st5_966  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[966]), .rdlo_in(a5_wr[982]),  .coef_in(coef[192]), .rdup_out(a6_wr[966]), .rdlo_out(a6_wr[982]));
			radix2 #(.width(width)) rd_st5_967  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[967]), .rdlo_in(a5_wr[983]),  .coef_in(coef[224]), .rdup_out(a6_wr[967]), .rdlo_out(a6_wr[983]));
			radix2 #(.width(width)) rd_st5_968  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[968]), .rdlo_in(a5_wr[984]),  .coef_in(coef[256]), .rdup_out(a6_wr[968]), .rdlo_out(a6_wr[984]));
			radix2 #(.width(width)) rd_st5_969  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[969]), .rdlo_in(a5_wr[985]),  .coef_in(coef[288]), .rdup_out(a6_wr[969]), .rdlo_out(a6_wr[985]));
			radix2 #(.width(width)) rd_st5_970  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[970]), .rdlo_in(a5_wr[986]),  .coef_in(coef[320]), .rdup_out(a6_wr[970]), .rdlo_out(a6_wr[986]));
			radix2 #(.width(width)) rd_st5_971  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[971]), .rdlo_in(a5_wr[987]),  .coef_in(coef[352]), .rdup_out(a6_wr[971]), .rdlo_out(a6_wr[987]));
			radix2 #(.width(width)) rd_st5_972  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[972]), .rdlo_in(a5_wr[988]),  .coef_in(coef[384]), .rdup_out(a6_wr[972]), .rdlo_out(a6_wr[988]));
			radix2 #(.width(width)) rd_st5_973  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[973]), .rdlo_in(a5_wr[989]),  .coef_in(coef[416]), .rdup_out(a6_wr[973]), .rdlo_out(a6_wr[989]));
			radix2 #(.width(width)) rd_st5_974  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[974]), .rdlo_in(a5_wr[990]),  .coef_in(coef[448]), .rdup_out(a6_wr[974]), .rdlo_out(a6_wr[990]));
			radix2 #(.width(width)) rd_st5_975  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[975]), .rdlo_in(a5_wr[991]),  .coef_in(coef[480]), .rdup_out(a6_wr[975]), .rdlo_out(a6_wr[991]));
			radix2 #(.width(width)) rd_st5_992  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[992]), .rdlo_in(a5_wr[1008]),  .coef_in(coef[0]), .rdup_out(a6_wr[992]), .rdlo_out(a6_wr[1008]));
			radix2 #(.width(width)) rd_st5_993  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[993]), .rdlo_in(a5_wr[1009]),  .coef_in(coef[32]), .rdup_out(a6_wr[993]), .rdlo_out(a6_wr[1009]));
			radix2 #(.width(width)) rd_st5_994  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[994]), .rdlo_in(a5_wr[1010]),  .coef_in(coef[64]), .rdup_out(a6_wr[994]), .rdlo_out(a6_wr[1010]));
			radix2 #(.width(width)) rd_st5_995  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[995]), .rdlo_in(a5_wr[1011]),  .coef_in(coef[96]), .rdup_out(a6_wr[995]), .rdlo_out(a6_wr[1011]));
			radix2 #(.width(width)) rd_st5_996  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[996]), .rdlo_in(a5_wr[1012]),  .coef_in(coef[128]), .rdup_out(a6_wr[996]), .rdlo_out(a6_wr[1012]));
			radix2 #(.width(width)) rd_st5_997  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[997]), .rdlo_in(a5_wr[1013]),  .coef_in(coef[160]), .rdup_out(a6_wr[997]), .rdlo_out(a6_wr[1013]));
			radix2 #(.width(width)) rd_st5_998  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[998]), .rdlo_in(a5_wr[1014]),  .coef_in(coef[192]), .rdup_out(a6_wr[998]), .rdlo_out(a6_wr[1014]));
			radix2 #(.width(width)) rd_st5_999  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[999]), .rdlo_in(a5_wr[1015]),  .coef_in(coef[224]), .rdup_out(a6_wr[999]), .rdlo_out(a6_wr[1015]));
			radix2 #(.width(width)) rd_st5_1000  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1000]), .rdlo_in(a5_wr[1016]),  .coef_in(coef[256]), .rdup_out(a6_wr[1000]), .rdlo_out(a6_wr[1016]));
			radix2 #(.width(width)) rd_st5_1001  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1001]), .rdlo_in(a5_wr[1017]),  .coef_in(coef[288]), .rdup_out(a6_wr[1001]), .rdlo_out(a6_wr[1017]));
			radix2 #(.width(width)) rd_st5_1002  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1002]), .rdlo_in(a5_wr[1018]),  .coef_in(coef[320]), .rdup_out(a6_wr[1002]), .rdlo_out(a6_wr[1018]));
			radix2 #(.width(width)) rd_st5_1003  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1003]), .rdlo_in(a5_wr[1019]),  .coef_in(coef[352]), .rdup_out(a6_wr[1003]), .rdlo_out(a6_wr[1019]));
			radix2 #(.width(width)) rd_st5_1004  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1004]), .rdlo_in(a5_wr[1020]),  .coef_in(coef[384]), .rdup_out(a6_wr[1004]), .rdlo_out(a6_wr[1020]));
			radix2 #(.width(width)) rd_st5_1005  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1005]), .rdlo_in(a5_wr[1021]),  .coef_in(coef[416]), .rdup_out(a6_wr[1005]), .rdlo_out(a6_wr[1021]));
			radix2 #(.width(width)) rd_st5_1006  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1006]), .rdlo_in(a5_wr[1022]),  .coef_in(coef[448]), .rdup_out(a6_wr[1006]), .rdlo_out(a6_wr[1022]));
			radix2 #(.width(width)) rd_st5_1007  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1007]), .rdlo_in(a5_wr[1023]),  .coef_in(coef[480]), .rdup_out(a6_wr[1007]), .rdlo_out(a6_wr[1023]));

		//--- radix stage 6
			radix2 #(.width(width)) rd_st6_0   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[0]), .rdlo_in(a6_wr[8]),  .coef_in(coef[0]), .rdup_out(a7_wr[0]), .rdlo_out(a7_wr[8]));
			radix2 #(.width(width)) rd_st6_1   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1]), .rdlo_in(a6_wr[9]),  .coef_in(coef[64]), .rdup_out(a7_wr[1]), .rdlo_out(a7_wr[9]));
			radix2 #(.width(width)) rd_st6_2   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[2]), .rdlo_in(a6_wr[10]),  .coef_in(coef[128]), .rdup_out(a7_wr[2]), .rdlo_out(a7_wr[10]));
			radix2 #(.width(width)) rd_st6_3   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[3]), .rdlo_in(a6_wr[11]),  .coef_in(coef[192]), .rdup_out(a7_wr[3]), .rdlo_out(a7_wr[11]));
			radix2 #(.width(width)) rd_st6_4   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[4]), .rdlo_in(a6_wr[12]),  .coef_in(coef[256]), .rdup_out(a7_wr[4]), .rdlo_out(a7_wr[12]));
			radix2 #(.width(width)) rd_st6_5   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[5]), .rdlo_in(a6_wr[13]),  .coef_in(coef[320]), .rdup_out(a7_wr[5]), .rdlo_out(a7_wr[13]));
			radix2 #(.width(width)) rd_st6_6   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[6]), .rdlo_in(a6_wr[14]),  .coef_in(coef[384]), .rdup_out(a7_wr[6]), .rdlo_out(a7_wr[14]));
			radix2 #(.width(width)) rd_st6_7   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[7]), .rdlo_in(a6_wr[15]),  .coef_in(coef[448]), .rdup_out(a7_wr[7]), .rdlo_out(a7_wr[15]));
			radix2 #(.width(width)) rd_st6_16  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[16]), .rdlo_in(a6_wr[24]),  .coef_in(coef[0]), .rdup_out(a7_wr[16]), .rdlo_out(a7_wr[24]));
			radix2 #(.width(width)) rd_st6_17  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[17]), .rdlo_in(a6_wr[25]),  .coef_in(coef[64]), .rdup_out(a7_wr[17]), .rdlo_out(a7_wr[25]));
			radix2 #(.width(width)) rd_st6_18  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[18]), .rdlo_in(a6_wr[26]),  .coef_in(coef[128]), .rdup_out(a7_wr[18]), .rdlo_out(a7_wr[26]));
			radix2 #(.width(width)) rd_st6_19  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[19]), .rdlo_in(a6_wr[27]),  .coef_in(coef[192]), .rdup_out(a7_wr[19]), .rdlo_out(a7_wr[27]));
			radix2 #(.width(width)) rd_st6_20  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[20]), .rdlo_in(a6_wr[28]),  .coef_in(coef[256]), .rdup_out(a7_wr[20]), .rdlo_out(a7_wr[28]));
			radix2 #(.width(width)) rd_st6_21  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[21]), .rdlo_in(a6_wr[29]),  .coef_in(coef[320]), .rdup_out(a7_wr[21]), .rdlo_out(a7_wr[29]));
			radix2 #(.width(width)) rd_st6_22  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[22]), .rdlo_in(a6_wr[30]),  .coef_in(coef[384]), .rdup_out(a7_wr[22]), .rdlo_out(a7_wr[30]));
			radix2 #(.width(width)) rd_st6_23  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[23]), .rdlo_in(a6_wr[31]),  .coef_in(coef[448]), .rdup_out(a7_wr[23]), .rdlo_out(a7_wr[31]));
			radix2 #(.width(width)) rd_st6_32  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[32]), .rdlo_in(a6_wr[40]),  .coef_in(coef[0]), .rdup_out(a7_wr[32]), .rdlo_out(a7_wr[40]));
			radix2 #(.width(width)) rd_st6_33  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[33]), .rdlo_in(a6_wr[41]),  .coef_in(coef[64]), .rdup_out(a7_wr[33]), .rdlo_out(a7_wr[41]));
			radix2 #(.width(width)) rd_st6_34  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[34]), .rdlo_in(a6_wr[42]),  .coef_in(coef[128]), .rdup_out(a7_wr[34]), .rdlo_out(a7_wr[42]));
			radix2 #(.width(width)) rd_st6_35  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[35]), .rdlo_in(a6_wr[43]),  .coef_in(coef[192]), .rdup_out(a7_wr[35]), .rdlo_out(a7_wr[43]));
			radix2 #(.width(width)) rd_st6_36  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[36]), .rdlo_in(a6_wr[44]),  .coef_in(coef[256]), .rdup_out(a7_wr[36]), .rdlo_out(a7_wr[44]));
			radix2 #(.width(width)) rd_st6_37  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[37]), .rdlo_in(a6_wr[45]),  .coef_in(coef[320]), .rdup_out(a7_wr[37]), .rdlo_out(a7_wr[45]));
			radix2 #(.width(width)) rd_st6_38  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[38]), .rdlo_in(a6_wr[46]),  .coef_in(coef[384]), .rdup_out(a7_wr[38]), .rdlo_out(a7_wr[46]));
			radix2 #(.width(width)) rd_st6_39  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[39]), .rdlo_in(a6_wr[47]),  .coef_in(coef[448]), .rdup_out(a7_wr[39]), .rdlo_out(a7_wr[47]));
			radix2 #(.width(width)) rd_st6_48  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[48]), .rdlo_in(a6_wr[56]),  .coef_in(coef[0]), .rdup_out(a7_wr[48]), .rdlo_out(a7_wr[56]));
			radix2 #(.width(width)) rd_st6_49  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[49]), .rdlo_in(a6_wr[57]),  .coef_in(coef[64]), .rdup_out(a7_wr[49]), .rdlo_out(a7_wr[57]));
			radix2 #(.width(width)) rd_st6_50  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[50]), .rdlo_in(a6_wr[58]),  .coef_in(coef[128]), .rdup_out(a7_wr[50]), .rdlo_out(a7_wr[58]));
			radix2 #(.width(width)) rd_st6_51  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[51]), .rdlo_in(a6_wr[59]),  .coef_in(coef[192]), .rdup_out(a7_wr[51]), .rdlo_out(a7_wr[59]));
			radix2 #(.width(width)) rd_st6_52  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[52]), .rdlo_in(a6_wr[60]),  .coef_in(coef[256]), .rdup_out(a7_wr[52]), .rdlo_out(a7_wr[60]));
			radix2 #(.width(width)) rd_st6_53  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[53]), .rdlo_in(a6_wr[61]),  .coef_in(coef[320]), .rdup_out(a7_wr[53]), .rdlo_out(a7_wr[61]));
			radix2 #(.width(width)) rd_st6_54  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[54]), .rdlo_in(a6_wr[62]),  .coef_in(coef[384]), .rdup_out(a7_wr[54]), .rdlo_out(a7_wr[62]));
			radix2 #(.width(width)) rd_st6_55  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[55]), .rdlo_in(a6_wr[63]),  .coef_in(coef[448]), .rdup_out(a7_wr[55]), .rdlo_out(a7_wr[63]));
			radix2 #(.width(width)) rd_st6_64  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[64]), .rdlo_in(a6_wr[72]),  .coef_in(coef[0]), .rdup_out(a7_wr[64]), .rdlo_out(a7_wr[72]));
			radix2 #(.width(width)) rd_st6_65  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[65]), .rdlo_in(a6_wr[73]),  .coef_in(coef[64]), .rdup_out(a7_wr[65]), .rdlo_out(a7_wr[73]));
			radix2 #(.width(width)) rd_st6_66  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[66]), .rdlo_in(a6_wr[74]),  .coef_in(coef[128]), .rdup_out(a7_wr[66]), .rdlo_out(a7_wr[74]));
			radix2 #(.width(width)) rd_st6_67  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[67]), .rdlo_in(a6_wr[75]),  .coef_in(coef[192]), .rdup_out(a7_wr[67]), .rdlo_out(a7_wr[75]));
			radix2 #(.width(width)) rd_st6_68  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[68]), .rdlo_in(a6_wr[76]),  .coef_in(coef[256]), .rdup_out(a7_wr[68]), .rdlo_out(a7_wr[76]));
			radix2 #(.width(width)) rd_st6_69  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[69]), .rdlo_in(a6_wr[77]),  .coef_in(coef[320]), .rdup_out(a7_wr[69]), .rdlo_out(a7_wr[77]));
			radix2 #(.width(width)) rd_st6_70  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[70]), .rdlo_in(a6_wr[78]),  .coef_in(coef[384]), .rdup_out(a7_wr[70]), .rdlo_out(a7_wr[78]));
			radix2 #(.width(width)) rd_st6_71  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[71]), .rdlo_in(a6_wr[79]),  .coef_in(coef[448]), .rdup_out(a7_wr[71]), .rdlo_out(a7_wr[79]));
			radix2 #(.width(width)) rd_st6_80  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[80]), .rdlo_in(a6_wr[88]),  .coef_in(coef[0]), .rdup_out(a7_wr[80]), .rdlo_out(a7_wr[88]));
			radix2 #(.width(width)) rd_st6_81  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[81]), .rdlo_in(a6_wr[89]),  .coef_in(coef[64]), .rdup_out(a7_wr[81]), .rdlo_out(a7_wr[89]));
			radix2 #(.width(width)) rd_st6_82  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[82]), .rdlo_in(a6_wr[90]),  .coef_in(coef[128]), .rdup_out(a7_wr[82]), .rdlo_out(a7_wr[90]));
			radix2 #(.width(width)) rd_st6_83  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[83]), .rdlo_in(a6_wr[91]),  .coef_in(coef[192]), .rdup_out(a7_wr[83]), .rdlo_out(a7_wr[91]));
			radix2 #(.width(width)) rd_st6_84  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[84]), .rdlo_in(a6_wr[92]),  .coef_in(coef[256]), .rdup_out(a7_wr[84]), .rdlo_out(a7_wr[92]));
			radix2 #(.width(width)) rd_st6_85  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[85]), .rdlo_in(a6_wr[93]),  .coef_in(coef[320]), .rdup_out(a7_wr[85]), .rdlo_out(a7_wr[93]));
			radix2 #(.width(width)) rd_st6_86  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[86]), .rdlo_in(a6_wr[94]),  .coef_in(coef[384]), .rdup_out(a7_wr[86]), .rdlo_out(a7_wr[94]));
			radix2 #(.width(width)) rd_st6_87  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[87]), .rdlo_in(a6_wr[95]),  .coef_in(coef[448]), .rdup_out(a7_wr[87]), .rdlo_out(a7_wr[95]));
			radix2 #(.width(width)) rd_st6_96  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[96]), .rdlo_in(a6_wr[104]),  .coef_in(coef[0]), .rdup_out(a7_wr[96]), .rdlo_out(a7_wr[104]));
			radix2 #(.width(width)) rd_st6_97  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[97]), .rdlo_in(a6_wr[105]),  .coef_in(coef[64]), .rdup_out(a7_wr[97]), .rdlo_out(a7_wr[105]));
			radix2 #(.width(width)) rd_st6_98  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[98]), .rdlo_in(a6_wr[106]),  .coef_in(coef[128]), .rdup_out(a7_wr[98]), .rdlo_out(a7_wr[106]));
			radix2 #(.width(width)) rd_st6_99  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[99]), .rdlo_in(a6_wr[107]),  .coef_in(coef[192]), .rdup_out(a7_wr[99]), .rdlo_out(a7_wr[107]));
			radix2 #(.width(width)) rd_st6_100  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[100]), .rdlo_in(a6_wr[108]),  .coef_in(coef[256]), .rdup_out(a7_wr[100]), .rdlo_out(a7_wr[108]));
			radix2 #(.width(width)) rd_st6_101  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[101]), .rdlo_in(a6_wr[109]),  .coef_in(coef[320]), .rdup_out(a7_wr[101]), .rdlo_out(a7_wr[109]));
			radix2 #(.width(width)) rd_st6_102  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[102]), .rdlo_in(a6_wr[110]),  .coef_in(coef[384]), .rdup_out(a7_wr[102]), .rdlo_out(a7_wr[110]));
			radix2 #(.width(width)) rd_st6_103  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[103]), .rdlo_in(a6_wr[111]),  .coef_in(coef[448]), .rdup_out(a7_wr[103]), .rdlo_out(a7_wr[111]));
			radix2 #(.width(width)) rd_st6_112  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[112]), .rdlo_in(a6_wr[120]),  .coef_in(coef[0]), .rdup_out(a7_wr[112]), .rdlo_out(a7_wr[120]));
			radix2 #(.width(width)) rd_st6_113  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[113]), .rdlo_in(a6_wr[121]),  .coef_in(coef[64]), .rdup_out(a7_wr[113]), .rdlo_out(a7_wr[121]));
			radix2 #(.width(width)) rd_st6_114  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[114]), .rdlo_in(a6_wr[122]),  .coef_in(coef[128]), .rdup_out(a7_wr[114]), .rdlo_out(a7_wr[122]));
			radix2 #(.width(width)) rd_st6_115  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[115]), .rdlo_in(a6_wr[123]),  .coef_in(coef[192]), .rdup_out(a7_wr[115]), .rdlo_out(a7_wr[123]));
			radix2 #(.width(width)) rd_st6_116  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[116]), .rdlo_in(a6_wr[124]),  .coef_in(coef[256]), .rdup_out(a7_wr[116]), .rdlo_out(a7_wr[124]));
			radix2 #(.width(width)) rd_st6_117  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[117]), .rdlo_in(a6_wr[125]),  .coef_in(coef[320]), .rdup_out(a7_wr[117]), .rdlo_out(a7_wr[125]));
			radix2 #(.width(width)) rd_st6_118  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[118]), .rdlo_in(a6_wr[126]),  .coef_in(coef[384]), .rdup_out(a7_wr[118]), .rdlo_out(a7_wr[126]));
			radix2 #(.width(width)) rd_st6_119  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[119]), .rdlo_in(a6_wr[127]),  .coef_in(coef[448]), .rdup_out(a7_wr[119]), .rdlo_out(a7_wr[127]));
			radix2 #(.width(width)) rd_st6_128  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[128]), .rdlo_in(a6_wr[136]),  .coef_in(coef[0]), .rdup_out(a7_wr[128]), .rdlo_out(a7_wr[136]));
			radix2 #(.width(width)) rd_st6_129  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[129]), .rdlo_in(a6_wr[137]),  .coef_in(coef[64]), .rdup_out(a7_wr[129]), .rdlo_out(a7_wr[137]));
			radix2 #(.width(width)) rd_st6_130  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[130]), .rdlo_in(a6_wr[138]),  .coef_in(coef[128]), .rdup_out(a7_wr[130]), .rdlo_out(a7_wr[138]));
			radix2 #(.width(width)) rd_st6_131  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[131]), .rdlo_in(a6_wr[139]),  .coef_in(coef[192]), .rdup_out(a7_wr[131]), .rdlo_out(a7_wr[139]));
			radix2 #(.width(width)) rd_st6_132  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[132]), .rdlo_in(a6_wr[140]),  .coef_in(coef[256]), .rdup_out(a7_wr[132]), .rdlo_out(a7_wr[140]));
			radix2 #(.width(width)) rd_st6_133  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[133]), .rdlo_in(a6_wr[141]),  .coef_in(coef[320]), .rdup_out(a7_wr[133]), .rdlo_out(a7_wr[141]));
			radix2 #(.width(width)) rd_st6_134  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[134]), .rdlo_in(a6_wr[142]),  .coef_in(coef[384]), .rdup_out(a7_wr[134]), .rdlo_out(a7_wr[142]));
			radix2 #(.width(width)) rd_st6_135  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[135]), .rdlo_in(a6_wr[143]),  .coef_in(coef[448]), .rdup_out(a7_wr[135]), .rdlo_out(a7_wr[143]));
			radix2 #(.width(width)) rd_st6_144  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[144]), .rdlo_in(a6_wr[152]),  .coef_in(coef[0]), .rdup_out(a7_wr[144]), .rdlo_out(a7_wr[152]));
			radix2 #(.width(width)) rd_st6_145  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[145]), .rdlo_in(a6_wr[153]),  .coef_in(coef[64]), .rdup_out(a7_wr[145]), .rdlo_out(a7_wr[153]));
			radix2 #(.width(width)) rd_st6_146  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[146]), .rdlo_in(a6_wr[154]),  .coef_in(coef[128]), .rdup_out(a7_wr[146]), .rdlo_out(a7_wr[154]));
			radix2 #(.width(width)) rd_st6_147  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[147]), .rdlo_in(a6_wr[155]),  .coef_in(coef[192]), .rdup_out(a7_wr[147]), .rdlo_out(a7_wr[155]));
			radix2 #(.width(width)) rd_st6_148  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[148]), .rdlo_in(a6_wr[156]),  .coef_in(coef[256]), .rdup_out(a7_wr[148]), .rdlo_out(a7_wr[156]));
			radix2 #(.width(width)) rd_st6_149  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[149]), .rdlo_in(a6_wr[157]),  .coef_in(coef[320]), .rdup_out(a7_wr[149]), .rdlo_out(a7_wr[157]));
			radix2 #(.width(width)) rd_st6_150  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[150]), .rdlo_in(a6_wr[158]),  .coef_in(coef[384]), .rdup_out(a7_wr[150]), .rdlo_out(a7_wr[158]));
			radix2 #(.width(width)) rd_st6_151  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[151]), .rdlo_in(a6_wr[159]),  .coef_in(coef[448]), .rdup_out(a7_wr[151]), .rdlo_out(a7_wr[159]));
			radix2 #(.width(width)) rd_st6_160  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[160]), .rdlo_in(a6_wr[168]),  .coef_in(coef[0]), .rdup_out(a7_wr[160]), .rdlo_out(a7_wr[168]));
			radix2 #(.width(width)) rd_st6_161  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[161]), .rdlo_in(a6_wr[169]),  .coef_in(coef[64]), .rdup_out(a7_wr[161]), .rdlo_out(a7_wr[169]));
			radix2 #(.width(width)) rd_st6_162  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[162]), .rdlo_in(a6_wr[170]),  .coef_in(coef[128]), .rdup_out(a7_wr[162]), .rdlo_out(a7_wr[170]));
			radix2 #(.width(width)) rd_st6_163  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[163]), .rdlo_in(a6_wr[171]),  .coef_in(coef[192]), .rdup_out(a7_wr[163]), .rdlo_out(a7_wr[171]));
			radix2 #(.width(width)) rd_st6_164  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[164]), .rdlo_in(a6_wr[172]),  .coef_in(coef[256]), .rdup_out(a7_wr[164]), .rdlo_out(a7_wr[172]));
			radix2 #(.width(width)) rd_st6_165  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[165]), .rdlo_in(a6_wr[173]),  .coef_in(coef[320]), .rdup_out(a7_wr[165]), .rdlo_out(a7_wr[173]));
			radix2 #(.width(width)) rd_st6_166  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[166]), .rdlo_in(a6_wr[174]),  .coef_in(coef[384]), .rdup_out(a7_wr[166]), .rdlo_out(a7_wr[174]));
			radix2 #(.width(width)) rd_st6_167  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[167]), .rdlo_in(a6_wr[175]),  .coef_in(coef[448]), .rdup_out(a7_wr[167]), .rdlo_out(a7_wr[175]));
			radix2 #(.width(width)) rd_st6_176  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[176]), .rdlo_in(a6_wr[184]),  .coef_in(coef[0]), .rdup_out(a7_wr[176]), .rdlo_out(a7_wr[184]));
			radix2 #(.width(width)) rd_st6_177  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[177]), .rdlo_in(a6_wr[185]),  .coef_in(coef[64]), .rdup_out(a7_wr[177]), .rdlo_out(a7_wr[185]));
			radix2 #(.width(width)) rd_st6_178  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[178]), .rdlo_in(a6_wr[186]),  .coef_in(coef[128]), .rdup_out(a7_wr[178]), .rdlo_out(a7_wr[186]));
			radix2 #(.width(width)) rd_st6_179  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[179]), .rdlo_in(a6_wr[187]),  .coef_in(coef[192]), .rdup_out(a7_wr[179]), .rdlo_out(a7_wr[187]));
			radix2 #(.width(width)) rd_st6_180  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[180]), .rdlo_in(a6_wr[188]),  .coef_in(coef[256]), .rdup_out(a7_wr[180]), .rdlo_out(a7_wr[188]));
			radix2 #(.width(width)) rd_st6_181  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[181]), .rdlo_in(a6_wr[189]),  .coef_in(coef[320]), .rdup_out(a7_wr[181]), .rdlo_out(a7_wr[189]));
			radix2 #(.width(width)) rd_st6_182  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[182]), .rdlo_in(a6_wr[190]),  .coef_in(coef[384]), .rdup_out(a7_wr[182]), .rdlo_out(a7_wr[190]));
			radix2 #(.width(width)) rd_st6_183  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[183]), .rdlo_in(a6_wr[191]),  .coef_in(coef[448]), .rdup_out(a7_wr[183]), .rdlo_out(a7_wr[191]));
			radix2 #(.width(width)) rd_st6_192  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[192]), .rdlo_in(a6_wr[200]),  .coef_in(coef[0]), .rdup_out(a7_wr[192]), .rdlo_out(a7_wr[200]));
			radix2 #(.width(width)) rd_st6_193  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[193]), .rdlo_in(a6_wr[201]),  .coef_in(coef[64]), .rdup_out(a7_wr[193]), .rdlo_out(a7_wr[201]));
			radix2 #(.width(width)) rd_st6_194  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[194]), .rdlo_in(a6_wr[202]),  .coef_in(coef[128]), .rdup_out(a7_wr[194]), .rdlo_out(a7_wr[202]));
			radix2 #(.width(width)) rd_st6_195  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[195]), .rdlo_in(a6_wr[203]),  .coef_in(coef[192]), .rdup_out(a7_wr[195]), .rdlo_out(a7_wr[203]));
			radix2 #(.width(width)) rd_st6_196  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[196]), .rdlo_in(a6_wr[204]),  .coef_in(coef[256]), .rdup_out(a7_wr[196]), .rdlo_out(a7_wr[204]));
			radix2 #(.width(width)) rd_st6_197  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[197]), .rdlo_in(a6_wr[205]),  .coef_in(coef[320]), .rdup_out(a7_wr[197]), .rdlo_out(a7_wr[205]));
			radix2 #(.width(width)) rd_st6_198  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[198]), .rdlo_in(a6_wr[206]),  .coef_in(coef[384]), .rdup_out(a7_wr[198]), .rdlo_out(a7_wr[206]));
			radix2 #(.width(width)) rd_st6_199  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[199]), .rdlo_in(a6_wr[207]),  .coef_in(coef[448]), .rdup_out(a7_wr[199]), .rdlo_out(a7_wr[207]));
			radix2 #(.width(width)) rd_st6_208  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[208]), .rdlo_in(a6_wr[216]),  .coef_in(coef[0]), .rdup_out(a7_wr[208]), .rdlo_out(a7_wr[216]));
			radix2 #(.width(width)) rd_st6_209  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[209]), .rdlo_in(a6_wr[217]),  .coef_in(coef[64]), .rdup_out(a7_wr[209]), .rdlo_out(a7_wr[217]));
			radix2 #(.width(width)) rd_st6_210  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[210]), .rdlo_in(a6_wr[218]),  .coef_in(coef[128]), .rdup_out(a7_wr[210]), .rdlo_out(a7_wr[218]));
			radix2 #(.width(width)) rd_st6_211  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[211]), .rdlo_in(a6_wr[219]),  .coef_in(coef[192]), .rdup_out(a7_wr[211]), .rdlo_out(a7_wr[219]));
			radix2 #(.width(width)) rd_st6_212  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[212]), .rdlo_in(a6_wr[220]),  .coef_in(coef[256]), .rdup_out(a7_wr[212]), .rdlo_out(a7_wr[220]));
			radix2 #(.width(width)) rd_st6_213  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[213]), .rdlo_in(a6_wr[221]),  .coef_in(coef[320]), .rdup_out(a7_wr[213]), .rdlo_out(a7_wr[221]));
			radix2 #(.width(width)) rd_st6_214  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[214]), .rdlo_in(a6_wr[222]),  .coef_in(coef[384]), .rdup_out(a7_wr[214]), .rdlo_out(a7_wr[222]));
			radix2 #(.width(width)) rd_st6_215  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[215]), .rdlo_in(a6_wr[223]),  .coef_in(coef[448]), .rdup_out(a7_wr[215]), .rdlo_out(a7_wr[223]));
			radix2 #(.width(width)) rd_st6_224  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[224]), .rdlo_in(a6_wr[232]),  .coef_in(coef[0]), .rdup_out(a7_wr[224]), .rdlo_out(a7_wr[232]));
			radix2 #(.width(width)) rd_st6_225  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[225]), .rdlo_in(a6_wr[233]),  .coef_in(coef[64]), .rdup_out(a7_wr[225]), .rdlo_out(a7_wr[233]));
			radix2 #(.width(width)) rd_st6_226  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[226]), .rdlo_in(a6_wr[234]),  .coef_in(coef[128]), .rdup_out(a7_wr[226]), .rdlo_out(a7_wr[234]));
			radix2 #(.width(width)) rd_st6_227  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[227]), .rdlo_in(a6_wr[235]),  .coef_in(coef[192]), .rdup_out(a7_wr[227]), .rdlo_out(a7_wr[235]));
			radix2 #(.width(width)) rd_st6_228  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[228]), .rdlo_in(a6_wr[236]),  .coef_in(coef[256]), .rdup_out(a7_wr[228]), .rdlo_out(a7_wr[236]));
			radix2 #(.width(width)) rd_st6_229  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[229]), .rdlo_in(a6_wr[237]),  .coef_in(coef[320]), .rdup_out(a7_wr[229]), .rdlo_out(a7_wr[237]));
			radix2 #(.width(width)) rd_st6_230  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[230]), .rdlo_in(a6_wr[238]),  .coef_in(coef[384]), .rdup_out(a7_wr[230]), .rdlo_out(a7_wr[238]));
			radix2 #(.width(width)) rd_st6_231  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[231]), .rdlo_in(a6_wr[239]),  .coef_in(coef[448]), .rdup_out(a7_wr[231]), .rdlo_out(a7_wr[239]));
			radix2 #(.width(width)) rd_st6_240  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[240]), .rdlo_in(a6_wr[248]),  .coef_in(coef[0]), .rdup_out(a7_wr[240]), .rdlo_out(a7_wr[248]));
			radix2 #(.width(width)) rd_st6_241  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[241]), .rdlo_in(a6_wr[249]),  .coef_in(coef[64]), .rdup_out(a7_wr[241]), .rdlo_out(a7_wr[249]));
			radix2 #(.width(width)) rd_st6_242  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[242]), .rdlo_in(a6_wr[250]),  .coef_in(coef[128]), .rdup_out(a7_wr[242]), .rdlo_out(a7_wr[250]));
			radix2 #(.width(width)) rd_st6_243  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[243]), .rdlo_in(a6_wr[251]),  .coef_in(coef[192]), .rdup_out(a7_wr[243]), .rdlo_out(a7_wr[251]));
			radix2 #(.width(width)) rd_st6_244  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[244]), .rdlo_in(a6_wr[252]),  .coef_in(coef[256]), .rdup_out(a7_wr[244]), .rdlo_out(a7_wr[252]));
			radix2 #(.width(width)) rd_st6_245  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[245]), .rdlo_in(a6_wr[253]),  .coef_in(coef[320]), .rdup_out(a7_wr[245]), .rdlo_out(a7_wr[253]));
			radix2 #(.width(width)) rd_st6_246  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[246]), .rdlo_in(a6_wr[254]),  .coef_in(coef[384]), .rdup_out(a7_wr[246]), .rdlo_out(a7_wr[254]));
			radix2 #(.width(width)) rd_st6_247  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[247]), .rdlo_in(a6_wr[255]),  .coef_in(coef[448]), .rdup_out(a7_wr[247]), .rdlo_out(a7_wr[255]));
			radix2 #(.width(width)) rd_st6_256  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[256]), .rdlo_in(a6_wr[264]),  .coef_in(coef[0]), .rdup_out(a7_wr[256]), .rdlo_out(a7_wr[264]));
			radix2 #(.width(width)) rd_st6_257  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[257]), .rdlo_in(a6_wr[265]),  .coef_in(coef[64]), .rdup_out(a7_wr[257]), .rdlo_out(a7_wr[265]));
			radix2 #(.width(width)) rd_st6_258  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[258]), .rdlo_in(a6_wr[266]),  .coef_in(coef[128]), .rdup_out(a7_wr[258]), .rdlo_out(a7_wr[266]));
			radix2 #(.width(width)) rd_st6_259  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[259]), .rdlo_in(a6_wr[267]),  .coef_in(coef[192]), .rdup_out(a7_wr[259]), .rdlo_out(a7_wr[267]));
			radix2 #(.width(width)) rd_st6_260  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[260]), .rdlo_in(a6_wr[268]),  .coef_in(coef[256]), .rdup_out(a7_wr[260]), .rdlo_out(a7_wr[268]));
			radix2 #(.width(width)) rd_st6_261  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[261]), .rdlo_in(a6_wr[269]),  .coef_in(coef[320]), .rdup_out(a7_wr[261]), .rdlo_out(a7_wr[269]));
			radix2 #(.width(width)) rd_st6_262  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[262]), .rdlo_in(a6_wr[270]),  .coef_in(coef[384]), .rdup_out(a7_wr[262]), .rdlo_out(a7_wr[270]));
			radix2 #(.width(width)) rd_st6_263  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[263]), .rdlo_in(a6_wr[271]),  .coef_in(coef[448]), .rdup_out(a7_wr[263]), .rdlo_out(a7_wr[271]));
			radix2 #(.width(width)) rd_st6_272  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[272]), .rdlo_in(a6_wr[280]),  .coef_in(coef[0]), .rdup_out(a7_wr[272]), .rdlo_out(a7_wr[280]));
			radix2 #(.width(width)) rd_st6_273  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[273]), .rdlo_in(a6_wr[281]),  .coef_in(coef[64]), .rdup_out(a7_wr[273]), .rdlo_out(a7_wr[281]));
			radix2 #(.width(width)) rd_st6_274  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[274]), .rdlo_in(a6_wr[282]),  .coef_in(coef[128]), .rdup_out(a7_wr[274]), .rdlo_out(a7_wr[282]));
			radix2 #(.width(width)) rd_st6_275  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[275]), .rdlo_in(a6_wr[283]),  .coef_in(coef[192]), .rdup_out(a7_wr[275]), .rdlo_out(a7_wr[283]));
			radix2 #(.width(width)) rd_st6_276  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[276]), .rdlo_in(a6_wr[284]),  .coef_in(coef[256]), .rdup_out(a7_wr[276]), .rdlo_out(a7_wr[284]));
			radix2 #(.width(width)) rd_st6_277  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[277]), .rdlo_in(a6_wr[285]),  .coef_in(coef[320]), .rdup_out(a7_wr[277]), .rdlo_out(a7_wr[285]));
			radix2 #(.width(width)) rd_st6_278  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[278]), .rdlo_in(a6_wr[286]),  .coef_in(coef[384]), .rdup_out(a7_wr[278]), .rdlo_out(a7_wr[286]));
			radix2 #(.width(width)) rd_st6_279  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[279]), .rdlo_in(a6_wr[287]),  .coef_in(coef[448]), .rdup_out(a7_wr[279]), .rdlo_out(a7_wr[287]));
			radix2 #(.width(width)) rd_st6_288  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[288]), .rdlo_in(a6_wr[296]),  .coef_in(coef[0]), .rdup_out(a7_wr[288]), .rdlo_out(a7_wr[296]));
			radix2 #(.width(width)) rd_st6_289  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[289]), .rdlo_in(a6_wr[297]),  .coef_in(coef[64]), .rdup_out(a7_wr[289]), .rdlo_out(a7_wr[297]));
			radix2 #(.width(width)) rd_st6_290  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[290]), .rdlo_in(a6_wr[298]),  .coef_in(coef[128]), .rdup_out(a7_wr[290]), .rdlo_out(a7_wr[298]));
			radix2 #(.width(width)) rd_st6_291  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[291]), .rdlo_in(a6_wr[299]),  .coef_in(coef[192]), .rdup_out(a7_wr[291]), .rdlo_out(a7_wr[299]));
			radix2 #(.width(width)) rd_st6_292  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[292]), .rdlo_in(a6_wr[300]),  .coef_in(coef[256]), .rdup_out(a7_wr[292]), .rdlo_out(a7_wr[300]));
			radix2 #(.width(width)) rd_st6_293  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[293]), .rdlo_in(a6_wr[301]),  .coef_in(coef[320]), .rdup_out(a7_wr[293]), .rdlo_out(a7_wr[301]));
			radix2 #(.width(width)) rd_st6_294  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[294]), .rdlo_in(a6_wr[302]),  .coef_in(coef[384]), .rdup_out(a7_wr[294]), .rdlo_out(a7_wr[302]));
			radix2 #(.width(width)) rd_st6_295  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[295]), .rdlo_in(a6_wr[303]),  .coef_in(coef[448]), .rdup_out(a7_wr[295]), .rdlo_out(a7_wr[303]));
			radix2 #(.width(width)) rd_st6_304  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[304]), .rdlo_in(a6_wr[312]),  .coef_in(coef[0]), .rdup_out(a7_wr[304]), .rdlo_out(a7_wr[312]));
			radix2 #(.width(width)) rd_st6_305  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[305]), .rdlo_in(a6_wr[313]),  .coef_in(coef[64]), .rdup_out(a7_wr[305]), .rdlo_out(a7_wr[313]));
			radix2 #(.width(width)) rd_st6_306  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[306]), .rdlo_in(a6_wr[314]),  .coef_in(coef[128]), .rdup_out(a7_wr[306]), .rdlo_out(a7_wr[314]));
			radix2 #(.width(width)) rd_st6_307  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[307]), .rdlo_in(a6_wr[315]),  .coef_in(coef[192]), .rdup_out(a7_wr[307]), .rdlo_out(a7_wr[315]));
			radix2 #(.width(width)) rd_st6_308  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[308]), .rdlo_in(a6_wr[316]),  .coef_in(coef[256]), .rdup_out(a7_wr[308]), .rdlo_out(a7_wr[316]));
			radix2 #(.width(width)) rd_st6_309  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[309]), .rdlo_in(a6_wr[317]),  .coef_in(coef[320]), .rdup_out(a7_wr[309]), .rdlo_out(a7_wr[317]));
			radix2 #(.width(width)) rd_st6_310  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[310]), .rdlo_in(a6_wr[318]),  .coef_in(coef[384]), .rdup_out(a7_wr[310]), .rdlo_out(a7_wr[318]));
			radix2 #(.width(width)) rd_st6_311  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[311]), .rdlo_in(a6_wr[319]),  .coef_in(coef[448]), .rdup_out(a7_wr[311]), .rdlo_out(a7_wr[319]));
			radix2 #(.width(width)) rd_st6_320  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[320]), .rdlo_in(a6_wr[328]),  .coef_in(coef[0]), .rdup_out(a7_wr[320]), .rdlo_out(a7_wr[328]));
			radix2 #(.width(width)) rd_st6_321  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[321]), .rdlo_in(a6_wr[329]),  .coef_in(coef[64]), .rdup_out(a7_wr[321]), .rdlo_out(a7_wr[329]));
			radix2 #(.width(width)) rd_st6_322  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[322]), .rdlo_in(a6_wr[330]),  .coef_in(coef[128]), .rdup_out(a7_wr[322]), .rdlo_out(a7_wr[330]));
			radix2 #(.width(width)) rd_st6_323  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[323]), .rdlo_in(a6_wr[331]),  .coef_in(coef[192]), .rdup_out(a7_wr[323]), .rdlo_out(a7_wr[331]));
			radix2 #(.width(width)) rd_st6_324  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[324]), .rdlo_in(a6_wr[332]),  .coef_in(coef[256]), .rdup_out(a7_wr[324]), .rdlo_out(a7_wr[332]));
			radix2 #(.width(width)) rd_st6_325  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[325]), .rdlo_in(a6_wr[333]),  .coef_in(coef[320]), .rdup_out(a7_wr[325]), .rdlo_out(a7_wr[333]));
			radix2 #(.width(width)) rd_st6_326  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[326]), .rdlo_in(a6_wr[334]),  .coef_in(coef[384]), .rdup_out(a7_wr[326]), .rdlo_out(a7_wr[334]));
			radix2 #(.width(width)) rd_st6_327  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[327]), .rdlo_in(a6_wr[335]),  .coef_in(coef[448]), .rdup_out(a7_wr[327]), .rdlo_out(a7_wr[335]));
			radix2 #(.width(width)) rd_st6_336  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[336]), .rdlo_in(a6_wr[344]),  .coef_in(coef[0]), .rdup_out(a7_wr[336]), .rdlo_out(a7_wr[344]));
			radix2 #(.width(width)) rd_st6_337  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[337]), .rdlo_in(a6_wr[345]),  .coef_in(coef[64]), .rdup_out(a7_wr[337]), .rdlo_out(a7_wr[345]));
			radix2 #(.width(width)) rd_st6_338  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[338]), .rdlo_in(a6_wr[346]),  .coef_in(coef[128]), .rdup_out(a7_wr[338]), .rdlo_out(a7_wr[346]));
			radix2 #(.width(width)) rd_st6_339  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[339]), .rdlo_in(a6_wr[347]),  .coef_in(coef[192]), .rdup_out(a7_wr[339]), .rdlo_out(a7_wr[347]));
			radix2 #(.width(width)) rd_st6_340  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[340]), .rdlo_in(a6_wr[348]),  .coef_in(coef[256]), .rdup_out(a7_wr[340]), .rdlo_out(a7_wr[348]));
			radix2 #(.width(width)) rd_st6_341  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[341]), .rdlo_in(a6_wr[349]),  .coef_in(coef[320]), .rdup_out(a7_wr[341]), .rdlo_out(a7_wr[349]));
			radix2 #(.width(width)) rd_st6_342  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[342]), .rdlo_in(a6_wr[350]),  .coef_in(coef[384]), .rdup_out(a7_wr[342]), .rdlo_out(a7_wr[350]));
			radix2 #(.width(width)) rd_st6_343  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[343]), .rdlo_in(a6_wr[351]),  .coef_in(coef[448]), .rdup_out(a7_wr[343]), .rdlo_out(a7_wr[351]));
			radix2 #(.width(width)) rd_st6_352  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[352]), .rdlo_in(a6_wr[360]),  .coef_in(coef[0]), .rdup_out(a7_wr[352]), .rdlo_out(a7_wr[360]));
			radix2 #(.width(width)) rd_st6_353  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[353]), .rdlo_in(a6_wr[361]),  .coef_in(coef[64]), .rdup_out(a7_wr[353]), .rdlo_out(a7_wr[361]));
			radix2 #(.width(width)) rd_st6_354  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[354]), .rdlo_in(a6_wr[362]),  .coef_in(coef[128]), .rdup_out(a7_wr[354]), .rdlo_out(a7_wr[362]));
			radix2 #(.width(width)) rd_st6_355  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[355]), .rdlo_in(a6_wr[363]),  .coef_in(coef[192]), .rdup_out(a7_wr[355]), .rdlo_out(a7_wr[363]));
			radix2 #(.width(width)) rd_st6_356  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[356]), .rdlo_in(a6_wr[364]),  .coef_in(coef[256]), .rdup_out(a7_wr[356]), .rdlo_out(a7_wr[364]));
			radix2 #(.width(width)) rd_st6_357  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[357]), .rdlo_in(a6_wr[365]),  .coef_in(coef[320]), .rdup_out(a7_wr[357]), .rdlo_out(a7_wr[365]));
			radix2 #(.width(width)) rd_st6_358  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[358]), .rdlo_in(a6_wr[366]),  .coef_in(coef[384]), .rdup_out(a7_wr[358]), .rdlo_out(a7_wr[366]));
			radix2 #(.width(width)) rd_st6_359  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[359]), .rdlo_in(a6_wr[367]),  .coef_in(coef[448]), .rdup_out(a7_wr[359]), .rdlo_out(a7_wr[367]));
			radix2 #(.width(width)) rd_st6_368  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[368]), .rdlo_in(a6_wr[376]),  .coef_in(coef[0]), .rdup_out(a7_wr[368]), .rdlo_out(a7_wr[376]));
			radix2 #(.width(width)) rd_st6_369  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[369]), .rdlo_in(a6_wr[377]),  .coef_in(coef[64]), .rdup_out(a7_wr[369]), .rdlo_out(a7_wr[377]));
			radix2 #(.width(width)) rd_st6_370  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[370]), .rdlo_in(a6_wr[378]),  .coef_in(coef[128]), .rdup_out(a7_wr[370]), .rdlo_out(a7_wr[378]));
			radix2 #(.width(width)) rd_st6_371  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[371]), .rdlo_in(a6_wr[379]),  .coef_in(coef[192]), .rdup_out(a7_wr[371]), .rdlo_out(a7_wr[379]));
			radix2 #(.width(width)) rd_st6_372  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[372]), .rdlo_in(a6_wr[380]),  .coef_in(coef[256]), .rdup_out(a7_wr[372]), .rdlo_out(a7_wr[380]));
			radix2 #(.width(width)) rd_st6_373  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[373]), .rdlo_in(a6_wr[381]),  .coef_in(coef[320]), .rdup_out(a7_wr[373]), .rdlo_out(a7_wr[381]));
			radix2 #(.width(width)) rd_st6_374  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[374]), .rdlo_in(a6_wr[382]),  .coef_in(coef[384]), .rdup_out(a7_wr[374]), .rdlo_out(a7_wr[382]));
			radix2 #(.width(width)) rd_st6_375  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[375]), .rdlo_in(a6_wr[383]),  .coef_in(coef[448]), .rdup_out(a7_wr[375]), .rdlo_out(a7_wr[383]));
			radix2 #(.width(width)) rd_st6_384  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[384]), .rdlo_in(a6_wr[392]),  .coef_in(coef[0]), .rdup_out(a7_wr[384]), .rdlo_out(a7_wr[392]));
			radix2 #(.width(width)) rd_st6_385  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[385]), .rdlo_in(a6_wr[393]),  .coef_in(coef[64]), .rdup_out(a7_wr[385]), .rdlo_out(a7_wr[393]));
			radix2 #(.width(width)) rd_st6_386  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[386]), .rdlo_in(a6_wr[394]),  .coef_in(coef[128]), .rdup_out(a7_wr[386]), .rdlo_out(a7_wr[394]));
			radix2 #(.width(width)) rd_st6_387  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[387]), .rdlo_in(a6_wr[395]),  .coef_in(coef[192]), .rdup_out(a7_wr[387]), .rdlo_out(a7_wr[395]));
			radix2 #(.width(width)) rd_st6_388  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[388]), .rdlo_in(a6_wr[396]),  .coef_in(coef[256]), .rdup_out(a7_wr[388]), .rdlo_out(a7_wr[396]));
			radix2 #(.width(width)) rd_st6_389  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[389]), .rdlo_in(a6_wr[397]),  .coef_in(coef[320]), .rdup_out(a7_wr[389]), .rdlo_out(a7_wr[397]));
			radix2 #(.width(width)) rd_st6_390  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[390]), .rdlo_in(a6_wr[398]),  .coef_in(coef[384]), .rdup_out(a7_wr[390]), .rdlo_out(a7_wr[398]));
			radix2 #(.width(width)) rd_st6_391  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[391]), .rdlo_in(a6_wr[399]),  .coef_in(coef[448]), .rdup_out(a7_wr[391]), .rdlo_out(a7_wr[399]));
			radix2 #(.width(width)) rd_st6_400  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[400]), .rdlo_in(a6_wr[408]),  .coef_in(coef[0]), .rdup_out(a7_wr[400]), .rdlo_out(a7_wr[408]));
			radix2 #(.width(width)) rd_st6_401  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[401]), .rdlo_in(a6_wr[409]),  .coef_in(coef[64]), .rdup_out(a7_wr[401]), .rdlo_out(a7_wr[409]));
			radix2 #(.width(width)) rd_st6_402  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[402]), .rdlo_in(a6_wr[410]),  .coef_in(coef[128]), .rdup_out(a7_wr[402]), .rdlo_out(a7_wr[410]));
			radix2 #(.width(width)) rd_st6_403  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[403]), .rdlo_in(a6_wr[411]),  .coef_in(coef[192]), .rdup_out(a7_wr[403]), .rdlo_out(a7_wr[411]));
			radix2 #(.width(width)) rd_st6_404  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[404]), .rdlo_in(a6_wr[412]),  .coef_in(coef[256]), .rdup_out(a7_wr[404]), .rdlo_out(a7_wr[412]));
			radix2 #(.width(width)) rd_st6_405  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[405]), .rdlo_in(a6_wr[413]),  .coef_in(coef[320]), .rdup_out(a7_wr[405]), .rdlo_out(a7_wr[413]));
			radix2 #(.width(width)) rd_st6_406  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[406]), .rdlo_in(a6_wr[414]),  .coef_in(coef[384]), .rdup_out(a7_wr[406]), .rdlo_out(a7_wr[414]));
			radix2 #(.width(width)) rd_st6_407  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[407]), .rdlo_in(a6_wr[415]),  .coef_in(coef[448]), .rdup_out(a7_wr[407]), .rdlo_out(a7_wr[415]));
			radix2 #(.width(width)) rd_st6_416  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[416]), .rdlo_in(a6_wr[424]),  .coef_in(coef[0]), .rdup_out(a7_wr[416]), .rdlo_out(a7_wr[424]));
			radix2 #(.width(width)) rd_st6_417  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[417]), .rdlo_in(a6_wr[425]),  .coef_in(coef[64]), .rdup_out(a7_wr[417]), .rdlo_out(a7_wr[425]));
			radix2 #(.width(width)) rd_st6_418  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[418]), .rdlo_in(a6_wr[426]),  .coef_in(coef[128]), .rdup_out(a7_wr[418]), .rdlo_out(a7_wr[426]));
			radix2 #(.width(width)) rd_st6_419  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[419]), .rdlo_in(a6_wr[427]),  .coef_in(coef[192]), .rdup_out(a7_wr[419]), .rdlo_out(a7_wr[427]));
			radix2 #(.width(width)) rd_st6_420  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[420]), .rdlo_in(a6_wr[428]),  .coef_in(coef[256]), .rdup_out(a7_wr[420]), .rdlo_out(a7_wr[428]));
			radix2 #(.width(width)) rd_st6_421  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[421]), .rdlo_in(a6_wr[429]),  .coef_in(coef[320]), .rdup_out(a7_wr[421]), .rdlo_out(a7_wr[429]));
			radix2 #(.width(width)) rd_st6_422  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[422]), .rdlo_in(a6_wr[430]),  .coef_in(coef[384]), .rdup_out(a7_wr[422]), .rdlo_out(a7_wr[430]));
			radix2 #(.width(width)) rd_st6_423  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[423]), .rdlo_in(a6_wr[431]),  .coef_in(coef[448]), .rdup_out(a7_wr[423]), .rdlo_out(a7_wr[431]));
			radix2 #(.width(width)) rd_st6_432  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[432]), .rdlo_in(a6_wr[440]),  .coef_in(coef[0]), .rdup_out(a7_wr[432]), .rdlo_out(a7_wr[440]));
			radix2 #(.width(width)) rd_st6_433  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[433]), .rdlo_in(a6_wr[441]),  .coef_in(coef[64]), .rdup_out(a7_wr[433]), .rdlo_out(a7_wr[441]));
			radix2 #(.width(width)) rd_st6_434  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[434]), .rdlo_in(a6_wr[442]),  .coef_in(coef[128]), .rdup_out(a7_wr[434]), .rdlo_out(a7_wr[442]));
			radix2 #(.width(width)) rd_st6_435  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[435]), .rdlo_in(a6_wr[443]),  .coef_in(coef[192]), .rdup_out(a7_wr[435]), .rdlo_out(a7_wr[443]));
			radix2 #(.width(width)) rd_st6_436  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[436]), .rdlo_in(a6_wr[444]),  .coef_in(coef[256]), .rdup_out(a7_wr[436]), .rdlo_out(a7_wr[444]));
			radix2 #(.width(width)) rd_st6_437  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[437]), .rdlo_in(a6_wr[445]),  .coef_in(coef[320]), .rdup_out(a7_wr[437]), .rdlo_out(a7_wr[445]));
			radix2 #(.width(width)) rd_st6_438  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[438]), .rdlo_in(a6_wr[446]),  .coef_in(coef[384]), .rdup_out(a7_wr[438]), .rdlo_out(a7_wr[446]));
			radix2 #(.width(width)) rd_st6_439  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[439]), .rdlo_in(a6_wr[447]),  .coef_in(coef[448]), .rdup_out(a7_wr[439]), .rdlo_out(a7_wr[447]));
			radix2 #(.width(width)) rd_st6_448  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[448]), .rdlo_in(a6_wr[456]),  .coef_in(coef[0]), .rdup_out(a7_wr[448]), .rdlo_out(a7_wr[456]));
			radix2 #(.width(width)) rd_st6_449  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[449]), .rdlo_in(a6_wr[457]),  .coef_in(coef[64]), .rdup_out(a7_wr[449]), .rdlo_out(a7_wr[457]));
			radix2 #(.width(width)) rd_st6_450  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[450]), .rdlo_in(a6_wr[458]),  .coef_in(coef[128]), .rdup_out(a7_wr[450]), .rdlo_out(a7_wr[458]));
			radix2 #(.width(width)) rd_st6_451  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[451]), .rdlo_in(a6_wr[459]),  .coef_in(coef[192]), .rdup_out(a7_wr[451]), .rdlo_out(a7_wr[459]));
			radix2 #(.width(width)) rd_st6_452  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[452]), .rdlo_in(a6_wr[460]),  .coef_in(coef[256]), .rdup_out(a7_wr[452]), .rdlo_out(a7_wr[460]));
			radix2 #(.width(width)) rd_st6_453  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[453]), .rdlo_in(a6_wr[461]),  .coef_in(coef[320]), .rdup_out(a7_wr[453]), .rdlo_out(a7_wr[461]));
			radix2 #(.width(width)) rd_st6_454  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[454]), .rdlo_in(a6_wr[462]),  .coef_in(coef[384]), .rdup_out(a7_wr[454]), .rdlo_out(a7_wr[462]));
			radix2 #(.width(width)) rd_st6_455  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[455]), .rdlo_in(a6_wr[463]),  .coef_in(coef[448]), .rdup_out(a7_wr[455]), .rdlo_out(a7_wr[463]));
			radix2 #(.width(width)) rd_st6_464  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[464]), .rdlo_in(a6_wr[472]),  .coef_in(coef[0]), .rdup_out(a7_wr[464]), .rdlo_out(a7_wr[472]));
			radix2 #(.width(width)) rd_st6_465  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[465]), .rdlo_in(a6_wr[473]),  .coef_in(coef[64]), .rdup_out(a7_wr[465]), .rdlo_out(a7_wr[473]));
			radix2 #(.width(width)) rd_st6_466  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[466]), .rdlo_in(a6_wr[474]),  .coef_in(coef[128]), .rdup_out(a7_wr[466]), .rdlo_out(a7_wr[474]));
			radix2 #(.width(width)) rd_st6_467  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[467]), .rdlo_in(a6_wr[475]),  .coef_in(coef[192]), .rdup_out(a7_wr[467]), .rdlo_out(a7_wr[475]));
			radix2 #(.width(width)) rd_st6_468  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[468]), .rdlo_in(a6_wr[476]),  .coef_in(coef[256]), .rdup_out(a7_wr[468]), .rdlo_out(a7_wr[476]));
			radix2 #(.width(width)) rd_st6_469  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[469]), .rdlo_in(a6_wr[477]),  .coef_in(coef[320]), .rdup_out(a7_wr[469]), .rdlo_out(a7_wr[477]));
			radix2 #(.width(width)) rd_st6_470  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[470]), .rdlo_in(a6_wr[478]),  .coef_in(coef[384]), .rdup_out(a7_wr[470]), .rdlo_out(a7_wr[478]));
			radix2 #(.width(width)) rd_st6_471  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[471]), .rdlo_in(a6_wr[479]),  .coef_in(coef[448]), .rdup_out(a7_wr[471]), .rdlo_out(a7_wr[479]));
			radix2 #(.width(width)) rd_st6_480  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[480]), .rdlo_in(a6_wr[488]),  .coef_in(coef[0]), .rdup_out(a7_wr[480]), .rdlo_out(a7_wr[488]));
			radix2 #(.width(width)) rd_st6_481  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[481]), .rdlo_in(a6_wr[489]),  .coef_in(coef[64]), .rdup_out(a7_wr[481]), .rdlo_out(a7_wr[489]));
			radix2 #(.width(width)) rd_st6_482  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[482]), .rdlo_in(a6_wr[490]),  .coef_in(coef[128]), .rdup_out(a7_wr[482]), .rdlo_out(a7_wr[490]));
			radix2 #(.width(width)) rd_st6_483  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[483]), .rdlo_in(a6_wr[491]),  .coef_in(coef[192]), .rdup_out(a7_wr[483]), .rdlo_out(a7_wr[491]));
			radix2 #(.width(width)) rd_st6_484  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[484]), .rdlo_in(a6_wr[492]),  .coef_in(coef[256]), .rdup_out(a7_wr[484]), .rdlo_out(a7_wr[492]));
			radix2 #(.width(width)) rd_st6_485  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[485]), .rdlo_in(a6_wr[493]),  .coef_in(coef[320]), .rdup_out(a7_wr[485]), .rdlo_out(a7_wr[493]));
			radix2 #(.width(width)) rd_st6_486  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[486]), .rdlo_in(a6_wr[494]),  .coef_in(coef[384]), .rdup_out(a7_wr[486]), .rdlo_out(a7_wr[494]));
			radix2 #(.width(width)) rd_st6_487  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[487]), .rdlo_in(a6_wr[495]),  .coef_in(coef[448]), .rdup_out(a7_wr[487]), .rdlo_out(a7_wr[495]));
			radix2 #(.width(width)) rd_st6_496  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[496]), .rdlo_in(a6_wr[504]),  .coef_in(coef[0]), .rdup_out(a7_wr[496]), .rdlo_out(a7_wr[504]));
			radix2 #(.width(width)) rd_st6_497  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[497]), .rdlo_in(a6_wr[505]),  .coef_in(coef[64]), .rdup_out(a7_wr[497]), .rdlo_out(a7_wr[505]));
			radix2 #(.width(width)) rd_st6_498  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[498]), .rdlo_in(a6_wr[506]),  .coef_in(coef[128]), .rdup_out(a7_wr[498]), .rdlo_out(a7_wr[506]));
			radix2 #(.width(width)) rd_st6_499  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[499]), .rdlo_in(a6_wr[507]),  .coef_in(coef[192]), .rdup_out(a7_wr[499]), .rdlo_out(a7_wr[507]));
			radix2 #(.width(width)) rd_st6_500  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[500]), .rdlo_in(a6_wr[508]),  .coef_in(coef[256]), .rdup_out(a7_wr[500]), .rdlo_out(a7_wr[508]));
			radix2 #(.width(width)) rd_st6_501  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[501]), .rdlo_in(a6_wr[509]),  .coef_in(coef[320]), .rdup_out(a7_wr[501]), .rdlo_out(a7_wr[509]));
			radix2 #(.width(width)) rd_st6_502  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[502]), .rdlo_in(a6_wr[510]),  .coef_in(coef[384]), .rdup_out(a7_wr[502]), .rdlo_out(a7_wr[510]));
			radix2 #(.width(width)) rd_st6_503  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[503]), .rdlo_in(a6_wr[511]),  .coef_in(coef[448]), .rdup_out(a7_wr[503]), .rdlo_out(a7_wr[511]));
			radix2 #(.width(width)) rd_st6_512  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[512]), .rdlo_in(a6_wr[520]),  .coef_in(coef[0]), .rdup_out(a7_wr[512]), .rdlo_out(a7_wr[520]));
			radix2 #(.width(width)) rd_st6_513  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[513]), .rdlo_in(a6_wr[521]),  .coef_in(coef[64]), .rdup_out(a7_wr[513]), .rdlo_out(a7_wr[521]));
			radix2 #(.width(width)) rd_st6_514  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[514]), .rdlo_in(a6_wr[522]),  .coef_in(coef[128]), .rdup_out(a7_wr[514]), .rdlo_out(a7_wr[522]));
			radix2 #(.width(width)) rd_st6_515  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[515]), .rdlo_in(a6_wr[523]),  .coef_in(coef[192]), .rdup_out(a7_wr[515]), .rdlo_out(a7_wr[523]));
			radix2 #(.width(width)) rd_st6_516  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[516]), .rdlo_in(a6_wr[524]),  .coef_in(coef[256]), .rdup_out(a7_wr[516]), .rdlo_out(a7_wr[524]));
			radix2 #(.width(width)) rd_st6_517  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[517]), .rdlo_in(a6_wr[525]),  .coef_in(coef[320]), .rdup_out(a7_wr[517]), .rdlo_out(a7_wr[525]));
			radix2 #(.width(width)) rd_st6_518  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[518]), .rdlo_in(a6_wr[526]),  .coef_in(coef[384]), .rdup_out(a7_wr[518]), .rdlo_out(a7_wr[526]));
			radix2 #(.width(width)) rd_st6_519  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[519]), .rdlo_in(a6_wr[527]),  .coef_in(coef[448]), .rdup_out(a7_wr[519]), .rdlo_out(a7_wr[527]));
			radix2 #(.width(width)) rd_st6_528  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[528]), .rdlo_in(a6_wr[536]),  .coef_in(coef[0]), .rdup_out(a7_wr[528]), .rdlo_out(a7_wr[536]));
			radix2 #(.width(width)) rd_st6_529  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[529]), .rdlo_in(a6_wr[537]),  .coef_in(coef[64]), .rdup_out(a7_wr[529]), .rdlo_out(a7_wr[537]));
			radix2 #(.width(width)) rd_st6_530  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[530]), .rdlo_in(a6_wr[538]),  .coef_in(coef[128]), .rdup_out(a7_wr[530]), .rdlo_out(a7_wr[538]));
			radix2 #(.width(width)) rd_st6_531  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[531]), .rdlo_in(a6_wr[539]),  .coef_in(coef[192]), .rdup_out(a7_wr[531]), .rdlo_out(a7_wr[539]));
			radix2 #(.width(width)) rd_st6_532  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[532]), .rdlo_in(a6_wr[540]),  .coef_in(coef[256]), .rdup_out(a7_wr[532]), .rdlo_out(a7_wr[540]));
			radix2 #(.width(width)) rd_st6_533  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[533]), .rdlo_in(a6_wr[541]),  .coef_in(coef[320]), .rdup_out(a7_wr[533]), .rdlo_out(a7_wr[541]));
			radix2 #(.width(width)) rd_st6_534  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[534]), .rdlo_in(a6_wr[542]),  .coef_in(coef[384]), .rdup_out(a7_wr[534]), .rdlo_out(a7_wr[542]));
			radix2 #(.width(width)) rd_st6_535  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[535]), .rdlo_in(a6_wr[543]),  .coef_in(coef[448]), .rdup_out(a7_wr[535]), .rdlo_out(a7_wr[543]));
			radix2 #(.width(width)) rd_st6_544  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[544]), .rdlo_in(a6_wr[552]),  .coef_in(coef[0]), .rdup_out(a7_wr[544]), .rdlo_out(a7_wr[552]));
			radix2 #(.width(width)) rd_st6_545  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[545]), .rdlo_in(a6_wr[553]),  .coef_in(coef[64]), .rdup_out(a7_wr[545]), .rdlo_out(a7_wr[553]));
			radix2 #(.width(width)) rd_st6_546  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[546]), .rdlo_in(a6_wr[554]),  .coef_in(coef[128]), .rdup_out(a7_wr[546]), .rdlo_out(a7_wr[554]));
			radix2 #(.width(width)) rd_st6_547  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[547]), .rdlo_in(a6_wr[555]),  .coef_in(coef[192]), .rdup_out(a7_wr[547]), .rdlo_out(a7_wr[555]));
			radix2 #(.width(width)) rd_st6_548  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[548]), .rdlo_in(a6_wr[556]),  .coef_in(coef[256]), .rdup_out(a7_wr[548]), .rdlo_out(a7_wr[556]));
			radix2 #(.width(width)) rd_st6_549  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[549]), .rdlo_in(a6_wr[557]),  .coef_in(coef[320]), .rdup_out(a7_wr[549]), .rdlo_out(a7_wr[557]));
			radix2 #(.width(width)) rd_st6_550  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[550]), .rdlo_in(a6_wr[558]),  .coef_in(coef[384]), .rdup_out(a7_wr[550]), .rdlo_out(a7_wr[558]));
			radix2 #(.width(width)) rd_st6_551  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[551]), .rdlo_in(a6_wr[559]),  .coef_in(coef[448]), .rdup_out(a7_wr[551]), .rdlo_out(a7_wr[559]));
			radix2 #(.width(width)) rd_st6_560  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[560]), .rdlo_in(a6_wr[568]),  .coef_in(coef[0]), .rdup_out(a7_wr[560]), .rdlo_out(a7_wr[568]));
			radix2 #(.width(width)) rd_st6_561  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[561]), .rdlo_in(a6_wr[569]),  .coef_in(coef[64]), .rdup_out(a7_wr[561]), .rdlo_out(a7_wr[569]));
			radix2 #(.width(width)) rd_st6_562  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[562]), .rdlo_in(a6_wr[570]),  .coef_in(coef[128]), .rdup_out(a7_wr[562]), .rdlo_out(a7_wr[570]));
			radix2 #(.width(width)) rd_st6_563  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[563]), .rdlo_in(a6_wr[571]),  .coef_in(coef[192]), .rdup_out(a7_wr[563]), .rdlo_out(a7_wr[571]));
			radix2 #(.width(width)) rd_st6_564  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[564]), .rdlo_in(a6_wr[572]),  .coef_in(coef[256]), .rdup_out(a7_wr[564]), .rdlo_out(a7_wr[572]));
			radix2 #(.width(width)) rd_st6_565  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[565]), .rdlo_in(a6_wr[573]),  .coef_in(coef[320]), .rdup_out(a7_wr[565]), .rdlo_out(a7_wr[573]));
			radix2 #(.width(width)) rd_st6_566  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[566]), .rdlo_in(a6_wr[574]),  .coef_in(coef[384]), .rdup_out(a7_wr[566]), .rdlo_out(a7_wr[574]));
			radix2 #(.width(width)) rd_st6_567  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[567]), .rdlo_in(a6_wr[575]),  .coef_in(coef[448]), .rdup_out(a7_wr[567]), .rdlo_out(a7_wr[575]));
			radix2 #(.width(width)) rd_st6_576  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[576]), .rdlo_in(a6_wr[584]),  .coef_in(coef[0]), .rdup_out(a7_wr[576]), .rdlo_out(a7_wr[584]));
			radix2 #(.width(width)) rd_st6_577  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[577]), .rdlo_in(a6_wr[585]),  .coef_in(coef[64]), .rdup_out(a7_wr[577]), .rdlo_out(a7_wr[585]));
			radix2 #(.width(width)) rd_st6_578  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[578]), .rdlo_in(a6_wr[586]),  .coef_in(coef[128]), .rdup_out(a7_wr[578]), .rdlo_out(a7_wr[586]));
			radix2 #(.width(width)) rd_st6_579  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[579]), .rdlo_in(a6_wr[587]),  .coef_in(coef[192]), .rdup_out(a7_wr[579]), .rdlo_out(a7_wr[587]));
			radix2 #(.width(width)) rd_st6_580  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[580]), .rdlo_in(a6_wr[588]),  .coef_in(coef[256]), .rdup_out(a7_wr[580]), .rdlo_out(a7_wr[588]));
			radix2 #(.width(width)) rd_st6_581  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[581]), .rdlo_in(a6_wr[589]),  .coef_in(coef[320]), .rdup_out(a7_wr[581]), .rdlo_out(a7_wr[589]));
			radix2 #(.width(width)) rd_st6_582  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[582]), .rdlo_in(a6_wr[590]),  .coef_in(coef[384]), .rdup_out(a7_wr[582]), .rdlo_out(a7_wr[590]));
			radix2 #(.width(width)) rd_st6_583  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[583]), .rdlo_in(a6_wr[591]),  .coef_in(coef[448]), .rdup_out(a7_wr[583]), .rdlo_out(a7_wr[591]));
			radix2 #(.width(width)) rd_st6_592  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[592]), .rdlo_in(a6_wr[600]),  .coef_in(coef[0]), .rdup_out(a7_wr[592]), .rdlo_out(a7_wr[600]));
			radix2 #(.width(width)) rd_st6_593  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[593]), .rdlo_in(a6_wr[601]),  .coef_in(coef[64]), .rdup_out(a7_wr[593]), .rdlo_out(a7_wr[601]));
			radix2 #(.width(width)) rd_st6_594  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[594]), .rdlo_in(a6_wr[602]),  .coef_in(coef[128]), .rdup_out(a7_wr[594]), .rdlo_out(a7_wr[602]));
			radix2 #(.width(width)) rd_st6_595  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[595]), .rdlo_in(a6_wr[603]),  .coef_in(coef[192]), .rdup_out(a7_wr[595]), .rdlo_out(a7_wr[603]));
			radix2 #(.width(width)) rd_st6_596  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[596]), .rdlo_in(a6_wr[604]),  .coef_in(coef[256]), .rdup_out(a7_wr[596]), .rdlo_out(a7_wr[604]));
			radix2 #(.width(width)) rd_st6_597  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[597]), .rdlo_in(a6_wr[605]),  .coef_in(coef[320]), .rdup_out(a7_wr[597]), .rdlo_out(a7_wr[605]));
			radix2 #(.width(width)) rd_st6_598  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[598]), .rdlo_in(a6_wr[606]),  .coef_in(coef[384]), .rdup_out(a7_wr[598]), .rdlo_out(a7_wr[606]));
			radix2 #(.width(width)) rd_st6_599  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[599]), .rdlo_in(a6_wr[607]),  .coef_in(coef[448]), .rdup_out(a7_wr[599]), .rdlo_out(a7_wr[607]));
			radix2 #(.width(width)) rd_st6_608  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[608]), .rdlo_in(a6_wr[616]),  .coef_in(coef[0]), .rdup_out(a7_wr[608]), .rdlo_out(a7_wr[616]));
			radix2 #(.width(width)) rd_st6_609  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[609]), .rdlo_in(a6_wr[617]),  .coef_in(coef[64]), .rdup_out(a7_wr[609]), .rdlo_out(a7_wr[617]));
			radix2 #(.width(width)) rd_st6_610  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[610]), .rdlo_in(a6_wr[618]),  .coef_in(coef[128]), .rdup_out(a7_wr[610]), .rdlo_out(a7_wr[618]));
			radix2 #(.width(width)) rd_st6_611  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[611]), .rdlo_in(a6_wr[619]),  .coef_in(coef[192]), .rdup_out(a7_wr[611]), .rdlo_out(a7_wr[619]));
			radix2 #(.width(width)) rd_st6_612  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[612]), .rdlo_in(a6_wr[620]),  .coef_in(coef[256]), .rdup_out(a7_wr[612]), .rdlo_out(a7_wr[620]));
			radix2 #(.width(width)) rd_st6_613  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[613]), .rdlo_in(a6_wr[621]),  .coef_in(coef[320]), .rdup_out(a7_wr[613]), .rdlo_out(a7_wr[621]));
			radix2 #(.width(width)) rd_st6_614  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[614]), .rdlo_in(a6_wr[622]),  .coef_in(coef[384]), .rdup_out(a7_wr[614]), .rdlo_out(a7_wr[622]));
			radix2 #(.width(width)) rd_st6_615  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[615]), .rdlo_in(a6_wr[623]),  .coef_in(coef[448]), .rdup_out(a7_wr[615]), .rdlo_out(a7_wr[623]));
			radix2 #(.width(width)) rd_st6_624  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[624]), .rdlo_in(a6_wr[632]),  .coef_in(coef[0]), .rdup_out(a7_wr[624]), .rdlo_out(a7_wr[632]));
			radix2 #(.width(width)) rd_st6_625  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[625]), .rdlo_in(a6_wr[633]),  .coef_in(coef[64]), .rdup_out(a7_wr[625]), .rdlo_out(a7_wr[633]));
			radix2 #(.width(width)) rd_st6_626  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[626]), .rdlo_in(a6_wr[634]),  .coef_in(coef[128]), .rdup_out(a7_wr[626]), .rdlo_out(a7_wr[634]));
			radix2 #(.width(width)) rd_st6_627  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[627]), .rdlo_in(a6_wr[635]),  .coef_in(coef[192]), .rdup_out(a7_wr[627]), .rdlo_out(a7_wr[635]));
			radix2 #(.width(width)) rd_st6_628  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[628]), .rdlo_in(a6_wr[636]),  .coef_in(coef[256]), .rdup_out(a7_wr[628]), .rdlo_out(a7_wr[636]));
			radix2 #(.width(width)) rd_st6_629  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[629]), .rdlo_in(a6_wr[637]),  .coef_in(coef[320]), .rdup_out(a7_wr[629]), .rdlo_out(a7_wr[637]));
			radix2 #(.width(width)) rd_st6_630  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[630]), .rdlo_in(a6_wr[638]),  .coef_in(coef[384]), .rdup_out(a7_wr[630]), .rdlo_out(a7_wr[638]));
			radix2 #(.width(width)) rd_st6_631  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[631]), .rdlo_in(a6_wr[639]),  .coef_in(coef[448]), .rdup_out(a7_wr[631]), .rdlo_out(a7_wr[639]));
			radix2 #(.width(width)) rd_st6_640  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[640]), .rdlo_in(a6_wr[648]),  .coef_in(coef[0]), .rdup_out(a7_wr[640]), .rdlo_out(a7_wr[648]));
			radix2 #(.width(width)) rd_st6_641  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[641]), .rdlo_in(a6_wr[649]),  .coef_in(coef[64]), .rdup_out(a7_wr[641]), .rdlo_out(a7_wr[649]));
			radix2 #(.width(width)) rd_st6_642  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[642]), .rdlo_in(a6_wr[650]),  .coef_in(coef[128]), .rdup_out(a7_wr[642]), .rdlo_out(a7_wr[650]));
			radix2 #(.width(width)) rd_st6_643  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[643]), .rdlo_in(a6_wr[651]),  .coef_in(coef[192]), .rdup_out(a7_wr[643]), .rdlo_out(a7_wr[651]));
			radix2 #(.width(width)) rd_st6_644  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[644]), .rdlo_in(a6_wr[652]),  .coef_in(coef[256]), .rdup_out(a7_wr[644]), .rdlo_out(a7_wr[652]));
			radix2 #(.width(width)) rd_st6_645  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[645]), .rdlo_in(a6_wr[653]),  .coef_in(coef[320]), .rdup_out(a7_wr[645]), .rdlo_out(a7_wr[653]));
			radix2 #(.width(width)) rd_st6_646  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[646]), .rdlo_in(a6_wr[654]),  .coef_in(coef[384]), .rdup_out(a7_wr[646]), .rdlo_out(a7_wr[654]));
			radix2 #(.width(width)) rd_st6_647  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[647]), .rdlo_in(a6_wr[655]),  .coef_in(coef[448]), .rdup_out(a7_wr[647]), .rdlo_out(a7_wr[655]));
			radix2 #(.width(width)) rd_st6_656  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[656]), .rdlo_in(a6_wr[664]),  .coef_in(coef[0]), .rdup_out(a7_wr[656]), .rdlo_out(a7_wr[664]));
			radix2 #(.width(width)) rd_st6_657  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[657]), .rdlo_in(a6_wr[665]),  .coef_in(coef[64]), .rdup_out(a7_wr[657]), .rdlo_out(a7_wr[665]));
			radix2 #(.width(width)) rd_st6_658  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[658]), .rdlo_in(a6_wr[666]),  .coef_in(coef[128]), .rdup_out(a7_wr[658]), .rdlo_out(a7_wr[666]));
			radix2 #(.width(width)) rd_st6_659  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[659]), .rdlo_in(a6_wr[667]),  .coef_in(coef[192]), .rdup_out(a7_wr[659]), .rdlo_out(a7_wr[667]));
			radix2 #(.width(width)) rd_st6_660  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[660]), .rdlo_in(a6_wr[668]),  .coef_in(coef[256]), .rdup_out(a7_wr[660]), .rdlo_out(a7_wr[668]));
			radix2 #(.width(width)) rd_st6_661  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[661]), .rdlo_in(a6_wr[669]),  .coef_in(coef[320]), .rdup_out(a7_wr[661]), .rdlo_out(a7_wr[669]));
			radix2 #(.width(width)) rd_st6_662  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[662]), .rdlo_in(a6_wr[670]),  .coef_in(coef[384]), .rdup_out(a7_wr[662]), .rdlo_out(a7_wr[670]));
			radix2 #(.width(width)) rd_st6_663  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[663]), .rdlo_in(a6_wr[671]),  .coef_in(coef[448]), .rdup_out(a7_wr[663]), .rdlo_out(a7_wr[671]));
			radix2 #(.width(width)) rd_st6_672  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[672]), .rdlo_in(a6_wr[680]),  .coef_in(coef[0]), .rdup_out(a7_wr[672]), .rdlo_out(a7_wr[680]));
			radix2 #(.width(width)) rd_st6_673  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[673]), .rdlo_in(a6_wr[681]),  .coef_in(coef[64]), .rdup_out(a7_wr[673]), .rdlo_out(a7_wr[681]));
			radix2 #(.width(width)) rd_st6_674  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[674]), .rdlo_in(a6_wr[682]),  .coef_in(coef[128]), .rdup_out(a7_wr[674]), .rdlo_out(a7_wr[682]));
			radix2 #(.width(width)) rd_st6_675  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[675]), .rdlo_in(a6_wr[683]),  .coef_in(coef[192]), .rdup_out(a7_wr[675]), .rdlo_out(a7_wr[683]));
			radix2 #(.width(width)) rd_st6_676  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[676]), .rdlo_in(a6_wr[684]),  .coef_in(coef[256]), .rdup_out(a7_wr[676]), .rdlo_out(a7_wr[684]));
			radix2 #(.width(width)) rd_st6_677  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[677]), .rdlo_in(a6_wr[685]),  .coef_in(coef[320]), .rdup_out(a7_wr[677]), .rdlo_out(a7_wr[685]));
			radix2 #(.width(width)) rd_st6_678  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[678]), .rdlo_in(a6_wr[686]),  .coef_in(coef[384]), .rdup_out(a7_wr[678]), .rdlo_out(a7_wr[686]));
			radix2 #(.width(width)) rd_st6_679  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[679]), .rdlo_in(a6_wr[687]),  .coef_in(coef[448]), .rdup_out(a7_wr[679]), .rdlo_out(a7_wr[687]));
			radix2 #(.width(width)) rd_st6_688  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[688]), .rdlo_in(a6_wr[696]),  .coef_in(coef[0]), .rdup_out(a7_wr[688]), .rdlo_out(a7_wr[696]));
			radix2 #(.width(width)) rd_st6_689  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[689]), .rdlo_in(a6_wr[697]),  .coef_in(coef[64]), .rdup_out(a7_wr[689]), .rdlo_out(a7_wr[697]));
			radix2 #(.width(width)) rd_st6_690  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[690]), .rdlo_in(a6_wr[698]),  .coef_in(coef[128]), .rdup_out(a7_wr[690]), .rdlo_out(a7_wr[698]));
			radix2 #(.width(width)) rd_st6_691  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[691]), .rdlo_in(a6_wr[699]),  .coef_in(coef[192]), .rdup_out(a7_wr[691]), .rdlo_out(a7_wr[699]));
			radix2 #(.width(width)) rd_st6_692  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[692]), .rdlo_in(a6_wr[700]),  .coef_in(coef[256]), .rdup_out(a7_wr[692]), .rdlo_out(a7_wr[700]));
			radix2 #(.width(width)) rd_st6_693  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[693]), .rdlo_in(a6_wr[701]),  .coef_in(coef[320]), .rdup_out(a7_wr[693]), .rdlo_out(a7_wr[701]));
			radix2 #(.width(width)) rd_st6_694  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[694]), .rdlo_in(a6_wr[702]),  .coef_in(coef[384]), .rdup_out(a7_wr[694]), .rdlo_out(a7_wr[702]));
			radix2 #(.width(width)) rd_st6_695  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[695]), .rdlo_in(a6_wr[703]),  .coef_in(coef[448]), .rdup_out(a7_wr[695]), .rdlo_out(a7_wr[703]));
			radix2 #(.width(width)) rd_st6_704  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[704]), .rdlo_in(a6_wr[712]),  .coef_in(coef[0]), .rdup_out(a7_wr[704]), .rdlo_out(a7_wr[712]));
			radix2 #(.width(width)) rd_st6_705  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[705]), .rdlo_in(a6_wr[713]),  .coef_in(coef[64]), .rdup_out(a7_wr[705]), .rdlo_out(a7_wr[713]));
			radix2 #(.width(width)) rd_st6_706  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[706]), .rdlo_in(a6_wr[714]),  .coef_in(coef[128]), .rdup_out(a7_wr[706]), .rdlo_out(a7_wr[714]));
			radix2 #(.width(width)) rd_st6_707  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[707]), .rdlo_in(a6_wr[715]),  .coef_in(coef[192]), .rdup_out(a7_wr[707]), .rdlo_out(a7_wr[715]));
			radix2 #(.width(width)) rd_st6_708  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[708]), .rdlo_in(a6_wr[716]),  .coef_in(coef[256]), .rdup_out(a7_wr[708]), .rdlo_out(a7_wr[716]));
			radix2 #(.width(width)) rd_st6_709  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[709]), .rdlo_in(a6_wr[717]),  .coef_in(coef[320]), .rdup_out(a7_wr[709]), .rdlo_out(a7_wr[717]));
			radix2 #(.width(width)) rd_st6_710  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[710]), .rdlo_in(a6_wr[718]),  .coef_in(coef[384]), .rdup_out(a7_wr[710]), .rdlo_out(a7_wr[718]));
			radix2 #(.width(width)) rd_st6_711  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[711]), .rdlo_in(a6_wr[719]),  .coef_in(coef[448]), .rdup_out(a7_wr[711]), .rdlo_out(a7_wr[719]));
			radix2 #(.width(width)) rd_st6_720  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[720]), .rdlo_in(a6_wr[728]),  .coef_in(coef[0]), .rdup_out(a7_wr[720]), .rdlo_out(a7_wr[728]));
			radix2 #(.width(width)) rd_st6_721  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[721]), .rdlo_in(a6_wr[729]),  .coef_in(coef[64]), .rdup_out(a7_wr[721]), .rdlo_out(a7_wr[729]));
			radix2 #(.width(width)) rd_st6_722  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[722]), .rdlo_in(a6_wr[730]),  .coef_in(coef[128]), .rdup_out(a7_wr[722]), .rdlo_out(a7_wr[730]));
			radix2 #(.width(width)) rd_st6_723  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[723]), .rdlo_in(a6_wr[731]),  .coef_in(coef[192]), .rdup_out(a7_wr[723]), .rdlo_out(a7_wr[731]));
			radix2 #(.width(width)) rd_st6_724  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[724]), .rdlo_in(a6_wr[732]),  .coef_in(coef[256]), .rdup_out(a7_wr[724]), .rdlo_out(a7_wr[732]));
			radix2 #(.width(width)) rd_st6_725  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[725]), .rdlo_in(a6_wr[733]),  .coef_in(coef[320]), .rdup_out(a7_wr[725]), .rdlo_out(a7_wr[733]));
			radix2 #(.width(width)) rd_st6_726  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[726]), .rdlo_in(a6_wr[734]),  .coef_in(coef[384]), .rdup_out(a7_wr[726]), .rdlo_out(a7_wr[734]));
			radix2 #(.width(width)) rd_st6_727  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[727]), .rdlo_in(a6_wr[735]),  .coef_in(coef[448]), .rdup_out(a7_wr[727]), .rdlo_out(a7_wr[735]));
			radix2 #(.width(width)) rd_st6_736  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[736]), .rdlo_in(a6_wr[744]),  .coef_in(coef[0]), .rdup_out(a7_wr[736]), .rdlo_out(a7_wr[744]));
			radix2 #(.width(width)) rd_st6_737  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[737]), .rdlo_in(a6_wr[745]),  .coef_in(coef[64]), .rdup_out(a7_wr[737]), .rdlo_out(a7_wr[745]));
			radix2 #(.width(width)) rd_st6_738  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[738]), .rdlo_in(a6_wr[746]),  .coef_in(coef[128]), .rdup_out(a7_wr[738]), .rdlo_out(a7_wr[746]));
			radix2 #(.width(width)) rd_st6_739  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[739]), .rdlo_in(a6_wr[747]),  .coef_in(coef[192]), .rdup_out(a7_wr[739]), .rdlo_out(a7_wr[747]));
			radix2 #(.width(width)) rd_st6_740  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[740]), .rdlo_in(a6_wr[748]),  .coef_in(coef[256]), .rdup_out(a7_wr[740]), .rdlo_out(a7_wr[748]));
			radix2 #(.width(width)) rd_st6_741  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[741]), .rdlo_in(a6_wr[749]),  .coef_in(coef[320]), .rdup_out(a7_wr[741]), .rdlo_out(a7_wr[749]));
			radix2 #(.width(width)) rd_st6_742  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[742]), .rdlo_in(a6_wr[750]),  .coef_in(coef[384]), .rdup_out(a7_wr[742]), .rdlo_out(a7_wr[750]));
			radix2 #(.width(width)) rd_st6_743  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[743]), .rdlo_in(a6_wr[751]),  .coef_in(coef[448]), .rdup_out(a7_wr[743]), .rdlo_out(a7_wr[751]));
			radix2 #(.width(width)) rd_st6_752  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[752]), .rdlo_in(a6_wr[760]),  .coef_in(coef[0]), .rdup_out(a7_wr[752]), .rdlo_out(a7_wr[760]));
			radix2 #(.width(width)) rd_st6_753  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[753]), .rdlo_in(a6_wr[761]),  .coef_in(coef[64]), .rdup_out(a7_wr[753]), .rdlo_out(a7_wr[761]));
			radix2 #(.width(width)) rd_st6_754  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[754]), .rdlo_in(a6_wr[762]),  .coef_in(coef[128]), .rdup_out(a7_wr[754]), .rdlo_out(a7_wr[762]));
			radix2 #(.width(width)) rd_st6_755  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[755]), .rdlo_in(a6_wr[763]),  .coef_in(coef[192]), .rdup_out(a7_wr[755]), .rdlo_out(a7_wr[763]));
			radix2 #(.width(width)) rd_st6_756  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[756]), .rdlo_in(a6_wr[764]),  .coef_in(coef[256]), .rdup_out(a7_wr[756]), .rdlo_out(a7_wr[764]));
			radix2 #(.width(width)) rd_st6_757  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[757]), .rdlo_in(a6_wr[765]),  .coef_in(coef[320]), .rdup_out(a7_wr[757]), .rdlo_out(a7_wr[765]));
			radix2 #(.width(width)) rd_st6_758  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[758]), .rdlo_in(a6_wr[766]),  .coef_in(coef[384]), .rdup_out(a7_wr[758]), .rdlo_out(a7_wr[766]));
			radix2 #(.width(width)) rd_st6_759  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[759]), .rdlo_in(a6_wr[767]),  .coef_in(coef[448]), .rdup_out(a7_wr[759]), .rdlo_out(a7_wr[767]));
			radix2 #(.width(width)) rd_st6_768  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[768]), .rdlo_in(a6_wr[776]),  .coef_in(coef[0]), .rdup_out(a7_wr[768]), .rdlo_out(a7_wr[776]));
			radix2 #(.width(width)) rd_st6_769  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[769]), .rdlo_in(a6_wr[777]),  .coef_in(coef[64]), .rdup_out(a7_wr[769]), .rdlo_out(a7_wr[777]));
			radix2 #(.width(width)) rd_st6_770  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[770]), .rdlo_in(a6_wr[778]),  .coef_in(coef[128]), .rdup_out(a7_wr[770]), .rdlo_out(a7_wr[778]));
			radix2 #(.width(width)) rd_st6_771  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[771]), .rdlo_in(a6_wr[779]),  .coef_in(coef[192]), .rdup_out(a7_wr[771]), .rdlo_out(a7_wr[779]));
			radix2 #(.width(width)) rd_st6_772  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[772]), .rdlo_in(a6_wr[780]),  .coef_in(coef[256]), .rdup_out(a7_wr[772]), .rdlo_out(a7_wr[780]));
			radix2 #(.width(width)) rd_st6_773  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[773]), .rdlo_in(a6_wr[781]),  .coef_in(coef[320]), .rdup_out(a7_wr[773]), .rdlo_out(a7_wr[781]));
			radix2 #(.width(width)) rd_st6_774  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[774]), .rdlo_in(a6_wr[782]),  .coef_in(coef[384]), .rdup_out(a7_wr[774]), .rdlo_out(a7_wr[782]));
			radix2 #(.width(width)) rd_st6_775  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[775]), .rdlo_in(a6_wr[783]),  .coef_in(coef[448]), .rdup_out(a7_wr[775]), .rdlo_out(a7_wr[783]));
			radix2 #(.width(width)) rd_st6_784  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[784]), .rdlo_in(a6_wr[792]),  .coef_in(coef[0]), .rdup_out(a7_wr[784]), .rdlo_out(a7_wr[792]));
			radix2 #(.width(width)) rd_st6_785  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[785]), .rdlo_in(a6_wr[793]),  .coef_in(coef[64]), .rdup_out(a7_wr[785]), .rdlo_out(a7_wr[793]));
			radix2 #(.width(width)) rd_st6_786  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[786]), .rdlo_in(a6_wr[794]),  .coef_in(coef[128]), .rdup_out(a7_wr[786]), .rdlo_out(a7_wr[794]));
			radix2 #(.width(width)) rd_st6_787  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[787]), .rdlo_in(a6_wr[795]),  .coef_in(coef[192]), .rdup_out(a7_wr[787]), .rdlo_out(a7_wr[795]));
			radix2 #(.width(width)) rd_st6_788  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[788]), .rdlo_in(a6_wr[796]),  .coef_in(coef[256]), .rdup_out(a7_wr[788]), .rdlo_out(a7_wr[796]));
			radix2 #(.width(width)) rd_st6_789  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[789]), .rdlo_in(a6_wr[797]),  .coef_in(coef[320]), .rdup_out(a7_wr[789]), .rdlo_out(a7_wr[797]));
			radix2 #(.width(width)) rd_st6_790  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[790]), .rdlo_in(a6_wr[798]),  .coef_in(coef[384]), .rdup_out(a7_wr[790]), .rdlo_out(a7_wr[798]));
			radix2 #(.width(width)) rd_st6_791  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[791]), .rdlo_in(a6_wr[799]),  .coef_in(coef[448]), .rdup_out(a7_wr[791]), .rdlo_out(a7_wr[799]));
			radix2 #(.width(width)) rd_st6_800  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[800]), .rdlo_in(a6_wr[808]),  .coef_in(coef[0]), .rdup_out(a7_wr[800]), .rdlo_out(a7_wr[808]));
			radix2 #(.width(width)) rd_st6_801  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[801]), .rdlo_in(a6_wr[809]),  .coef_in(coef[64]), .rdup_out(a7_wr[801]), .rdlo_out(a7_wr[809]));
			radix2 #(.width(width)) rd_st6_802  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[802]), .rdlo_in(a6_wr[810]),  .coef_in(coef[128]), .rdup_out(a7_wr[802]), .rdlo_out(a7_wr[810]));
			radix2 #(.width(width)) rd_st6_803  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[803]), .rdlo_in(a6_wr[811]),  .coef_in(coef[192]), .rdup_out(a7_wr[803]), .rdlo_out(a7_wr[811]));
			radix2 #(.width(width)) rd_st6_804  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[804]), .rdlo_in(a6_wr[812]),  .coef_in(coef[256]), .rdup_out(a7_wr[804]), .rdlo_out(a7_wr[812]));
			radix2 #(.width(width)) rd_st6_805  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[805]), .rdlo_in(a6_wr[813]),  .coef_in(coef[320]), .rdup_out(a7_wr[805]), .rdlo_out(a7_wr[813]));
			radix2 #(.width(width)) rd_st6_806  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[806]), .rdlo_in(a6_wr[814]),  .coef_in(coef[384]), .rdup_out(a7_wr[806]), .rdlo_out(a7_wr[814]));
			radix2 #(.width(width)) rd_st6_807  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[807]), .rdlo_in(a6_wr[815]),  .coef_in(coef[448]), .rdup_out(a7_wr[807]), .rdlo_out(a7_wr[815]));
			radix2 #(.width(width)) rd_st6_816  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[816]), .rdlo_in(a6_wr[824]),  .coef_in(coef[0]), .rdup_out(a7_wr[816]), .rdlo_out(a7_wr[824]));
			radix2 #(.width(width)) rd_st6_817  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[817]), .rdlo_in(a6_wr[825]),  .coef_in(coef[64]), .rdup_out(a7_wr[817]), .rdlo_out(a7_wr[825]));
			radix2 #(.width(width)) rd_st6_818  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[818]), .rdlo_in(a6_wr[826]),  .coef_in(coef[128]), .rdup_out(a7_wr[818]), .rdlo_out(a7_wr[826]));
			radix2 #(.width(width)) rd_st6_819  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[819]), .rdlo_in(a6_wr[827]),  .coef_in(coef[192]), .rdup_out(a7_wr[819]), .rdlo_out(a7_wr[827]));
			radix2 #(.width(width)) rd_st6_820  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[820]), .rdlo_in(a6_wr[828]),  .coef_in(coef[256]), .rdup_out(a7_wr[820]), .rdlo_out(a7_wr[828]));
			radix2 #(.width(width)) rd_st6_821  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[821]), .rdlo_in(a6_wr[829]),  .coef_in(coef[320]), .rdup_out(a7_wr[821]), .rdlo_out(a7_wr[829]));
			radix2 #(.width(width)) rd_st6_822  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[822]), .rdlo_in(a6_wr[830]),  .coef_in(coef[384]), .rdup_out(a7_wr[822]), .rdlo_out(a7_wr[830]));
			radix2 #(.width(width)) rd_st6_823  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[823]), .rdlo_in(a6_wr[831]),  .coef_in(coef[448]), .rdup_out(a7_wr[823]), .rdlo_out(a7_wr[831]));
			radix2 #(.width(width)) rd_st6_832  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[832]), .rdlo_in(a6_wr[840]),  .coef_in(coef[0]), .rdup_out(a7_wr[832]), .rdlo_out(a7_wr[840]));
			radix2 #(.width(width)) rd_st6_833  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[833]), .rdlo_in(a6_wr[841]),  .coef_in(coef[64]), .rdup_out(a7_wr[833]), .rdlo_out(a7_wr[841]));
			radix2 #(.width(width)) rd_st6_834  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[834]), .rdlo_in(a6_wr[842]),  .coef_in(coef[128]), .rdup_out(a7_wr[834]), .rdlo_out(a7_wr[842]));
			radix2 #(.width(width)) rd_st6_835  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[835]), .rdlo_in(a6_wr[843]),  .coef_in(coef[192]), .rdup_out(a7_wr[835]), .rdlo_out(a7_wr[843]));
			radix2 #(.width(width)) rd_st6_836  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[836]), .rdlo_in(a6_wr[844]),  .coef_in(coef[256]), .rdup_out(a7_wr[836]), .rdlo_out(a7_wr[844]));
			radix2 #(.width(width)) rd_st6_837  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[837]), .rdlo_in(a6_wr[845]),  .coef_in(coef[320]), .rdup_out(a7_wr[837]), .rdlo_out(a7_wr[845]));
			radix2 #(.width(width)) rd_st6_838  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[838]), .rdlo_in(a6_wr[846]),  .coef_in(coef[384]), .rdup_out(a7_wr[838]), .rdlo_out(a7_wr[846]));
			radix2 #(.width(width)) rd_st6_839  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[839]), .rdlo_in(a6_wr[847]),  .coef_in(coef[448]), .rdup_out(a7_wr[839]), .rdlo_out(a7_wr[847]));
			radix2 #(.width(width)) rd_st6_848  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[848]), .rdlo_in(a6_wr[856]),  .coef_in(coef[0]), .rdup_out(a7_wr[848]), .rdlo_out(a7_wr[856]));
			radix2 #(.width(width)) rd_st6_849  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[849]), .rdlo_in(a6_wr[857]),  .coef_in(coef[64]), .rdup_out(a7_wr[849]), .rdlo_out(a7_wr[857]));
			radix2 #(.width(width)) rd_st6_850  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[850]), .rdlo_in(a6_wr[858]),  .coef_in(coef[128]), .rdup_out(a7_wr[850]), .rdlo_out(a7_wr[858]));
			radix2 #(.width(width)) rd_st6_851  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[851]), .rdlo_in(a6_wr[859]),  .coef_in(coef[192]), .rdup_out(a7_wr[851]), .rdlo_out(a7_wr[859]));
			radix2 #(.width(width)) rd_st6_852  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[852]), .rdlo_in(a6_wr[860]),  .coef_in(coef[256]), .rdup_out(a7_wr[852]), .rdlo_out(a7_wr[860]));
			radix2 #(.width(width)) rd_st6_853  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[853]), .rdlo_in(a6_wr[861]),  .coef_in(coef[320]), .rdup_out(a7_wr[853]), .rdlo_out(a7_wr[861]));
			radix2 #(.width(width)) rd_st6_854  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[854]), .rdlo_in(a6_wr[862]),  .coef_in(coef[384]), .rdup_out(a7_wr[854]), .rdlo_out(a7_wr[862]));
			radix2 #(.width(width)) rd_st6_855  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[855]), .rdlo_in(a6_wr[863]),  .coef_in(coef[448]), .rdup_out(a7_wr[855]), .rdlo_out(a7_wr[863]));
			radix2 #(.width(width)) rd_st6_864  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[864]), .rdlo_in(a6_wr[872]),  .coef_in(coef[0]), .rdup_out(a7_wr[864]), .rdlo_out(a7_wr[872]));
			radix2 #(.width(width)) rd_st6_865  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[865]), .rdlo_in(a6_wr[873]),  .coef_in(coef[64]), .rdup_out(a7_wr[865]), .rdlo_out(a7_wr[873]));
			radix2 #(.width(width)) rd_st6_866  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[866]), .rdlo_in(a6_wr[874]),  .coef_in(coef[128]), .rdup_out(a7_wr[866]), .rdlo_out(a7_wr[874]));
			radix2 #(.width(width)) rd_st6_867  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[867]), .rdlo_in(a6_wr[875]),  .coef_in(coef[192]), .rdup_out(a7_wr[867]), .rdlo_out(a7_wr[875]));
			radix2 #(.width(width)) rd_st6_868  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[868]), .rdlo_in(a6_wr[876]),  .coef_in(coef[256]), .rdup_out(a7_wr[868]), .rdlo_out(a7_wr[876]));
			radix2 #(.width(width)) rd_st6_869  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[869]), .rdlo_in(a6_wr[877]),  .coef_in(coef[320]), .rdup_out(a7_wr[869]), .rdlo_out(a7_wr[877]));
			radix2 #(.width(width)) rd_st6_870  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[870]), .rdlo_in(a6_wr[878]),  .coef_in(coef[384]), .rdup_out(a7_wr[870]), .rdlo_out(a7_wr[878]));
			radix2 #(.width(width)) rd_st6_871  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[871]), .rdlo_in(a6_wr[879]),  .coef_in(coef[448]), .rdup_out(a7_wr[871]), .rdlo_out(a7_wr[879]));
			radix2 #(.width(width)) rd_st6_880  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[880]), .rdlo_in(a6_wr[888]),  .coef_in(coef[0]), .rdup_out(a7_wr[880]), .rdlo_out(a7_wr[888]));
			radix2 #(.width(width)) rd_st6_881  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[881]), .rdlo_in(a6_wr[889]),  .coef_in(coef[64]), .rdup_out(a7_wr[881]), .rdlo_out(a7_wr[889]));
			radix2 #(.width(width)) rd_st6_882  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[882]), .rdlo_in(a6_wr[890]),  .coef_in(coef[128]), .rdup_out(a7_wr[882]), .rdlo_out(a7_wr[890]));
			radix2 #(.width(width)) rd_st6_883  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[883]), .rdlo_in(a6_wr[891]),  .coef_in(coef[192]), .rdup_out(a7_wr[883]), .rdlo_out(a7_wr[891]));
			radix2 #(.width(width)) rd_st6_884  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[884]), .rdlo_in(a6_wr[892]),  .coef_in(coef[256]), .rdup_out(a7_wr[884]), .rdlo_out(a7_wr[892]));
			radix2 #(.width(width)) rd_st6_885  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[885]), .rdlo_in(a6_wr[893]),  .coef_in(coef[320]), .rdup_out(a7_wr[885]), .rdlo_out(a7_wr[893]));
			radix2 #(.width(width)) rd_st6_886  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[886]), .rdlo_in(a6_wr[894]),  .coef_in(coef[384]), .rdup_out(a7_wr[886]), .rdlo_out(a7_wr[894]));
			radix2 #(.width(width)) rd_st6_887  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[887]), .rdlo_in(a6_wr[895]),  .coef_in(coef[448]), .rdup_out(a7_wr[887]), .rdlo_out(a7_wr[895]));
			radix2 #(.width(width)) rd_st6_896  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[896]), .rdlo_in(a6_wr[904]),  .coef_in(coef[0]), .rdup_out(a7_wr[896]), .rdlo_out(a7_wr[904]));
			radix2 #(.width(width)) rd_st6_897  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[897]), .rdlo_in(a6_wr[905]),  .coef_in(coef[64]), .rdup_out(a7_wr[897]), .rdlo_out(a7_wr[905]));
			radix2 #(.width(width)) rd_st6_898  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[898]), .rdlo_in(a6_wr[906]),  .coef_in(coef[128]), .rdup_out(a7_wr[898]), .rdlo_out(a7_wr[906]));
			radix2 #(.width(width)) rd_st6_899  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[899]), .rdlo_in(a6_wr[907]),  .coef_in(coef[192]), .rdup_out(a7_wr[899]), .rdlo_out(a7_wr[907]));
			radix2 #(.width(width)) rd_st6_900  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[900]), .rdlo_in(a6_wr[908]),  .coef_in(coef[256]), .rdup_out(a7_wr[900]), .rdlo_out(a7_wr[908]));
			radix2 #(.width(width)) rd_st6_901  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[901]), .rdlo_in(a6_wr[909]),  .coef_in(coef[320]), .rdup_out(a7_wr[901]), .rdlo_out(a7_wr[909]));
			radix2 #(.width(width)) rd_st6_902  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[902]), .rdlo_in(a6_wr[910]),  .coef_in(coef[384]), .rdup_out(a7_wr[902]), .rdlo_out(a7_wr[910]));
			radix2 #(.width(width)) rd_st6_903  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[903]), .rdlo_in(a6_wr[911]),  .coef_in(coef[448]), .rdup_out(a7_wr[903]), .rdlo_out(a7_wr[911]));
			radix2 #(.width(width)) rd_st6_912  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[912]), .rdlo_in(a6_wr[920]),  .coef_in(coef[0]), .rdup_out(a7_wr[912]), .rdlo_out(a7_wr[920]));
			radix2 #(.width(width)) rd_st6_913  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[913]), .rdlo_in(a6_wr[921]),  .coef_in(coef[64]), .rdup_out(a7_wr[913]), .rdlo_out(a7_wr[921]));
			radix2 #(.width(width)) rd_st6_914  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[914]), .rdlo_in(a6_wr[922]),  .coef_in(coef[128]), .rdup_out(a7_wr[914]), .rdlo_out(a7_wr[922]));
			radix2 #(.width(width)) rd_st6_915  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[915]), .rdlo_in(a6_wr[923]),  .coef_in(coef[192]), .rdup_out(a7_wr[915]), .rdlo_out(a7_wr[923]));
			radix2 #(.width(width)) rd_st6_916  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[916]), .rdlo_in(a6_wr[924]),  .coef_in(coef[256]), .rdup_out(a7_wr[916]), .rdlo_out(a7_wr[924]));
			radix2 #(.width(width)) rd_st6_917  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[917]), .rdlo_in(a6_wr[925]),  .coef_in(coef[320]), .rdup_out(a7_wr[917]), .rdlo_out(a7_wr[925]));
			radix2 #(.width(width)) rd_st6_918  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[918]), .rdlo_in(a6_wr[926]),  .coef_in(coef[384]), .rdup_out(a7_wr[918]), .rdlo_out(a7_wr[926]));
			radix2 #(.width(width)) rd_st6_919  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[919]), .rdlo_in(a6_wr[927]),  .coef_in(coef[448]), .rdup_out(a7_wr[919]), .rdlo_out(a7_wr[927]));
			radix2 #(.width(width)) rd_st6_928  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[928]), .rdlo_in(a6_wr[936]),  .coef_in(coef[0]), .rdup_out(a7_wr[928]), .rdlo_out(a7_wr[936]));
			radix2 #(.width(width)) rd_st6_929  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[929]), .rdlo_in(a6_wr[937]),  .coef_in(coef[64]), .rdup_out(a7_wr[929]), .rdlo_out(a7_wr[937]));
			radix2 #(.width(width)) rd_st6_930  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[930]), .rdlo_in(a6_wr[938]),  .coef_in(coef[128]), .rdup_out(a7_wr[930]), .rdlo_out(a7_wr[938]));
			radix2 #(.width(width)) rd_st6_931  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[931]), .rdlo_in(a6_wr[939]),  .coef_in(coef[192]), .rdup_out(a7_wr[931]), .rdlo_out(a7_wr[939]));
			radix2 #(.width(width)) rd_st6_932  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[932]), .rdlo_in(a6_wr[940]),  .coef_in(coef[256]), .rdup_out(a7_wr[932]), .rdlo_out(a7_wr[940]));
			radix2 #(.width(width)) rd_st6_933  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[933]), .rdlo_in(a6_wr[941]),  .coef_in(coef[320]), .rdup_out(a7_wr[933]), .rdlo_out(a7_wr[941]));
			radix2 #(.width(width)) rd_st6_934  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[934]), .rdlo_in(a6_wr[942]),  .coef_in(coef[384]), .rdup_out(a7_wr[934]), .rdlo_out(a7_wr[942]));
			radix2 #(.width(width)) rd_st6_935  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[935]), .rdlo_in(a6_wr[943]),  .coef_in(coef[448]), .rdup_out(a7_wr[935]), .rdlo_out(a7_wr[943]));
			radix2 #(.width(width)) rd_st6_944  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[944]), .rdlo_in(a6_wr[952]),  .coef_in(coef[0]), .rdup_out(a7_wr[944]), .rdlo_out(a7_wr[952]));
			radix2 #(.width(width)) rd_st6_945  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[945]), .rdlo_in(a6_wr[953]),  .coef_in(coef[64]), .rdup_out(a7_wr[945]), .rdlo_out(a7_wr[953]));
			radix2 #(.width(width)) rd_st6_946  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[946]), .rdlo_in(a6_wr[954]),  .coef_in(coef[128]), .rdup_out(a7_wr[946]), .rdlo_out(a7_wr[954]));
			radix2 #(.width(width)) rd_st6_947  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[947]), .rdlo_in(a6_wr[955]),  .coef_in(coef[192]), .rdup_out(a7_wr[947]), .rdlo_out(a7_wr[955]));
			radix2 #(.width(width)) rd_st6_948  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[948]), .rdlo_in(a6_wr[956]),  .coef_in(coef[256]), .rdup_out(a7_wr[948]), .rdlo_out(a7_wr[956]));
			radix2 #(.width(width)) rd_st6_949  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[949]), .rdlo_in(a6_wr[957]),  .coef_in(coef[320]), .rdup_out(a7_wr[949]), .rdlo_out(a7_wr[957]));
			radix2 #(.width(width)) rd_st6_950  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[950]), .rdlo_in(a6_wr[958]),  .coef_in(coef[384]), .rdup_out(a7_wr[950]), .rdlo_out(a7_wr[958]));
			radix2 #(.width(width)) rd_st6_951  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[951]), .rdlo_in(a6_wr[959]),  .coef_in(coef[448]), .rdup_out(a7_wr[951]), .rdlo_out(a7_wr[959]));
			radix2 #(.width(width)) rd_st6_960  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[960]), .rdlo_in(a6_wr[968]),  .coef_in(coef[0]), .rdup_out(a7_wr[960]), .rdlo_out(a7_wr[968]));
			radix2 #(.width(width)) rd_st6_961  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[961]), .rdlo_in(a6_wr[969]),  .coef_in(coef[64]), .rdup_out(a7_wr[961]), .rdlo_out(a7_wr[969]));
			radix2 #(.width(width)) rd_st6_962  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[962]), .rdlo_in(a6_wr[970]),  .coef_in(coef[128]), .rdup_out(a7_wr[962]), .rdlo_out(a7_wr[970]));
			radix2 #(.width(width)) rd_st6_963  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[963]), .rdlo_in(a6_wr[971]),  .coef_in(coef[192]), .rdup_out(a7_wr[963]), .rdlo_out(a7_wr[971]));
			radix2 #(.width(width)) rd_st6_964  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[964]), .rdlo_in(a6_wr[972]),  .coef_in(coef[256]), .rdup_out(a7_wr[964]), .rdlo_out(a7_wr[972]));
			radix2 #(.width(width)) rd_st6_965  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[965]), .rdlo_in(a6_wr[973]),  .coef_in(coef[320]), .rdup_out(a7_wr[965]), .rdlo_out(a7_wr[973]));
			radix2 #(.width(width)) rd_st6_966  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[966]), .rdlo_in(a6_wr[974]),  .coef_in(coef[384]), .rdup_out(a7_wr[966]), .rdlo_out(a7_wr[974]));
			radix2 #(.width(width)) rd_st6_967  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[967]), .rdlo_in(a6_wr[975]),  .coef_in(coef[448]), .rdup_out(a7_wr[967]), .rdlo_out(a7_wr[975]));
			radix2 #(.width(width)) rd_st6_976  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[976]), .rdlo_in(a6_wr[984]),  .coef_in(coef[0]), .rdup_out(a7_wr[976]), .rdlo_out(a7_wr[984]));
			radix2 #(.width(width)) rd_st6_977  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[977]), .rdlo_in(a6_wr[985]),  .coef_in(coef[64]), .rdup_out(a7_wr[977]), .rdlo_out(a7_wr[985]));
			radix2 #(.width(width)) rd_st6_978  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[978]), .rdlo_in(a6_wr[986]),  .coef_in(coef[128]), .rdup_out(a7_wr[978]), .rdlo_out(a7_wr[986]));
			radix2 #(.width(width)) rd_st6_979  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[979]), .rdlo_in(a6_wr[987]),  .coef_in(coef[192]), .rdup_out(a7_wr[979]), .rdlo_out(a7_wr[987]));
			radix2 #(.width(width)) rd_st6_980  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[980]), .rdlo_in(a6_wr[988]),  .coef_in(coef[256]), .rdup_out(a7_wr[980]), .rdlo_out(a7_wr[988]));
			radix2 #(.width(width)) rd_st6_981  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[981]), .rdlo_in(a6_wr[989]),  .coef_in(coef[320]), .rdup_out(a7_wr[981]), .rdlo_out(a7_wr[989]));
			radix2 #(.width(width)) rd_st6_982  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[982]), .rdlo_in(a6_wr[990]),  .coef_in(coef[384]), .rdup_out(a7_wr[982]), .rdlo_out(a7_wr[990]));
			radix2 #(.width(width)) rd_st6_983  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[983]), .rdlo_in(a6_wr[991]),  .coef_in(coef[448]), .rdup_out(a7_wr[983]), .rdlo_out(a7_wr[991]));
			radix2 #(.width(width)) rd_st6_992  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[992]), .rdlo_in(a6_wr[1000]),  .coef_in(coef[0]), .rdup_out(a7_wr[992]), .rdlo_out(a7_wr[1000]));
			radix2 #(.width(width)) rd_st6_993  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[993]), .rdlo_in(a6_wr[1001]),  .coef_in(coef[64]), .rdup_out(a7_wr[993]), .rdlo_out(a7_wr[1001]));
			radix2 #(.width(width)) rd_st6_994  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[994]), .rdlo_in(a6_wr[1002]),  .coef_in(coef[128]), .rdup_out(a7_wr[994]), .rdlo_out(a7_wr[1002]));
			radix2 #(.width(width)) rd_st6_995  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[995]), .rdlo_in(a6_wr[1003]),  .coef_in(coef[192]), .rdup_out(a7_wr[995]), .rdlo_out(a7_wr[1003]));
			radix2 #(.width(width)) rd_st6_996  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[996]), .rdlo_in(a6_wr[1004]),  .coef_in(coef[256]), .rdup_out(a7_wr[996]), .rdlo_out(a7_wr[1004]));
			radix2 #(.width(width)) rd_st6_997  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[997]), .rdlo_in(a6_wr[1005]),  .coef_in(coef[320]), .rdup_out(a7_wr[997]), .rdlo_out(a7_wr[1005]));
			radix2 #(.width(width)) rd_st6_998  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[998]), .rdlo_in(a6_wr[1006]),  .coef_in(coef[384]), .rdup_out(a7_wr[998]), .rdlo_out(a7_wr[1006]));
			radix2 #(.width(width)) rd_st6_999  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[999]), .rdlo_in(a6_wr[1007]),  .coef_in(coef[448]), .rdup_out(a7_wr[999]), .rdlo_out(a7_wr[1007]));
			radix2 #(.width(width)) rd_st6_1008  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1008]), .rdlo_in(a6_wr[1016]),  .coef_in(coef[0]), .rdup_out(a7_wr[1008]), .rdlo_out(a7_wr[1016]));
			radix2 #(.width(width)) rd_st6_1009  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1009]), .rdlo_in(a6_wr[1017]),  .coef_in(coef[64]), .rdup_out(a7_wr[1009]), .rdlo_out(a7_wr[1017]));
			radix2 #(.width(width)) rd_st6_1010  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1010]), .rdlo_in(a6_wr[1018]),  .coef_in(coef[128]), .rdup_out(a7_wr[1010]), .rdlo_out(a7_wr[1018]));
			radix2 #(.width(width)) rd_st6_1011  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1011]), .rdlo_in(a6_wr[1019]),  .coef_in(coef[192]), .rdup_out(a7_wr[1011]), .rdlo_out(a7_wr[1019]));
			radix2 #(.width(width)) rd_st6_1012  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1012]), .rdlo_in(a6_wr[1020]),  .coef_in(coef[256]), .rdup_out(a7_wr[1012]), .rdlo_out(a7_wr[1020]));
			radix2 #(.width(width)) rd_st6_1013  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1013]), .rdlo_in(a6_wr[1021]),  .coef_in(coef[320]), .rdup_out(a7_wr[1013]), .rdlo_out(a7_wr[1021]));
			radix2 #(.width(width)) rd_st6_1014  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1014]), .rdlo_in(a6_wr[1022]),  .coef_in(coef[384]), .rdup_out(a7_wr[1014]), .rdlo_out(a7_wr[1022]));
			radix2 #(.width(width)) rd_st6_1015  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1015]), .rdlo_in(a6_wr[1023]),  .coef_in(coef[448]), .rdup_out(a7_wr[1015]), .rdlo_out(a7_wr[1023]));

		//--- radix stage 7
			radix2 #(.width(width)) rd_st7_0   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[0]), .rdlo_in(a7_wr[4]),  .coef_in(coef[0]), .rdup_out(a8_wr[0]), .rdlo_out(a8_wr[4]));
			radix2 #(.width(width)) rd_st7_1   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1]), .rdlo_in(a7_wr[5]),  .coef_in(coef[128]), .rdup_out(a8_wr[1]), .rdlo_out(a8_wr[5]));
			radix2 #(.width(width)) rd_st7_2   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[2]), .rdlo_in(a7_wr[6]),  .coef_in(coef[256]), .rdup_out(a8_wr[2]), .rdlo_out(a8_wr[6]));
			radix2 #(.width(width)) rd_st7_3   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[3]), .rdlo_in(a7_wr[7]),  .coef_in(coef[384]), .rdup_out(a8_wr[3]), .rdlo_out(a8_wr[7]));
			radix2 #(.width(width)) rd_st7_8   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[8]), .rdlo_in(a7_wr[12]),  .coef_in(coef[0]), .rdup_out(a8_wr[8]), .rdlo_out(a8_wr[12]));
			radix2 #(.width(width)) rd_st7_9   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[9]), .rdlo_in(a7_wr[13]),  .coef_in(coef[128]), .rdup_out(a8_wr[9]), .rdlo_out(a8_wr[13]));
			radix2 #(.width(width)) rd_st7_10  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[10]), .rdlo_in(a7_wr[14]),  .coef_in(coef[256]), .rdup_out(a8_wr[10]), .rdlo_out(a8_wr[14]));
			radix2 #(.width(width)) rd_st7_11  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[11]), .rdlo_in(a7_wr[15]),  .coef_in(coef[384]), .rdup_out(a8_wr[11]), .rdlo_out(a8_wr[15]));
			radix2 #(.width(width)) rd_st7_16  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[16]), .rdlo_in(a7_wr[20]),  .coef_in(coef[0]), .rdup_out(a8_wr[16]), .rdlo_out(a8_wr[20]));
			radix2 #(.width(width)) rd_st7_17  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[17]), .rdlo_in(a7_wr[21]),  .coef_in(coef[128]), .rdup_out(a8_wr[17]), .rdlo_out(a8_wr[21]));
			radix2 #(.width(width)) rd_st7_18  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[18]), .rdlo_in(a7_wr[22]),  .coef_in(coef[256]), .rdup_out(a8_wr[18]), .rdlo_out(a8_wr[22]));
			radix2 #(.width(width)) rd_st7_19  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[19]), .rdlo_in(a7_wr[23]),  .coef_in(coef[384]), .rdup_out(a8_wr[19]), .rdlo_out(a8_wr[23]));
			radix2 #(.width(width)) rd_st7_24  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[24]), .rdlo_in(a7_wr[28]),  .coef_in(coef[0]), .rdup_out(a8_wr[24]), .rdlo_out(a8_wr[28]));
			radix2 #(.width(width)) rd_st7_25  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[25]), .rdlo_in(a7_wr[29]),  .coef_in(coef[128]), .rdup_out(a8_wr[25]), .rdlo_out(a8_wr[29]));
			radix2 #(.width(width)) rd_st7_26  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[26]), .rdlo_in(a7_wr[30]),  .coef_in(coef[256]), .rdup_out(a8_wr[26]), .rdlo_out(a8_wr[30]));
			radix2 #(.width(width)) rd_st7_27  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[27]), .rdlo_in(a7_wr[31]),  .coef_in(coef[384]), .rdup_out(a8_wr[27]), .rdlo_out(a8_wr[31]));
			radix2 #(.width(width)) rd_st7_32  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[32]), .rdlo_in(a7_wr[36]),  .coef_in(coef[0]), .rdup_out(a8_wr[32]), .rdlo_out(a8_wr[36]));
			radix2 #(.width(width)) rd_st7_33  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[33]), .rdlo_in(a7_wr[37]),  .coef_in(coef[128]), .rdup_out(a8_wr[33]), .rdlo_out(a8_wr[37]));
			radix2 #(.width(width)) rd_st7_34  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[34]), .rdlo_in(a7_wr[38]),  .coef_in(coef[256]), .rdup_out(a8_wr[34]), .rdlo_out(a8_wr[38]));
			radix2 #(.width(width)) rd_st7_35  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[35]), .rdlo_in(a7_wr[39]),  .coef_in(coef[384]), .rdup_out(a8_wr[35]), .rdlo_out(a8_wr[39]));
			radix2 #(.width(width)) rd_st7_40  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[40]), .rdlo_in(a7_wr[44]),  .coef_in(coef[0]), .rdup_out(a8_wr[40]), .rdlo_out(a8_wr[44]));
			radix2 #(.width(width)) rd_st7_41  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[41]), .rdlo_in(a7_wr[45]),  .coef_in(coef[128]), .rdup_out(a8_wr[41]), .rdlo_out(a8_wr[45]));
			radix2 #(.width(width)) rd_st7_42  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[42]), .rdlo_in(a7_wr[46]),  .coef_in(coef[256]), .rdup_out(a8_wr[42]), .rdlo_out(a8_wr[46]));
			radix2 #(.width(width)) rd_st7_43  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[43]), .rdlo_in(a7_wr[47]),  .coef_in(coef[384]), .rdup_out(a8_wr[43]), .rdlo_out(a8_wr[47]));
			radix2 #(.width(width)) rd_st7_48  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[48]), .rdlo_in(a7_wr[52]),  .coef_in(coef[0]), .rdup_out(a8_wr[48]), .rdlo_out(a8_wr[52]));
			radix2 #(.width(width)) rd_st7_49  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[49]), .rdlo_in(a7_wr[53]),  .coef_in(coef[128]), .rdup_out(a8_wr[49]), .rdlo_out(a8_wr[53]));
			radix2 #(.width(width)) rd_st7_50  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[50]), .rdlo_in(a7_wr[54]),  .coef_in(coef[256]), .rdup_out(a8_wr[50]), .rdlo_out(a8_wr[54]));
			radix2 #(.width(width)) rd_st7_51  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[51]), .rdlo_in(a7_wr[55]),  .coef_in(coef[384]), .rdup_out(a8_wr[51]), .rdlo_out(a8_wr[55]));
			radix2 #(.width(width)) rd_st7_56  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[56]), .rdlo_in(a7_wr[60]),  .coef_in(coef[0]), .rdup_out(a8_wr[56]), .rdlo_out(a8_wr[60]));
			radix2 #(.width(width)) rd_st7_57  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[57]), .rdlo_in(a7_wr[61]),  .coef_in(coef[128]), .rdup_out(a8_wr[57]), .rdlo_out(a8_wr[61]));
			radix2 #(.width(width)) rd_st7_58  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[58]), .rdlo_in(a7_wr[62]),  .coef_in(coef[256]), .rdup_out(a8_wr[58]), .rdlo_out(a8_wr[62]));
			radix2 #(.width(width)) rd_st7_59  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[59]), .rdlo_in(a7_wr[63]),  .coef_in(coef[384]), .rdup_out(a8_wr[59]), .rdlo_out(a8_wr[63]));
			radix2 #(.width(width)) rd_st7_64  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[64]), .rdlo_in(a7_wr[68]),  .coef_in(coef[0]), .rdup_out(a8_wr[64]), .rdlo_out(a8_wr[68]));
			radix2 #(.width(width)) rd_st7_65  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[65]), .rdlo_in(a7_wr[69]),  .coef_in(coef[128]), .rdup_out(a8_wr[65]), .rdlo_out(a8_wr[69]));
			radix2 #(.width(width)) rd_st7_66  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[66]), .rdlo_in(a7_wr[70]),  .coef_in(coef[256]), .rdup_out(a8_wr[66]), .rdlo_out(a8_wr[70]));
			radix2 #(.width(width)) rd_st7_67  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[67]), .rdlo_in(a7_wr[71]),  .coef_in(coef[384]), .rdup_out(a8_wr[67]), .rdlo_out(a8_wr[71]));
			radix2 #(.width(width)) rd_st7_72  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[72]), .rdlo_in(a7_wr[76]),  .coef_in(coef[0]), .rdup_out(a8_wr[72]), .rdlo_out(a8_wr[76]));
			radix2 #(.width(width)) rd_st7_73  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[73]), .rdlo_in(a7_wr[77]),  .coef_in(coef[128]), .rdup_out(a8_wr[73]), .rdlo_out(a8_wr[77]));
			radix2 #(.width(width)) rd_st7_74  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[74]), .rdlo_in(a7_wr[78]),  .coef_in(coef[256]), .rdup_out(a8_wr[74]), .rdlo_out(a8_wr[78]));
			radix2 #(.width(width)) rd_st7_75  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[75]), .rdlo_in(a7_wr[79]),  .coef_in(coef[384]), .rdup_out(a8_wr[75]), .rdlo_out(a8_wr[79]));
			radix2 #(.width(width)) rd_st7_80  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[80]), .rdlo_in(a7_wr[84]),  .coef_in(coef[0]), .rdup_out(a8_wr[80]), .rdlo_out(a8_wr[84]));
			radix2 #(.width(width)) rd_st7_81  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[81]), .rdlo_in(a7_wr[85]),  .coef_in(coef[128]), .rdup_out(a8_wr[81]), .rdlo_out(a8_wr[85]));
			radix2 #(.width(width)) rd_st7_82  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[82]), .rdlo_in(a7_wr[86]),  .coef_in(coef[256]), .rdup_out(a8_wr[82]), .rdlo_out(a8_wr[86]));
			radix2 #(.width(width)) rd_st7_83  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[83]), .rdlo_in(a7_wr[87]),  .coef_in(coef[384]), .rdup_out(a8_wr[83]), .rdlo_out(a8_wr[87]));
			radix2 #(.width(width)) rd_st7_88  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[88]), .rdlo_in(a7_wr[92]),  .coef_in(coef[0]), .rdup_out(a8_wr[88]), .rdlo_out(a8_wr[92]));
			radix2 #(.width(width)) rd_st7_89  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[89]), .rdlo_in(a7_wr[93]),  .coef_in(coef[128]), .rdup_out(a8_wr[89]), .rdlo_out(a8_wr[93]));
			radix2 #(.width(width)) rd_st7_90  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[90]), .rdlo_in(a7_wr[94]),  .coef_in(coef[256]), .rdup_out(a8_wr[90]), .rdlo_out(a8_wr[94]));
			radix2 #(.width(width)) rd_st7_91  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[91]), .rdlo_in(a7_wr[95]),  .coef_in(coef[384]), .rdup_out(a8_wr[91]), .rdlo_out(a8_wr[95]));
			radix2 #(.width(width)) rd_st7_96  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[96]), .rdlo_in(a7_wr[100]),  .coef_in(coef[0]), .rdup_out(a8_wr[96]), .rdlo_out(a8_wr[100]));
			radix2 #(.width(width)) rd_st7_97  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[97]), .rdlo_in(a7_wr[101]),  .coef_in(coef[128]), .rdup_out(a8_wr[97]), .rdlo_out(a8_wr[101]));
			radix2 #(.width(width)) rd_st7_98  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[98]), .rdlo_in(a7_wr[102]),  .coef_in(coef[256]), .rdup_out(a8_wr[98]), .rdlo_out(a8_wr[102]));
			radix2 #(.width(width)) rd_st7_99  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[99]), .rdlo_in(a7_wr[103]),  .coef_in(coef[384]), .rdup_out(a8_wr[99]), .rdlo_out(a8_wr[103]));
			radix2 #(.width(width)) rd_st7_104  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[104]), .rdlo_in(a7_wr[108]),  .coef_in(coef[0]), .rdup_out(a8_wr[104]), .rdlo_out(a8_wr[108]));
			radix2 #(.width(width)) rd_st7_105  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[105]), .rdlo_in(a7_wr[109]),  .coef_in(coef[128]), .rdup_out(a8_wr[105]), .rdlo_out(a8_wr[109]));
			radix2 #(.width(width)) rd_st7_106  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[106]), .rdlo_in(a7_wr[110]),  .coef_in(coef[256]), .rdup_out(a8_wr[106]), .rdlo_out(a8_wr[110]));
			radix2 #(.width(width)) rd_st7_107  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[107]), .rdlo_in(a7_wr[111]),  .coef_in(coef[384]), .rdup_out(a8_wr[107]), .rdlo_out(a8_wr[111]));
			radix2 #(.width(width)) rd_st7_112  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[112]), .rdlo_in(a7_wr[116]),  .coef_in(coef[0]), .rdup_out(a8_wr[112]), .rdlo_out(a8_wr[116]));
			radix2 #(.width(width)) rd_st7_113  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[113]), .rdlo_in(a7_wr[117]),  .coef_in(coef[128]), .rdup_out(a8_wr[113]), .rdlo_out(a8_wr[117]));
			radix2 #(.width(width)) rd_st7_114  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[114]), .rdlo_in(a7_wr[118]),  .coef_in(coef[256]), .rdup_out(a8_wr[114]), .rdlo_out(a8_wr[118]));
			radix2 #(.width(width)) rd_st7_115  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[115]), .rdlo_in(a7_wr[119]),  .coef_in(coef[384]), .rdup_out(a8_wr[115]), .rdlo_out(a8_wr[119]));
			radix2 #(.width(width)) rd_st7_120  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[120]), .rdlo_in(a7_wr[124]),  .coef_in(coef[0]), .rdup_out(a8_wr[120]), .rdlo_out(a8_wr[124]));
			radix2 #(.width(width)) rd_st7_121  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[121]), .rdlo_in(a7_wr[125]),  .coef_in(coef[128]), .rdup_out(a8_wr[121]), .rdlo_out(a8_wr[125]));
			radix2 #(.width(width)) rd_st7_122  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[122]), .rdlo_in(a7_wr[126]),  .coef_in(coef[256]), .rdup_out(a8_wr[122]), .rdlo_out(a8_wr[126]));
			radix2 #(.width(width)) rd_st7_123  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[123]), .rdlo_in(a7_wr[127]),  .coef_in(coef[384]), .rdup_out(a8_wr[123]), .rdlo_out(a8_wr[127]));
			radix2 #(.width(width)) rd_st7_128  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[128]), .rdlo_in(a7_wr[132]),  .coef_in(coef[0]), .rdup_out(a8_wr[128]), .rdlo_out(a8_wr[132]));
			radix2 #(.width(width)) rd_st7_129  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[129]), .rdlo_in(a7_wr[133]),  .coef_in(coef[128]), .rdup_out(a8_wr[129]), .rdlo_out(a8_wr[133]));
			radix2 #(.width(width)) rd_st7_130  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[130]), .rdlo_in(a7_wr[134]),  .coef_in(coef[256]), .rdup_out(a8_wr[130]), .rdlo_out(a8_wr[134]));
			radix2 #(.width(width)) rd_st7_131  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[131]), .rdlo_in(a7_wr[135]),  .coef_in(coef[384]), .rdup_out(a8_wr[131]), .rdlo_out(a8_wr[135]));
			radix2 #(.width(width)) rd_st7_136  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[136]), .rdlo_in(a7_wr[140]),  .coef_in(coef[0]), .rdup_out(a8_wr[136]), .rdlo_out(a8_wr[140]));
			radix2 #(.width(width)) rd_st7_137  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[137]), .rdlo_in(a7_wr[141]),  .coef_in(coef[128]), .rdup_out(a8_wr[137]), .rdlo_out(a8_wr[141]));
			radix2 #(.width(width)) rd_st7_138  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[138]), .rdlo_in(a7_wr[142]),  .coef_in(coef[256]), .rdup_out(a8_wr[138]), .rdlo_out(a8_wr[142]));
			radix2 #(.width(width)) rd_st7_139  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[139]), .rdlo_in(a7_wr[143]),  .coef_in(coef[384]), .rdup_out(a8_wr[139]), .rdlo_out(a8_wr[143]));
			radix2 #(.width(width)) rd_st7_144  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[144]), .rdlo_in(a7_wr[148]),  .coef_in(coef[0]), .rdup_out(a8_wr[144]), .rdlo_out(a8_wr[148]));
			radix2 #(.width(width)) rd_st7_145  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[145]), .rdlo_in(a7_wr[149]),  .coef_in(coef[128]), .rdup_out(a8_wr[145]), .rdlo_out(a8_wr[149]));
			radix2 #(.width(width)) rd_st7_146  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[146]), .rdlo_in(a7_wr[150]),  .coef_in(coef[256]), .rdup_out(a8_wr[146]), .rdlo_out(a8_wr[150]));
			radix2 #(.width(width)) rd_st7_147  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[147]), .rdlo_in(a7_wr[151]),  .coef_in(coef[384]), .rdup_out(a8_wr[147]), .rdlo_out(a8_wr[151]));
			radix2 #(.width(width)) rd_st7_152  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[152]), .rdlo_in(a7_wr[156]),  .coef_in(coef[0]), .rdup_out(a8_wr[152]), .rdlo_out(a8_wr[156]));
			radix2 #(.width(width)) rd_st7_153  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[153]), .rdlo_in(a7_wr[157]),  .coef_in(coef[128]), .rdup_out(a8_wr[153]), .rdlo_out(a8_wr[157]));
			radix2 #(.width(width)) rd_st7_154  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[154]), .rdlo_in(a7_wr[158]),  .coef_in(coef[256]), .rdup_out(a8_wr[154]), .rdlo_out(a8_wr[158]));
			radix2 #(.width(width)) rd_st7_155  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[155]), .rdlo_in(a7_wr[159]),  .coef_in(coef[384]), .rdup_out(a8_wr[155]), .rdlo_out(a8_wr[159]));
			radix2 #(.width(width)) rd_st7_160  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[160]), .rdlo_in(a7_wr[164]),  .coef_in(coef[0]), .rdup_out(a8_wr[160]), .rdlo_out(a8_wr[164]));
			radix2 #(.width(width)) rd_st7_161  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[161]), .rdlo_in(a7_wr[165]),  .coef_in(coef[128]), .rdup_out(a8_wr[161]), .rdlo_out(a8_wr[165]));
			radix2 #(.width(width)) rd_st7_162  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[162]), .rdlo_in(a7_wr[166]),  .coef_in(coef[256]), .rdup_out(a8_wr[162]), .rdlo_out(a8_wr[166]));
			radix2 #(.width(width)) rd_st7_163  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[163]), .rdlo_in(a7_wr[167]),  .coef_in(coef[384]), .rdup_out(a8_wr[163]), .rdlo_out(a8_wr[167]));
			radix2 #(.width(width)) rd_st7_168  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[168]), .rdlo_in(a7_wr[172]),  .coef_in(coef[0]), .rdup_out(a8_wr[168]), .rdlo_out(a8_wr[172]));
			radix2 #(.width(width)) rd_st7_169  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[169]), .rdlo_in(a7_wr[173]),  .coef_in(coef[128]), .rdup_out(a8_wr[169]), .rdlo_out(a8_wr[173]));
			radix2 #(.width(width)) rd_st7_170  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[170]), .rdlo_in(a7_wr[174]),  .coef_in(coef[256]), .rdup_out(a8_wr[170]), .rdlo_out(a8_wr[174]));
			radix2 #(.width(width)) rd_st7_171  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[171]), .rdlo_in(a7_wr[175]),  .coef_in(coef[384]), .rdup_out(a8_wr[171]), .rdlo_out(a8_wr[175]));
			radix2 #(.width(width)) rd_st7_176  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[176]), .rdlo_in(a7_wr[180]),  .coef_in(coef[0]), .rdup_out(a8_wr[176]), .rdlo_out(a8_wr[180]));
			radix2 #(.width(width)) rd_st7_177  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[177]), .rdlo_in(a7_wr[181]),  .coef_in(coef[128]), .rdup_out(a8_wr[177]), .rdlo_out(a8_wr[181]));
			radix2 #(.width(width)) rd_st7_178  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[178]), .rdlo_in(a7_wr[182]),  .coef_in(coef[256]), .rdup_out(a8_wr[178]), .rdlo_out(a8_wr[182]));
			radix2 #(.width(width)) rd_st7_179  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[179]), .rdlo_in(a7_wr[183]),  .coef_in(coef[384]), .rdup_out(a8_wr[179]), .rdlo_out(a8_wr[183]));
			radix2 #(.width(width)) rd_st7_184  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[184]), .rdlo_in(a7_wr[188]),  .coef_in(coef[0]), .rdup_out(a8_wr[184]), .rdlo_out(a8_wr[188]));
			radix2 #(.width(width)) rd_st7_185  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[185]), .rdlo_in(a7_wr[189]),  .coef_in(coef[128]), .rdup_out(a8_wr[185]), .rdlo_out(a8_wr[189]));
			radix2 #(.width(width)) rd_st7_186  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[186]), .rdlo_in(a7_wr[190]),  .coef_in(coef[256]), .rdup_out(a8_wr[186]), .rdlo_out(a8_wr[190]));
			radix2 #(.width(width)) rd_st7_187  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[187]), .rdlo_in(a7_wr[191]),  .coef_in(coef[384]), .rdup_out(a8_wr[187]), .rdlo_out(a8_wr[191]));
			radix2 #(.width(width)) rd_st7_192  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[192]), .rdlo_in(a7_wr[196]),  .coef_in(coef[0]), .rdup_out(a8_wr[192]), .rdlo_out(a8_wr[196]));
			radix2 #(.width(width)) rd_st7_193  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[193]), .rdlo_in(a7_wr[197]),  .coef_in(coef[128]), .rdup_out(a8_wr[193]), .rdlo_out(a8_wr[197]));
			radix2 #(.width(width)) rd_st7_194  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[194]), .rdlo_in(a7_wr[198]),  .coef_in(coef[256]), .rdup_out(a8_wr[194]), .rdlo_out(a8_wr[198]));
			radix2 #(.width(width)) rd_st7_195  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[195]), .rdlo_in(a7_wr[199]),  .coef_in(coef[384]), .rdup_out(a8_wr[195]), .rdlo_out(a8_wr[199]));
			radix2 #(.width(width)) rd_st7_200  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[200]), .rdlo_in(a7_wr[204]),  .coef_in(coef[0]), .rdup_out(a8_wr[200]), .rdlo_out(a8_wr[204]));
			radix2 #(.width(width)) rd_st7_201  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[201]), .rdlo_in(a7_wr[205]),  .coef_in(coef[128]), .rdup_out(a8_wr[201]), .rdlo_out(a8_wr[205]));
			radix2 #(.width(width)) rd_st7_202  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[202]), .rdlo_in(a7_wr[206]),  .coef_in(coef[256]), .rdup_out(a8_wr[202]), .rdlo_out(a8_wr[206]));
			radix2 #(.width(width)) rd_st7_203  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[203]), .rdlo_in(a7_wr[207]),  .coef_in(coef[384]), .rdup_out(a8_wr[203]), .rdlo_out(a8_wr[207]));
			radix2 #(.width(width)) rd_st7_208  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[208]), .rdlo_in(a7_wr[212]),  .coef_in(coef[0]), .rdup_out(a8_wr[208]), .rdlo_out(a8_wr[212]));
			radix2 #(.width(width)) rd_st7_209  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[209]), .rdlo_in(a7_wr[213]),  .coef_in(coef[128]), .rdup_out(a8_wr[209]), .rdlo_out(a8_wr[213]));
			radix2 #(.width(width)) rd_st7_210  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[210]), .rdlo_in(a7_wr[214]),  .coef_in(coef[256]), .rdup_out(a8_wr[210]), .rdlo_out(a8_wr[214]));
			radix2 #(.width(width)) rd_st7_211  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[211]), .rdlo_in(a7_wr[215]),  .coef_in(coef[384]), .rdup_out(a8_wr[211]), .rdlo_out(a8_wr[215]));
			radix2 #(.width(width)) rd_st7_216  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[216]), .rdlo_in(a7_wr[220]),  .coef_in(coef[0]), .rdup_out(a8_wr[216]), .rdlo_out(a8_wr[220]));
			radix2 #(.width(width)) rd_st7_217  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[217]), .rdlo_in(a7_wr[221]),  .coef_in(coef[128]), .rdup_out(a8_wr[217]), .rdlo_out(a8_wr[221]));
			radix2 #(.width(width)) rd_st7_218  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[218]), .rdlo_in(a7_wr[222]),  .coef_in(coef[256]), .rdup_out(a8_wr[218]), .rdlo_out(a8_wr[222]));
			radix2 #(.width(width)) rd_st7_219  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[219]), .rdlo_in(a7_wr[223]),  .coef_in(coef[384]), .rdup_out(a8_wr[219]), .rdlo_out(a8_wr[223]));
			radix2 #(.width(width)) rd_st7_224  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[224]), .rdlo_in(a7_wr[228]),  .coef_in(coef[0]), .rdup_out(a8_wr[224]), .rdlo_out(a8_wr[228]));
			radix2 #(.width(width)) rd_st7_225  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[225]), .rdlo_in(a7_wr[229]),  .coef_in(coef[128]), .rdup_out(a8_wr[225]), .rdlo_out(a8_wr[229]));
			radix2 #(.width(width)) rd_st7_226  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[226]), .rdlo_in(a7_wr[230]),  .coef_in(coef[256]), .rdup_out(a8_wr[226]), .rdlo_out(a8_wr[230]));
			radix2 #(.width(width)) rd_st7_227  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[227]), .rdlo_in(a7_wr[231]),  .coef_in(coef[384]), .rdup_out(a8_wr[227]), .rdlo_out(a8_wr[231]));
			radix2 #(.width(width)) rd_st7_232  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[232]), .rdlo_in(a7_wr[236]),  .coef_in(coef[0]), .rdup_out(a8_wr[232]), .rdlo_out(a8_wr[236]));
			radix2 #(.width(width)) rd_st7_233  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[233]), .rdlo_in(a7_wr[237]),  .coef_in(coef[128]), .rdup_out(a8_wr[233]), .rdlo_out(a8_wr[237]));
			radix2 #(.width(width)) rd_st7_234  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[234]), .rdlo_in(a7_wr[238]),  .coef_in(coef[256]), .rdup_out(a8_wr[234]), .rdlo_out(a8_wr[238]));
			radix2 #(.width(width)) rd_st7_235  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[235]), .rdlo_in(a7_wr[239]),  .coef_in(coef[384]), .rdup_out(a8_wr[235]), .rdlo_out(a8_wr[239]));
			radix2 #(.width(width)) rd_st7_240  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[240]), .rdlo_in(a7_wr[244]),  .coef_in(coef[0]), .rdup_out(a8_wr[240]), .rdlo_out(a8_wr[244]));
			radix2 #(.width(width)) rd_st7_241  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[241]), .rdlo_in(a7_wr[245]),  .coef_in(coef[128]), .rdup_out(a8_wr[241]), .rdlo_out(a8_wr[245]));
			radix2 #(.width(width)) rd_st7_242  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[242]), .rdlo_in(a7_wr[246]),  .coef_in(coef[256]), .rdup_out(a8_wr[242]), .rdlo_out(a8_wr[246]));
			radix2 #(.width(width)) rd_st7_243  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[243]), .rdlo_in(a7_wr[247]),  .coef_in(coef[384]), .rdup_out(a8_wr[243]), .rdlo_out(a8_wr[247]));
			radix2 #(.width(width)) rd_st7_248  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[248]), .rdlo_in(a7_wr[252]),  .coef_in(coef[0]), .rdup_out(a8_wr[248]), .rdlo_out(a8_wr[252]));
			radix2 #(.width(width)) rd_st7_249  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[249]), .rdlo_in(a7_wr[253]),  .coef_in(coef[128]), .rdup_out(a8_wr[249]), .rdlo_out(a8_wr[253]));
			radix2 #(.width(width)) rd_st7_250  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[250]), .rdlo_in(a7_wr[254]),  .coef_in(coef[256]), .rdup_out(a8_wr[250]), .rdlo_out(a8_wr[254]));
			radix2 #(.width(width)) rd_st7_251  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[251]), .rdlo_in(a7_wr[255]),  .coef_in(coef[384]), .rdup_out(a8_wr[251]), .rdlo_out(a8_wr[255]));
			radix2 #(.width(width)) rd_st7_256  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[256]), .rdlo_in(a7_wr[260]),  .coef_in(coef[0]), .rdup_out(a8_wr[256]), .rdlo_out(a8_wr[260]));
			radix2 #(.width(width)) rd_st7_257  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[257]), .rdlo_in(a7_wr[261]),  .coef_in(coef[128]), .rdup_out(a8_wr[257]), .rdlo_out(a8_wr[261]));
			radix2 #(.width(width)) rd_st7_258  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[258]), .rdlo_in(a7_wr[262]),  .coef_in(coef[256]), .rdup_out(a8_wr[258]), .rdlo_out(a8_wr[262]));
			radix2 #(.width(width)) rd_st7_259  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[259]), .rdlo_in(a7_wr[263]),  .coef_in(coef[384]), .rdup_out(a8_wr[259]), .rdlo_out(a8_wr[263]));
			radix2 #(.width(width)) rd_st7_264  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[264]), .rdlo_in(a7_wr[268]),  .coef_in(coef[0]), .rdup_out(a8_wr[264]), .rdlo_out(a8_wr[268]));
			radix2 #(.width(width)) rd_st7_265  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[265]), .rdlo_in(a7_wr[269]),  .coef_in(coef[128]), .rdup_out(a8_wr[265]), .rdlo_out(a8_wr[269]));
			radix2 #(.width(width)) rd_st7_266  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[266]), .rdlo_in(a7_wr[270]),  .coef_in(coef[256]), .rdup_out(a8_wr[266]), .rdlo_out(a8_wr[270]));
			radix2 #(.width(width)) rd_st7_267  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[267]), .rdlo_in(a7_wr[271]),  .coef_in(coef[384]), .rdup_out(a8_wr[267]), .rdlo_out(a8_wr[271]));
			radix2 #(.width(width)) rd_st7_272  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[272]), .rdlo_in(a7_wr[276]),  .coef_in(coef[0]), .rdup_out(a8_wr[272]), .rdlo_out(a8_wr[276]));
			radix2 #(.width(width)) rd_st7_273  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[273]), .rdlo_in(a7_wr[277]),  .coef_in(coef[128]), .rdup_out(a8_wr[273]), .rdlo_out(a8_wr[277]));
			radix2 #(.width(width)) rd_st7_274  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[274]), .rdlo_in(a7_wr[278]),  .coef_in(coef[256]), .rdup_out(a8_wr[274]), .rdlo_out(a8_wr[278]));
			radix2 #(.width(width)) rd_st7_275  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[275]), .rdlo_in(a7_wr[279]),  .coef_in(coef[384]), .rdup_out(a8_wr[275]), .rdlo_out(a8_wr[279]));
			radix2 #(.width(width)) rd_st7_280  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[280]), .rdlo_in(a7_wr[284]),  .coef_in(coef[0]), .rdup_out(a8_wr[280]), .rdlo_out(a8_wr[284]));
			radix2 #(.width(width)) rd_st7_281  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[281]), .rdlo_in(a7_wr[285]),  .coef_in(coef[128]), .rdup_out(a8_wr[281]), .rdlo_out(a8_wr[285]));
			radix2 #(.width(width)) rd_st7_282  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[282]), .rdlo_in(a7_wr[286]),  .coef_in(coef[256]), .rdup_out(a8_wr[282]), .rdlo_out(a8_wr[286]));
			radix2 #(.width(width)) rd_st7_283  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[283]), .rdlo_in(a7_wr[287]),  .coef_in(coef[384]), .rdup_out(a8_wr[283]), .rdlo_out(a8_wr[287]));
			radix2 #(.width(width)) rd_st7_288  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[288]), .rdlo_in(a7_wr[292]),  .coef_in(coef[0]), .rdup_out(a8_wr[288]), .rdlo_out(a8_wr[292]));
			radix2 #(.width(width)) rd_st7_289  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[289]), .rdlo_in(a7_wr[293]),  .coef_in(coef[128]), .rdup_out(a8_wr[289]), .rdlo_out(a8_wr[293]));
			radix2 #(.width(width)) rd_st7_290  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[290]), .rdlo_in(a7_wr[294]),  .coef_in(coef[256]), .rdup_out(a8_wr[290]), .rdlo_out(a8_wr[294]));
			radix2 #(.width(width)) rd_st7_291  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[291]), .rdlo_in(a7_wr[295]),  .coef_in(coef[384]), .rdup_out(a8_wr[291]), .rdlo_out(a8_wr[295]));
			radix2 #(.width(width)) rd_st7_296  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[296]), .rdlo_in(a7_wr[300]),  .coef_in(coef[0]), .rdup_out(a8_wr[296]), .rdlo_out(a8_wr[300]));
			radix2 #(.width(width)) rd_st7_297  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[297]), .rdlo_in(a7_wr[301]),  .coef_in(coef[128]), .rdup_out(a8_wr[297]), .rdlo_out(a8_wr[301]));
			radix2 #(.width(width)) rd_st7_298  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[298]), .rdlo_in(a7_wr[302]),  .coef_in(coef[256]), .rdup_out(a8_wr[298]), .rdlo_out(a8_wr[302]));
			radix2 #(.width(width)) rd_st7_299  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[299]), .rdlo_in(a7_wr[303]),  .coef_in(coef[384]), .rdup_out(a8_wr[299]), .rdlo_out(a8_wr[303]));
			radix2 #(.width(width)) rd_st7_304  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[304]), .rdlo_in(a7_wr[308]),  .coef_in(coef[0]), .rdup_out(a8_wr[304]), .rdlo_out(a8_wr[308]));
			radix2 #(.width(width)) rd_st7_305  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[305]), .rdlo_in(a7_wr[309]),  .coef_in(coef[128]), .rdup_out(a8_wr[305]), .rdlo_out(a8_wr[309]));
			radix2 #(.width(width)) rd_st7_306  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[306]), .rdlo_in(a7_wr[310]),  .coef_in(coef[256]), .rdup_out(a8_wr[306]), .rdlo_out(a8_wr[310]));
			radix2 #(.width(width)) rd_st7_307  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[307]), .rdlo_in(a7_wr[311]),  .coef_in(coef[384]), .rdup_out(a8_wr[307]), .rdlo_out(a8_wr[311]));
			radix2 #(.width(width)) rd_st7_312  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[312]), .rdlo_in(a7_wr[316]),  .coef_in(coef[0]), .rdup_out(a8_wr[312]), .rdlo_out(a8_wr[316]));
			radix2 #(.width(width)) rd_st7_313  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[313]), .rdlo_in(a7_wr[317]),  .coef_in(coef[128]), .rdup_out(a8_wr[313]), .rdlo_out(a8_wr[317]));
			radix2 #(.width(width)) rd_st7_314  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[314]), .rdlo_in(a7_wr[318]),  .coef_in(coef[256]), .rdup_out(a8_wr[314]), .rdlo_out(a8_wr[318]));
			radix2 #(.width(width)) rd_st7_315  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[315]), .rdlo_in(a7_wr[319]),  .coef_in(coef[384]), .rdup_out(a8_wr[315]), .rdlo_out(a8_wr[319]));
			radix2 #(.width(width)) rd_st7_320  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[320]), .rdlo_in(a7_wr[324]),  .coef_in(coef[0]), .rdup_out(a8_wr[320]), .rdlo_out(a8_wr[324]));
			radix2 #(.width(width)) rd_st7_321  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[321]), .rdlo_in(a7_wr[325]),  .coef_in(coef[128]), .rdup_out(a8_wr[321]), .rdlo_out(a8_wr[325]));
			radix2 #(.width(width)) rd_st7_322  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[322]), .rdlo_in(a7_wr[326]),  .coef_in(coef[256]), .rdup_out(a8_wr[322]), .rdlo_out(a8_wr[326]));
			radix2 #(.width(width)) rd_st7_323  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[323]), .rdlo_in(a7_wr[327]),  .coef_in(coef[384]), .rdup_out(a8_wr[323]), .rdlo_out(a8_wr[327]));
			radix2 #(.width(width)) rd_st7_328  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[328]), .rdlo_in(a7_wr[332]),  .coef_in(coef[0]), .rdup_out(a8_wr[328]), .rdlo_out(a8_wr[332]));
			radix2 #(.width(width)) rd_st7_329  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[329]), .rdlo_in(a7_wr[333]),  .coef_in(coef[128]), .rdup_out(a8_wr[329]), .rdlo_out(a8_wr[333]));
			radix2 #(.width(width)) rd_st7_330  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[330]), .rdlo_in(a7_wr[334]),  .coef_in(coef[256]), .rdup_out(a8_wr[330]), .rdlo_out(a8_wr[334]));
			radix2 #(.width(width)) rd_st7_331  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[331]), .rdlo_in(a7_wr[335]),  .coef_in(coef[384]), .rdup_out(a8_wr[331]), .rdlo_out(a8_wr[335]));
			radix2 #(.width(width)) rd_st7_336  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[336]), .rdlo_in(a7_wr[340]),  .coef_in(coef[0]), .rdup_out(a8_wr[336]), .rdlo_out(a8_wr[340]));
			radix2 #(.width(width)) rd_st7_337  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[337]), .rdlo_in(a7_wr[341]),  .coef_in(coef[128]), .rdup_out(a8_wr[337]), .rdlo_out(a8_wr[341]));
			radix2 #(.width(width)) rd_st7_338  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[338]), .rdlo_in(a7_wr[342]),  .coef_in(coef[256]), .rdup_out(a8_wr[338]), .rdlo_out(a8_wr[342]));
			radix2 #(.width(width)) rd_st7_339  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[339]), .rdlo_in(a7_wr[343]),  .coef_in(coef[384]), .rdup_out(a8_wr[339]), .rdlo_out(a8_wr[343]));
			radix2 #(.width(width)) rd_st7_344  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[344]), .rdlo_in(a7_wr[348]),  .coef_in(coef[0]), .rdup_out(a8_wr[344]), .rdlo_out(a8_wr[348]));
			radix2 #(.width(width)) rd_st7_345  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[345]), .rdlo_in(a7_wr[349]),  .coef_in(coef[128]), .rdup_out(a8_wr[345]), .rdlo_out(a8_wr[349]));
			radix2 #(.width(width)) rd_st7_346  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[346]), .rdlo_in(a7_wr[350]),  .coef_in(coef[256]), .rdup_out(a8_wr[346]), .rdlo_out(a8_wr[350]));
			radix2 #(.width(width)) rd_st7_347  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[347]), .rdlo_in(a7_wr[351]),  .coef_in(coef[384]), .rdup_out(a8_wr[347]), .rdlo_out(a8_wr[351]));
			radix2 #(.width(width)) rd_st7_352  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[352]), .rdlo_in(a7_wr[356]),  .coef_in(coef[0]), .rdup_out(a8_wr[352]), .rdlo_out(a8_wr[356]));
			radix2 #(.width(width)) rd_st7_353  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[353]), .rdlo_in(a7_wr[357]),  .coef_in(coef[128]), .rdup_out(a8_wr[353]), .rdlo_out(a8_wr[357]));
			radix2 #(.width(width)) rd_st7_354  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[354]), .rdlo_in(a7_wr[358]),  .coef_in(coef[256]), .rdup_out(a8_wr[354]), .rdlo_out(a8_wr[358]));
			radix2 #(.width(width)) rd_st7_355  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[355]), .rdlo_in(a7_wr[359]),  .coef_in(coef[384]), .rdup_out(a8_wr[355]), .rdlo_out(a8_wr[359]));
			radix2 #(.width(width)) rd_st7_360  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[360]), .rdlo_in(a7_wr[364]),  .coef_in(coef[0]), .rdup_out(a8_wr[360]), .rdlo_out(a8_wr[364]));
			radix2 #(.width(width)) rd_st7_361  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[361]), .rdlo_in(a7_wr[365]),  .coef_in(coef[128]), .rdup_out(a8_wr[361]), .rdlo_out(a8_wr[365]));
			radix2 #(.width(width)) rd_st7_362  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[362]), .rdlo_in(a7_wr[366]),  .coef_in(coef[256]), .rdup_out(a8_wr[362]), .rdlo_out(a8_wr[366]));
			radix2 #(.width(width)) rd_st7_363  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[363]), .rdlo_in(a7_wr[367]),  .coef_in(coef[384]), .rdup_out(a8_wr[363]), .rdlo_out(a8_wr[367]));
			radix2 #(.width(width)) rd_st7_368  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[368]), .rdlo_in(a7_wr[372]),  .coef_in(coef[0]), .rdup_out(a8_wr[368]), .rdlo_out(a8_wr[372]));
			radix2 #(.width(width)) rd_st7_369  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[369]), .rdlo_in(a7_wr[373]),  .coef_in(coef[128]), .rdup_out(a8_wr[369]), .rdlo_out(a8_wr[373]));
			radix2 #(.width(width)) rd_st7_370  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[370]), .rdlo_in(a7_wr[374]),  .coef_in(coef[256]), .rdup_out(a8_wr[370]), .rdlo_out(a8_wr[374]));
			radix2 #(.width(width)) rd_st7_371  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[371]), .rdlo_in(a7_wr[375]),  .coef_in(coef[384]), .rdup_out(a8_wr[371]), .rdlo_out(a8_wr[375]));
			radix2 #(.width(width)) rd_st7_376  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[376]), .rdlo_in(a7_wr[380]),  .coef_in(coef[0]), .rdup_out(a8_wr[376]), .rdlo_out(a8_wr[380]));
			radix2 #(.width(width)) rd_st7_377  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[377]), .rdlo_in(a7_wr[381]),  .coef_in(coef[128]), .rdup_out(a8_wr[377]), .rdlo_out(a8_wr[381]));
			radix2 #(.width(width)) rd_st7_378  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[378]), .rdlo_in(a7_wr[382]),  .coef_in(coef[256]), .rdup_out(a8_wr[378]), .rdlo_out(a8_wr[382]));
			radix2 #(.width(width)) rd_st7_379  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[379]), .rdlo_in(a7_wr[383]),  .coef_in(coef[384]), .rdup_out(a8_wr[379]), .rdlo_out(a8_wr[383]));
			radix2 #(.width(width)) rd_st7_384  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[384]), .rdlo_in(a7_wr[388]),  .coef_in(coef[0]), .rdup_out(a8_wr[384]), .rdlo_out(a8_wr[388]));
			radix2 #(.width(width)) rd_st7_385  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[385]), .rdlo_in(a7_wr[389]),  .coef_in(coef[128]), .rdup_out(a8_wr[385]), .rdlo_out(a8_wr[389]));
			radix2 #(.width(width)) rd_st7_386  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[386]), .rdlo_in(a7_wr[390]),  .coef_in(coef[256]), .rdup_out(a8_wr[386]), .rdlo_out(a8_wr[390]));
			radix2 #(.width(width)) rd_st7_387  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[387]), .rdlo_in(a7_wr[391]),  .coef_in(coef[384]), .rdup_out(a8_wr[387]), .rdlo_out(a8_wr[391]));
			radix2 #(.width(width)) rd_st7_392  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[392]), .rdlo_in(a7_wr[396]),  .coef_in(coef[0]), .rdup_out(a8_wr[392]), .rdlo_out(a8_wr[396]));
			radix2 #(.width(width)) rd_st7_393  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[393]), .rdlo_in(a7_wr[397]),  .coef_in(coef[128]), .rdup_out(a8_wr[393]), .rdlo_out(a8_wr[397]));
			radix2 #(.width(width)) rd_st7_394  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[394]), .rdlo_in(a7_wr[398]),  .coef_in(coef[256]), .rdup_out(a8_wr[394]), .rdlo_out(a8_wr[398]));
			radix2 #(.width(width)) rd_st7_395  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[395]), .rdlo_in(a7_wr[399]),  .coef_in(coef[384]), .rdup_out(a8_wr[395]), .rdlo_out(a8_wr[399]));
			radix2 #(.width(width)) rd_st7_400  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[400]), .rdlo_in(a7_wr[404]),  .coef_in(coef[0]), .rdup_out(a8_wr[400]), .rdlo_out(a8_wr[404]));
			radix2 #(.width(width)) rd_st7_401  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[401]), .rdlo_in(a7_wr[405]),  .coef_in(coef[128]), .rdup_out(a8_wr[401]), .rdlo_out(a8_wr[405]));
			radix2 #(.width(width)) rd_st7_402  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[402]), .rdlo_in(a7_wr[406]),  .coef_in(coef[256]), .rdup_out(a8_wr[402]), .rdlo_out(a8_wr[406]));
			radix2 #(.width(width)) rd_st7_403  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[403]), .rdlo_in(a7_wr[407]),  .coef_in(coef[384]), .rdup_out(a8_wr[403]), .rdlo_out(a8_wr[407]));
			radix2 #(.width(width)) rd_st7_408  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[408]), .rdlo_in(a7_wr[412]),  .coef_in(coef[0]), .rdup_out(a8_wr[408]), .rdlo_out(a8_wr[412]));
			radix2 #(.width(width)) rd_st7_409  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[409]), .rdlo_in(a7_wr[413]),  .coef_in(coef[128]), .rdup_out(a8_wr[409]), .rdlo_out(a8_wr[413]));
			radix2 #(.width(width)) rd_st7_410  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[410]), .rdlo_in(a7_wr[414]),  .coef_in(coef[256]), .rdup_out(a8_wr[410]), .rdlo_out(a8_wr[414]));
			radix2 #(.width(width)) rd_st7_411  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[411]), .rdlo_in(a7_wr[415]),  .coef_in(coef[384]), .rdup_out(a8_wr[411]), .rdlo_out(a8_wr[415]));
			radix2 #(.width(width)) rd_st7_416  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[416]), .rdlo_in(a7_wr[420]),  .coef_in(coef[0]), .rdup_out(a8_wr[416]), .rdlo_out(a8_wr[420]));
			radix2 #(.width(width)) rd_st7_417  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[417]), .rdlo_in(a7_wr[421]),  .coef_in(coef[128]), .rdup_out(a8_wr[417]), .rdlo_out(a8_wr[421]));
			radix2 #(.width(width)) rd_st7_418  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[418]), .rdlo_in(a7_wr[422]),  .coef_in(coef[256]), .rdup_out(a8_wr[418]), .rdlo_out(a8_wr[422]));
			radix2 #(.width(width)) rd_st7_419  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[419]), .rdlo_in(a7_wr[423]),  .coef_in(coef[384]), .rdup_out(a8_wr[419]), .rdlo_out(a8_wr[423]));
			radix2 #(.width(width)) rd_st7_424  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[424]), .rdlo_in(a7_wr[428]),  .coef_in(coef[0]), .rdup_out(a8_wr[424]), .rdlo_out(a8_wr[428]));
			radix2 #(.width(width)) rd_st7_425  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[425]), .rdlo_in(a7_wr[429]),  .coef_in(coef[128]), .rdup_out(a8_wr[425]), .rdlo_out(a8_wr[429]));
			radix2 #(.width(width)) rd_st7_426  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[426]), .rdlo_in(a7_wr[430]),  .coef_in(coef[256]), .rdup_out(a8_wr[426]), .rdlo_out(a8_wr[430]));
			radix2 #(.width(width)) rd_st7_427  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[427]), .rdlo_in(a7_wr[431]),  .coef_in(coef[384]), .rdup_out(a8_wr[427]), .rdlo_out(a8_wr[431]));
			radix2 #(.width(width)) rd_st7_432  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[432]), .rdlo_in(a7_wr[436]),  .coef_in(coef[0]), .rdup_out(a8_wr[432]), .rdlo_out(a8_wr[436]));
			radix2 #(.width(width)) rd_st7_433  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[433]), .rdlo_in(a7_wr[437]),  .coef_in(coef[128]), .rdup_out(a8_wr[433]), .rdlo_out(a8_wr[437]));
			radix2 #(.width(width)) rd_st7_434  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[434]), .rdlo_in(a7_wr[438]),  .coef_in(coef[256]), .rdup_out(a8_wr[434]), .rdlo_out(a8_wr[438]));
			radix2 #(.width(width)) rd_st7_435  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[435]), .rdlo_in(a7_wr[439]),  .coef_in(coef[384]), .rdup_out(a8_wr[435]), .rdlo_out(a8_wr[439]));
			radix2 #(.width(width)) rd_st7_440  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[440]), .rdlo_in(a7_wr[444]),  .coef_in(coef[0]), .rdup_out(a8_wr[440]), .rdlo_out(a8_wr[444]));
			radix2 #(.width(width)) rd_st7_441  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[441]), .rdlo_in(a7_wr[445]),  .coef_in(coef[128]), .rdup_out(a8_wr[441]), .rdlo_out(a8_wr[445]));
			radix2 #(.width(width)) rd_st7_442  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[442]), .rdlo_in(a7_wr[446]),  .coef_in(coef[256]), .rdup_out(a8_wr[442]), .rdlo_out(a8_wr[446]));
			radix2 #(.width(width)) rd_st7_443  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[443]), .rdlo_in(a7_wr[447]),  .coef_in(coef[384]), .rdup_out(a8_wr[443]), .rdlo_out(a8_wr[447]));
			radix2 #(.width(width)) rd_st7_448  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[448]), .rdlo_in(a7_wr[452]),  .coef_in(coef[0]), .rdup_out(a8_wr[448]), .rdlo_out(a8_wr[452]));
			radix2 #(.width(width)) rd_st7_449  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[449]), .rdlo_in(a7_wr[453]),  .coef_in(coef[128]), .rdup_out(a8_wr[449]), .rdlo_out(a8_wr[453]));
			radix2 #(.width(width)) rd_st7_450  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[450]), .rdlo_in(a7_wr[454]),  .coef_in(coef[256]), .rdup_out(a8_wr[450]), .rdlo_out(a8_wr[454]));
			radix2 #(.width(width)) rd_st7_451  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[451]), .rdlo_in(a7_wr[455]),  .coef_in(coef[384]), .rdup_out(a8_wr[451]), .rdlo_out(a8_wr[455]));
			radix2 #(.width(width)) rd_st7_456  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[456]), .rdlo_in(a7_wr[460]),  .coef_in(coef[0]), .rdup_out(a8_wr[456]), .rdlo_out(a8_wr[460]));
			radix2 #(.width(width)) rd_st7_457  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[457]), .rdlo_in(a7_wr[461]),  .coef_in(coef[128]), .rdup_out(a8_wr[457]), .rdlo_out(a8_wr[461]));
			radix2 #(.width(width)) rd_st7_458  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[458]), .rdlo_in(a7_wr[462]),  .coef_in(coef[256]), .rdup_out(a8_wr[458]), .rdlo_out(a8_wr[462]));
			radix2 #(.width(width)) rd_st7_459  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[459]), .rdlo_in(a7_wr[463]),  .coef_in(coef[384]), .rdup_out(a8_wr[459]), .rdlo_out(a8_wr[463]));
			radix2 #(.width(width)) rd_st7_464  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[464]), .rdlo_in(a7_wr[468]),  .coef_in(coef[0]), .rdup_out(a8_wr[464]), .rdlo_out(a8_wr[468]));
			radix2 #(.width(width)) rd_st7_465  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[465]), .rdlo_in(a7_wr[469]),  .coef_in(coef[128]), .rdup_out(a8_wr[465]), .rdlo_out(a8_wr[469]));
			radix2 #(.width(width)) rd_st7_466  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[466]), .rdlo_in(a7_wr[470]),  .coef_in(coef[256]), .rdup_out(a8_wr[466]), .rdlo_out(a8_wr[470]));
			radix2 #(.width(width)) rd_st7_467  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[467]), .rdlo_in(a7_wr[471]),  .coef_in(coef[384]), .rdup_out(a8_wr[467]), .rdlo_out(a8_wr[471]));
			radix2 #(.width(width)) rd_st7_472  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[472]), .rdlo_in(a7_wr[476]),  .coef_in(coef[0]), .rdup_out(a8_wr[472]), .rdlo_out(a8_wr[476]));
			radix2 #(.width(width)) rd_st7_473  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[473]), .rdlo_in(a7_wr[477]),  .coef_in(coef[128]), .rdup_out(a8_wr[473]), .rdlo_out(a8_wr[477]));
			radix2 #(.width(width)) rd_st7_474  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[474]), .rdlo_in(a7_wr[478]),  .coef_in(coef[256]), .rdup_out(a8_wr[474]), .rdlo_out(a8_wr[478]));
			radix2 #(.width(width)) rd_st7_475  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[475]), .rdlo_in(a7_wr[479]),  .coef_in(coef[384]), .rdup_out(a8_wr[475]), .rdlo_out(a8_wr[479]));
			radix2 #(.width(width)) rd_st7_480  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[480]), .rdlo_in(a7_wr[484]),  .coef_in(coef[0]), .rdup_out(a8_wr[480]), .rdlo_out(a8_wr[484]));
			radix2 #(.width(width)) rd_st7_481  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[481]), .rdlo_in(a7_wr[485]),  .coef_in(coef[128]), .rdup_out(a8_wr[481]), .rdlo_out(a8_wr[485]));
			radix2 #(.width(width)) rd_st7_482  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[482]), .rdlo_in(a7_wr[486]),  .coef_in(coef[256]), .rdup_out(a8_wr[482]), .rdlo_out(a8_wr[486]));
			radix2 #(.width(width)) rd_st7_483  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[483]), .rdlo_in(a7_wr[487]),  .coef_in(coef[384]), .rdup_out(a8_wr[483]), .rdlo_out(a8_wr[487]));
			radix2 #(.width(width)) rd_st7_488  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[488]), .rdlo_in(a7_wr[492]),  .coef_in(coef[0]), .rdup_out(a8_wr[488]), .rdlo_out(a8_wr[492]));
			radix2 #(.width(width)) rd_st7_489  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[489]), .rdlo_in(a7_wr[493]),  .coef_in(coef[128]), .rdup_out(a8_wr[489]), .rdlo_out(a8_wr[493]));
			radix2 #(.width(width)) rd_st7_490  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[490]), .rdlo_in(a7_wr[494]),  .coef_in(coef[256]), .rdup_out(a8_wr[490]), .rdlo_out(a8_wr[494]));
			radix2 #(.width(width)) rd_st7_491  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[491]), .rdlo_in(a7_wr[495]),  .coef_in(coef[384]), .rdup_out(a8_wr[491]), .rdlo_out(a8_wr[495]));
			radix2 #(.width(width)) rd_st7_496  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[496]), .rdlo_in(a7_wr[500]),  .coef_in(coef[0]), .rdup_out(a8_wr[496]), .rdlo_out(a8_wr[500]));
			radix2 #(.width(width)) rd_st7_497  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[497]), .rdlo_in(a7_wr[501]),  .coef_in(coef[128]), .rdup_out(a8_wr[497]), .rdlo_out(a8_wr[501]));
			radix2 #(.width(width)) rd_st7_498  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[498]), .rdlo_in(a7_wr[502]),  .coef_in(coef[256]), .rdup_out(a8_wr[498]), .rdlo_out(a8_wr[502]));
			radix2 #(.width(width)) rd_st7_499  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[499]), .rdlo_in(a7_wr[503]),  .coef_in(coef[384]), .rdup_out(a8_wr[499]), .rdlo_out(a8_wr[503]));
			radix2 #(.width(width)) rd_st7_504  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[504]), .rdlo_in(a7_wr[508]),  .coef_in(coef[0]), .rdup_out(a8_wr[504]), .rdlo_out(a8_wr[508]));
			radix2 #(.width(width)) rd_st7_505  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[505]), .rdlo_in(a7_wr[509]),  .coef_in(coef[128]), .rdup_out(a8_wr[505]), .rdlo_out(a8_wr[509]));
			radix2 #(.width(width)) rd_st7_506  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[506]), .rdlo_in(a7_wr[510]),  .coef_in(coef[256]), .rdup_out(a8_wr[506]), .rdlo_out(a8_wr[510]));
			radix2 #(.width(width)) rd_st7_507  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[507]), .rdlo_in(a7_wr[511]),  .coef_in(coef[384]), .rdup_out(a8_wr[507]), .rdlo_out(a8_wr[511]));
			radix2 #(.width(width)) rd_st7_512  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[512]), .rdlo_in(a7_wr[516]),  .coef_in(coef[0]), .rdup_out(a8_wr[512]), .rdlo_out(a8_wr[516]));
			radix2 #(.width(width)) rd_st7_513  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[513]), .rdlo_in(a7_wr[517]),  .coef_in(coef[128]), .rdup_out(a8_wr[513]), .rdlo_out(a8_wr[517]));
			radix2 #(.width(width)) rd_st7_514  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[514]), .rdlo_in(a7_wr[518]),  .coef_in(coef[256]), .rdup_out(a8_wr[514]), .rdlo_out(a8_wr[518]));
			radix2 #(.width(width)) rd_st7_515  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[515]), .rdlo_in(a7_wr[519]),  .coef_in(coef[384]), .rdup_out(a8_wr[515]), .rdlo_out(a8_wr[519]));
			radix2 #(.width(width)) rd_st7_520  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[520]), .rdlo_in(a7_wr[524]),  .coef_in(coef[0]), .rdup_out(a8_wr[520]), .rdlo_out(a8_wr[524]));
			radix2 #(.width(width)) rd_st7_521  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[521]), .rdlo_in(a7_wr[525]),  .coef_in(coef[128]), .rdup_out(a8_wr[521]), .rdlo_out(a8_wr[525]));
			radix2 #(.width(width)) rd_st7_522  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[522]), .rdlo_in(a7_wr[526]),  .coef_in(coef[256]), .rdup_out(a8_wr[522]), .rdlo_out(a8_wr[526]));
			radix2 #(.width(width)) rd_st7_523  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[523]), .rdlo_in(a7_wr[527]),  .coef_in(coef[384]), .rdup_out(a8_wr[523]), .rdlo_out(a8_wr[527]));
			radix2 #(.width(width)) rd_st7_528  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[528]), .rdlo_in(a7_wr[532]),  .coef_in(coef[0]), .rdup_out(a8_wr[528]), .rdlo_out(a8_wr[532]));
			radix2 #(.width(width)) rd_st7_529  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[529]), .rdlo_in(a7_wr[533]),  .coef_in(coef[128]), .rdup_out(a8_wr[529]), .rdlo_out(a8_wr[533]));
			radix2 #(.width(width)) rd_st7_530  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[530]), .rdlo_in(a7_wr[534]),  .coef_in(coef[256]), .rdup_out(a8_wr[530]), .rdlo_out(a8_wr[534]));
			radix2 #(.width(width)) rd_st7_531  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[531]), .rdlo_in(a7_wr[535]),  .coef_in(coef[384]), .rdup_out(a8_wr[531]), .rdlo_out(a8_wr[535]));
			radix2 #(.width(width)) rd_st7_536  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[536]), .rdlo_in(a7_wr[540]),  .coef_in(coef[0]), .rdup_out(a8_wr[536]), .rdlo_out(a8_wr[540]));
			radix2 #(.width(width)) rd_st7_537  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[537]), .rdlo_in(a7_wr[541]),  .coef_in(coef[128]), .rdup_out(a8_wr[537]), .rdlo_out(a8_wr[541]));
			radix2 #(.width(width)) rd_st7_538  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[538]), .rdlo_in(a7_wr[542]),  .coef_in(coef[256]), .rdup_out(a8_wr[538]), .rdlo_out(a8_wr[542]));
			radix2 #(.width(width)) rd_st7_539  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[539]), .rdlo_in(a7_wr[543]),  .coef_in(coef[384]), .rdup_out(a8_wr[539]), .rdlo_out(a8_wr[543]));
			radix2 #(.width(width)) rd_st7_544  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[544]), .rdlo_in(a7_wr[548]),  .coef_in(coef[0]), .rdup_out(a8_wr[544]), .rdlo_out(a8_wr[548]));
			radix2 #(.width(width)) rd_st7_545  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[545]), .rdlo_in(a7_wr[549]),  .coef_in(coef[128]), .rdup_out(a8_wr[545]), .rdlo_out(a8_wr[549]));
			radix2 #(.width(width)) rd_st7_546  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[546]), .rdlo_in(a7_wr[550]),  .coef_in(coef[256]), .rdup_out(a8_wr[546]), .rdlo_out(a8_wr[550]));
			radix2 #(.width(width)) rd_st7_547  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[547]), .rdlo_in(a7_wr[551]),  .coef_in(coef[384]), .rdup_out(a8_wr[547]), .rdlo_out(a8_wr[551]));
			radix2 #(.width(width)) rd_st7_552  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[552]), .rdlo_in(a7_wr[556]),  .coef_in(coef[0]), .rdup_out(a8_wr[552]), .rdlo_out(a8_wr[556]));
			radix2 #(.width(width)) rd_st7_553  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[553]), .rdlo_in(a7_wr[557]),  .coef_in(coef[128]), .rdup_out(a8_wr[553]), .rdlo_out(a8_wr[557]));
			radix2 #(.width(width)) rd_st7_554  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[554]), .rdlo_in(a7_wr[558]),  .coef_in(coef[256]), .rdup_out(a8_wr[554]), .rdlo_out(a8_wr[558]));
			radix2 #(.width(width)) rd_st7_555  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[555]), .rdlo_in(a7_wr[559]),  .coef_in(coef[384]), .rdup_out(a8_wr[555]), .rdlo_out(a8_wr[559]));
			radix2 #(.width(width)) rd_st7_560  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[560]), .rdlo_in(a7_wr[564]),  .coef_in(coef[0]), .rdup_out(a8_wr[560]), .rdlo_out(a8_wr[564]));
			radix2 #(.width(width)) rd_st7_561  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[561]), .rdlo_in(a7_wr[565]),  .coef_in(coef[128]), .rdup_out(a8_wr[561]), .rdlo_out(a8_wr[565]));
			radix2 #(.width(width)) rd_st7_562  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[562]), .rdlo_in(a7_wr[566]),  .coef_in(coef[256]), .rdup_out(a8_wr[562]), .rdlo_out(a8_wr[566]));
			radix2 #(.width(width)) rd_st7_563  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[563]), .rdlo_in(a7_wr[567]),  .coef_in(coef[384]), .rdup_out(a8_wr[563]), .rdlo_out(a8_wr[567]));
			radix2 #(.width(width)) rd_st7_568  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[568]), .rdlo_in(a7_wr[572]),  .coef_in(coef[0]), .rdup_out(a8_wr[568]), .rdlo_out(a8_wr[572]));
			radix2 #(.width(width)) rd_st7_569  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[569]), .rdlo_in(a7_wr[573]),  .coef_in(coef[128]), .rdup_out(a8_wr[569]), .rdlo_out(a8_wr[573]));
			radix2 #(.width(width)) rd_st7_570  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[570]), .rdlo_in(a7_wr[574]),  .coef_in(coef[256]), .rdup_out(a8_wr[570]), .rdlo_out(a8_wr[574]));
			radix2 #(.width(width)) rd_st7_571  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[571]), .rdlo_in(a7_wr[575]),  .coef_in(coef[384]), .rdup_out(a8_wr[571]), .rdlo_out(a8_wr[575]));
			radix2 #(.width(width)) rd_st7_576  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[576]), .rdlo_in(a7_wr[580]),  .coef_in(coef[0]), .rdup_out(a8_wr[576]), .rdlo_out(a8_wr[580]));
			radix2 #(.width(width)) rd_st7_577  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[577]), .rdlo_in(a7_wr[581]),  .coef_in(coef[128]), .rdup_out(a8_wr[577]), .rdlo_out(a8_wr[581]));
			radix2 #(.width(width)) rd_st7_578  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[578]), .rdlo_in(a7_wr[582]),  .coef_in(coef[256]), .rdup_out(a8_wr[578]), .rdlo_out(a8_wr[582]));
			radix2 #(.width(width)) rd_st7_579  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[579]), .rdlo_in(a7_wr[583]),  .coef_in(coef[384]), .rdup_out(a8_wr[579]), .rdlo_out(a8_wr[583]));
			radix2 #(.width(width)) rd_st7_584  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[584]), .rdlo_in(a7_wr[588]),  .coef_in(coef[0]), .rdup_out(a8_wr[584]), .rdlo_out(a8_wr[588]));
			radix2 #(.width(width)) rd_st7_585  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[585]), .rdlo_in(a7_wr[589]),  .coef_in(coef[128]), .rdup_out(a8_wr[585]), .rdlo_out(a8_wr[589]));
			radix2 #(.width(width)) rd_st7_586  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[586]), .rdlo_in(a7_wr[590]),  .coef_in(coef[256]), .rdup_out(a8_wr[586]), .rdlo_out(a8_wr[590]));
			radix2 #(.width(width)) rd_st7_587  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[587]), .rdlo_in(a7_wr[591]),  .coef_in(coef[384]), .rdup_out(a8_wr[587]), .rdlo_out(a8_wr[591]));
			radix2 #(.width(width)) rd_st7_592  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[592]), .rdlo_in(a7_wr[596]),  .coef_in(coef[0]), .rdup_out(a8_wr[592]), .rdlo_out(a8_wr[596]));
			radix2 #(.width(width)) rd_st7_593  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[593]), .rdlo_in(a7_wr[597]),  .coef_in(coef[128]), .rdup_out(a8_wr[593]), .rdlo_out(a8_wr[597]));
			radix2 #(.width(width)) rd_st7_594  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[594]), .rdlo_in(a7_wr[598]),  .coef_in(coef[256]), .rdup_out(a8_wr[594]), .rdlo_out(a8_wr[598]));
			radix2 #(.width(width)) rd_st7_595  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[595]), .rdlo_in(a7_wr[599]),  .coef_in(coef[384]), .rdup_out(a8_wr[595]), .rdlo_out(a8_wr[599]));
			radix2 #(.width(width)) rd_st7_600  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[600]), .rdlo_in(a7_wr[604]),  .coef_in(coef[0]), .rdup_out(a8_wr[600]), .rdlo_out(a8_wr[604]));
			radix2 #(.width(width)) rd_st7_601  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[601]), .rdlo_in(a7_wr[605]),  .coef_in(coef[128]), .rdup_out(a8_wr[601]), .rdlo_out(a8_wr[605]));
			radix2 #(.width(width)) rd_st7_602  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[602]), .rdlo_in(a7_wr[606]),  .coef_in(coef[256]), .rdup_out(a8_wr[602]), .rdlo_out(a8_wr[606]));
			radix2 #(.width(width)) rd_st7_603  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[603]), .rdlo_in(a7_wr[607]),  .coef_in(coef[384]), .rdup_out(a8_wr[603]), .rdlo_out(a8_wr[607]));
			radix2 #(.width(width)) rd_st7_608  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[608]), .rdlo_in(a7_wr[612]),  .coef_in(coef[0]), .rdup_out(a8_wr[608]), .rdlo_out(a8_wr[612]));
			radix2 #(.width(width)) rd_st7_609  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[609]), .rdlo_in(a7_wr[613]),  .coef_in(coef[128]), .rdup_out(a8_wr[609]), .rdlo_out(a8_wr[613]));
			radix2 #(.width(width)) rd_st7_610  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[610]), .rdlo_in(a7_wr[614]),  .coef_in(coef[256]), .rdup_out(a8_wr[610]), .rdlo_out(a8_wr[614]));
			radix2 #(.width(width)) rd_st7_611  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[611]), .rdlo_in(a7_wr[615]),  .coef_in(coef[384]), .rdup_out(a8_wr[611]), .rdlo_out(a8_wr[615]));
			radix2 #(.width(width)) rd_st7_616  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[616]), .rdlo_in(a7_wr[620]),  .coef_in(coef[0]), .rdup_out(a8_wr[616]), .rdlo_out(a8_wr[620]));
			radix2 #(.width(width)) rd_st7_617  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[617]), .rdlo_in(a7_wr[621]),  .coef_in(coef[128]), .rdup_out(a8_wr[617]), .rdlo_out(a8_wr[621]));
			radix2 #(.width(width)) rd_st7_618  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[618]), .rdlo_in(a7_wr[622]),  .coef_in(coef[256]), .rdup_out(a8_wr[618]), .rdlo_out(a8_wr[622]));
			radix2 #(.width(width)) rd_st7_619  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[619]), .rdlo_in(a7_wr[623]),  .coef_in(coef[384]), .rdup_out(a8_wr[619]), .rdlo_out(a8_wr[623]));
			radix2 #(.width(width)) rd_st7_624  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[624]), .rdlo_in(a7_wr[628]),  .coef_in(coef[0]), .rdup_out(a8_wr[624]), .rdlo_out(a8_wr[628]));
			radix2 #(.width(width)) rd_st7_625  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[625]), .rdlo_in(a7_wr[629]),  .coef_in(coef[128]), .rdup_out(a8_wr[625]), .rdlo_out(a8_wr[629]));
			radix2 #(.width(width)) rd_st7_626  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[626]), .rdlo_in(a7_wr[630]),  .coef_in(coef[256]), .rdup_out(a8_wr[626]), .rdlo_out(a8_wr[630]));
			radix2 #(.width(width)) rd_st7_627  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[627]), .rdlo_in(a7_wr[631]),  .coef_in(coef[384]), .rdup_out(a8_wr[627]), .rdlo_out(a8_wr[631]));
			radix2 #(.width(width)) rd_st7_632  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[632]), .rdlo_in(a7_wr[636]),  .coef_in(coef[0]), .rdup_out(a8_wr[632]), .rdlo_out(a8_wr[636]));
			radix2 #(.width(width)) rd_st7_633  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[633]), .rdlo_in(a7_wr[637]),  .coef_in(coef[128]), .rdup_out(a8_wr[633]), .rdlo_out(a8_wr[637]));
			radix2 #(.width(width)) rd_st7_634  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[634]), .rdlo_in(a7_wr[638]),  .coef_in(coef[256]), .rdup_out(a8_wr[634]), .rdlo_out(a8_wr[638]));
			radix2 #(.width(width)) rd_st7_635  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[635]), .rdlo_in(a7_wr[639]),  .coef_in(coef[384]), .rdup_out(a8_wr[635]), .rdlo_out(a8_wr[639]));
			radix2 #(.width(width)) rd_st7_640  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[640]), .rdlo_in(a7_wr[644]),  .coef_in(coef[0]), .rdup_out(a8_wr[640]), .rdlo_out(a8_wr[644]));
			radix2 #(.width(width)) rd_st7_641  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[641]), .rdlo_in(a7_wr[645]),  .coef_in(coef[128]), .rdup_out(a8_wr[641]), .rdlo_out(a8_wr[645]));
			radix2 #(.width(width)) rd_st7_642  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[642]), .rdlo_in(a7_wr[646]),  .coef_in(coef[256]), .rdup_out(a8_wr[642]), .rdlo_out(a8_wr[646]));
			radix2 #(.width(width)) rd_st7_643  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[643]), .rdlo_in(a7_wr[647]),  .coef_in(coef[384]), .rdup_out(a8_wr[643]), .rdlo_out(a8_wr[647]));
			radix2 #(.width(width)) rd_st7_648  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[648]), .rdlo_in(a7_wr[652]),  .coef_in(coef[0]), .rdup_out(a8_wr[648]), .rdlo_out(a8_wr[652]));
			radix2 #(.width(width)) rd_st7_649  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[649]), .rdlo_in(a7_wr[653]),  .coef_in(coef[128]), .rdup_out(a8_wr[649]), .rdlo_out(a8_wr[653]));
			radix2 #(.width(width)) rd_st7_650  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[650]), .rdlo_in(a7_wr[654]),  .coef_in(coef[256]), .rdup_out(a8_wr[650]), .rdlo_out(a8_wr[654]));
			radix2 #(.width(width)) rd_st7_651  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[651]), .rdlo_in(a7_wr[655]),  .coef_in(coef[384]), .rdup_out(a8_wr[651]), .rdlo_out(a8_wr[655]));
			radix2 #(.width(width)) rd_st7_656  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[656]), .rdlo_in(a7_wr[660]),  .coef_in(coef[0]), .rdup_out(a8_wr[656]), .rdlo_out(a8_wr[660]));
			radix2 #(.width(width)) rd_st7_657  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[657]), .rdlo_in(a7_wr[661]),  .coef_in(coef[128]), .rdup_out(a8_wr[657]), .rdlo_out(a8_wr[661]));
			radix2 #(.width(width)) rd_st7_658  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[658]), .rdlo_in(a7_wr[662]),  .coef_in(coef[256]), .rdup_out(a8_wr[658]), .rdlo_out(a8_wr[662]));
			radix2 #(.width(width)) rd_st7_659  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[659]), .rdlo_in(a7_wr[663]),  .coef_in(coef[384]), .rdup_out(a8_wr[659]), .rdlo_out(a8_wr[663]));
			radix2 #(.width(width)) rd_st7_664  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[664]), .rdlo_in(a7_wr[668]),  .coef_in(coef[0]), .rdup_out(a8_wr[664]), .rdlo_out(a8_wr[668]));
			radix2 #(.width(width)) rd_st7_665  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[665]), .rdlo_in(a7_wr[669]),  .coef_in(coef[128]), .rdup_out(a8_wr[665]), .rdlo_out(a8_wr[669]));
			radix2 #(.width(width)) rd_st7_666  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[666]), .rdlo_in(a7_wr[670]),  .coef_in(coef[256]), .rdup_out(a8_wr[666]), .rdlo_out(a8_wr[670]));
			radix2 #(.width(width)) rd_st7_667  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[667]), .rdlo_in(a7_wr[671]),  .coef_in(coef[384]), .rdup_out(a8_wr[667]), .rdlo_out(a8_wr[671]));
			radix2 #(.width(width)) rd_st7_672  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[672]), .rdlo_in(a7_wr[676]),  .coef_in(coef[0]), .rdup_out(a8_wr[672]), .rdlo_out(a8_wr[676]));
			radix2 #(.width(width)) rd_st7_673  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[673]), .rdlo_in(a7_wr[677]),  .coef_in(coef[128]), .rdup_out(a8_wr[673]), .rdlo_out(a8_wr[677]));
			radix2 #(.width(width)) rd_st7_674  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[674]), .rdlo_in(a7_wr[678]),  .coef_in(coef[256]), .rdup_out(a8_wr[674]), .rdlo_out(a8_wr[678]));
			radix2 #(.width(width)) rd_st7_675  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[675]), .rdlo_in(a7_wr[679]),  .coef_in(coef[384]), .rdup_out(a8_wr[675]), .rdlo_out(a8_wr[679]));
			radix2 #(.width(width)) rd_st7_680  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[680]), .rdlo_in(a7_wr[684]),  .coef_in(coef[0]), .rdup_out(a8_wr[680]), .rdlo_out(a8_wr[684]));
			radix2 #(.width(width)) rd_st7_681  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[681]), .rdlo_in(a7_wr[685]),  .coef_in(coef[128]), .rdup_out(a8_wr[681]), .rdlo_out(a8_wr[685]));
			radix2 #(.width(width)) rd_st7_682  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[682]), .rdlo_in(a7_wr[686]),  .coef_in(coef[256]), .rdup_out(a8_wr[682]), .rdlo_out(a8_wr[686]));
			radix2 #(.width(width)) rd_st7_683  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[683]), .rdlo_in(a7_wr[687]),  .coef_in(coef[384]), .rdup_out(a8_wr[683]), .rdlo_out(a8_wr[687]));
			radix2 #(.width(width)) rd_st7_688  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[688]), .rdlo_in(a7_wr[692]),  .coef_in(coef[0]), .rdup_out(a8_wr[688]), .rdlo_out(a8_wr[692]));
			radix2 #(.width(width)) rd_st7_689  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[689]), .rdlo_in(a7_wr[693]),  .coef_in(coef[128]), .rdup_out(a8_wr[689]), .rdlo_out(a8_wr[693]));
			radix2 #(.width(width)) rd_st7_690  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[690]), .rdlo_in(a7_wr[694]),  .coef_in(coef[256]), .rdup_out(a8_wr[690]), .rdlo_out(a8_wr[694]));
			radix2 #(.width(width)) rd_st7_691  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[691]), .rdlo_in(a7_wr[695]),  .coef_in(coef[384]), .rdup_out(a8_wr[691]), .rdlo_out(a8_wr[695]));
			radix2 #(.width(width)) rd_st7_696  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[696]), .rdlo_in(a7_wr[700]),  .coef_in(coef[0]), .rdup_out(a8_wr[696]), .rdlo_out(a8_wr[700]));
			radix2 #(.width(width)) rd_st7_697  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[697]), .rdlo_in(a7_wr[701]),  .coef_in(coef[128]), .rdup_out(a8_wr[697]), .rdlo_out(a8_wr[701]));
			radix2 #(.width(width)) rd_st7_698  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[698]), .rdlo_in(a7_wr[702]),  .coef_in(coef[256]), .rdup_out(a8_wr[698]), .rdlo_out(a8_wr[702]));
			radix2 #(.width(width)) rd_st7_699  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[699]), .rdlo_in(a7_wr[703]),  .coef_in(coef[384]), .rdup_out(a8_wr[699]), .rdlo_out(a8_wr[703]));
			radix2 #(.width(width)) rd_st7_704  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[704]), .rdlo_in(a7_wr[708]),  .coef_in(coef[0]), .rdup_out(a8_wr[704]), .rdlo_out(a8_wr[708]));
			radix2 #(.width(width)) rd_st7_705  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[705]), .rdlo_in(a7_wr[709]),  .coef_in(coef[128]), .rdup_out(a8_wr[705]), .rdlo_out(a8_wr[709]));
			radix2 #(.width(width)) rd_st7_706  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[706]), .rdlo_in(a7_wr[710]),  .coef_in(coef[256]), .rdup_out(a8_wr[706]), .rdlo_out(a8_wr[710]));
			radix2 #(.width(width)) rd_st7_707  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[707]), .rdlo_in(a7_wr[711]),  .coef_in(coef[384]), .rdup_out(a8_wr[707]), .rdlo_out(a8_wr[711]));
			radix2 #(.width(width)) rd_st7_712  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[712]), .rdlo_in(a7_wr[716]),  .coef_in(coef[0]), .rdup_out(a8_wr[712]), .rdlo_out(a8_wr[716]));
			radix2 #(.width(width)) rd_st7_713  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[713]), .rdlo_in(a7_wr[717]),  .coef_in(coef[128]), .rdup_out(a8_wr[713]), .rdlo_out(a8_wr[717]));
			radix2 #(.width(width)) rd_st7_714  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[714]), .rdlo_in(a7_wr[718]),  .coef_in(coef[256]), .rdup_out(a8_wr[714]), .rdlo_out(a8_wr[718]));
			radix2 #(.width(width)) rd_st7_715  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[715]), .rdlo_in(a7_wr[719]),  .coef_in(coef[384]), .rdup_out(a8_wr[715]), .rdlo_out(a8_wr[719]));
			radix2 #(.width(width)) rd_st7_720  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[720]), .rdlo_in(a7_wr[724]),  .coef_in(coef[0]), .rdup_out(a8_wr[720]), .rdlo_out(a8_wr[724]));
			radix2 #(.width(width)) rd_st7_721  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[721]), .rdlo_in(a7_wr[725]),  .coef_in(coef[128]), .rdup_out(a8_wr[721]), .rdlo_out(a8_wr[725]));
			radix2 #(.width(width)) rd_st7_722  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[722]), .rdlo_in(a7_wr[726]),  .coef_in(coef[256]), .rdup_out(a8_wr[722]), .rdlo_out(a8_wr[726]));
			radix2 #(.width(width)) rd_st7_723  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[723]), .rdlo_in(a7_wr[727]),  .coef_in(coef[384]), .rdup_out(a8_wr[723]), .rdlo_out(a8_wr[727]));
			radix2 #(.width(width)) rd_st7_728  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[728]), .rdlo_in(a7_wr[732]),  .coef_in(coef[0]), .rdup_out(a8_wr[728]), .rdlo_out(a8_wr[732]));
			radix2 #(.width(width)) rd_st7_729  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[729]), .rdlo_in(a7_wr[733]),  .coef_in(coef[128]), .rdup_out(a8_wr[729]), .rdlo_out(a8_wr[733]));
			radix2 #(.width(width)) rd_st7_730  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[730]), .rdlo_in(a7_wr[734]),  .coef_in(coef[256]), .rdup_out(a8_wr[730]), .rdlo_out(a8_wr[734]));
			radix2 #(.width(width)) rd_st7_731  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[731]), .rdlo_in(a7_wr[735]),  .coef_in(coef[384]), .rdup_out(a8_wr[731]), .rdlo_out(a8_wr[735]));
			radix2 #(.width(width)) rd_st7_736  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[736]), .rdlo_in(a7_wr[740]),  .coef_in(coef[0]), .rdup_out(a8_wr[736]), .rdlo_out(a8_wr[740]));
			radix2 #(.width(width)) rd_st7_737  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[737]), .rdlo_in(a7_wr[741]),  .coef_in(coef[128]), .rdup_out(a8_wr[737]), .rdlo_out(a8_wr[741]));
			radix2 #(.width(width)) rd_st7_738  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[738]), .rdlo_in(a7_wr[742]),  .coef_in(coef[256]), .rdup_out(a8_wr[738]), .rdlo_out(a8_wr[742]));
			radix2 #(.width(width)) rd_st7_739  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[739]), .rdlo_in(a7_wr[743]),  .coef_in(coef[384]), .rdup_out(a8_wr[739]), .rdlo_out(a8_wr[743]));
			radix2 #(.width(width)) rd_st7_744  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[744]), .rdlo_in(a7_wr[748]),  .coef_in(coef[0]), .rdup_out(a8_wr[744]), .rdlo_out(a8_wr[748]));
			radix2 #(.width(width)) rd_st7_745  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[745]), .rdlo_in(a7_wr[749]),  .coef_in(coef[128]), .rdup_out(a8_wr[745]), .rdlo_out(a8_wr[749]));
			radix2 #(.width(width)) rd_st7_746  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[746]), .rdlo_in(a7_wr[750]),  .coef_in(coef[256]), .rdup_out(a8_wr[746]), .rdlo_out(a8_wr[750]));
			radix2 #(.width(width)) rd_st7_747  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[747]), .rdlo_in(a7_wr[751]),  .coef_in(coef[384]), .rdup_out(a8_wr[747]), .rdlo_out(a8_wr[751]));
			radix2 #(.width(width)) rd_st7_752  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[752]), .rdlo_in(a7_wr[756]),  .coef_in(coef[0]), .rdup_out(a8_wr[752]), .rdlo_out(a8_wr[756]));
			radix2 #(.width(width)) rd_st7_753  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[753]), .rdlo_in(a7_wr[757]),  .coef_in(coef[128]), .rdup_out(a8_wr[753]), .rdlo_out(a8_wr[757]));
			radix2 #(.width(width)) rd_st7_754  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[754]), .rdlo_in(a7_wr[758]),  .coef_in(coef[256]), .rdup_out(a8_wr[754]), .rdlo_out(a8_wr[758]));
			radix2 #(.width(width)) rd_st7_755  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[755]), .rdlo_in(a7_wr[759]),  .coef_in(coef[384]), .rdup_out(a8_wr[755]), .rdlo_out(a8_wr[759]));
			radix2 #(.width(width)) rd_st7_760  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[760]), .rdlo_in(a7_wr[764]),  .coef_in(coef[0]), .rdup_out(a8_wr[760]), .rdlo_out(a8_wr[764]));
			radix2 #(.width(width)) rd_st7_761  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[761]), .rdlo_in(a7_wr[765]),  .coef_in(coef[128]), .rdup_out(a8_wr[761]), .rdlo_out(a8_wr[765]));
			radix2 #(.width(width)) rd_st7_762  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[762]), .rdlo_in(a7_wr[766]),  .coef_in(coef[256]), .rdup_out(a8_wr[762]), .rdlo_out(a8_wr[766]));
			radix2 #(.width(width)) rd_st7_763  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[763]), .rdlo_in(a7_wr[767]),  .coef_in(coef[384]), .rdup_out(a8_wr[763]), .rdlo_out(a8_wr[767]));
			radix2 #(.width(width)) rd_st7_768  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[768]), .rdlo_in(a7_wr[772]),  .coef_in(coef[0]), .rdup_out(a8_wr[768]), .rdlo_out(a8_wr[772]));
			radix2 #(.width(width)) rd_st7_769  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[769]), .rdlo_in(a7_wr[773]),  .coef_in(coef[128]), .rdup_out(a8_wr[769]), .rdlo_out(a8_wr[773]));
			radix2 #(.width(width)) rd_st7_770  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[770]), .rdlo_in(a7_wr[774]),  .coef_in(coef[256]), .rdup_out(a8_wr[770]), .rdlo_out(a8_wr[774]));
			radix2 #(.width(width)) rd_st7_771  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[771]), .rdlo_in(a7_wr[775]),  .coef_in(coef[384]), .rdup_out(a8_wr[771]), .rdlo_out(a8_wr[775]));
			radix2 #(.width(width)) rd_st7_776  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[776]), .rdlo_in(a7_wr[780]),  .coef_in(coef[0]), .rdup_out(a8_wr[776]), .rdlo_out(a8_wr[780]));
			radix2 #(.width(width)) rd_st7_777  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[777]), .rdlo_in(a7_wr[781]),  .coef_in(coef[128]), .rdup_out(a8_wr[777]), .rdlo_out(a8_wr[781]));
			radix2 #(.width(width)) rd_st7_778  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[778]), .rdlo_in(a7_wr[782]),  .coef_in(coef[256]), .rdup_out(a8_wr[778]), .rdlo_out(a8_wr[782]));
			radix2 #(.width(width)) rd_st7_779  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[779]), .rdlo_in(a7_wr[783]),  .coef_in(coef[384]), .rdup_out(a8_wr[779]), .rdlo_out(a8_wr[783]));
			radix2 #(.width(width)) rd_st7_784  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[784]), .rdlo_in(a7_wr[788]),  .coef_in(coef[0]), .rdup_out(a8_wr[784]), .rdlo_out(a8_wr[788]));
			radix2 #(.width(width)) rd_st7_785  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[785]), .rdlo_in(a7_wr[789]),  .coef_in(coef[128]), .rdup_out(a8_wr[785]), .rdlo_out(a8_wr[789]));
			radix2 #(.width(width)) rd_st7_786  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[786]), .rdlo_in(a7_wr[790]),  .coef_in(coef[256]), .rdup_out(a8_wr[786]), .rdlo_out(a8_wr[790]));
			radix2 #(.width(width)) rd_st7_787  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[787]), .rdlo_in(a7_wr[791]),  .coef_in(coef[384]), .rdup_out(a8_wr[787]), .rdlo_out(a8_wr[791]));
			radix2 #(.width(width)) rd_st7_792  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[792]), .rdlo_in(a7_wr[796]),  .coef_in(coef[0]), .rdup_out(a8_wr[792]), .rdlo_out(a8_wr[796]));
			radix2 #(.width(width)) rd_st7_793  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[793]), .rdlo_in(a7_wr[797]),  .coef_in(coef[128]), .rdup_out(a8_wr[793]), .rdlo_out(a8_wr[797]));
			radix2 #(.width(width)) rd_st7_794  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[794]), .rdlo_in(a7_wr[798]),  .coef_in(coef[256]), .rdup_out(a8_wr[794]), .rdlo_out(a8_wr[798]));
			radix2 #(.width(width)) rd_st7_795  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[795]), .rdlo_in(a7_wr[799]),  .coef_in(coef[384]), .rdup_out(a8_wr[795]), .rdlo_out(a8_wr[799]));
			radix2 #(.width(width)) rd_st7_800  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[800]), .rdlo_in(a7_wr[804]),  .coef_in(coef[0]), .rdup_out(a8_wr[800]), .rdlo_out(a8_wr[804]));
			radix2 #(.width(width)) rd_st7_801  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[801]), .rdlo_in(a7_wr[805]),  .coef_in(coef[128]), .rdup_out(a8_wr[801]), .rdlo_out(a8_wr[805]));
			radix2 #(.width(width)) rd_st7_802  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[802]), .rdlo_in(a7_wr[806]),  .coef_in(coef[256]), .rdup_out(a8_wr[802]), .rdlo_out(a8_wr[806]));
			radix2 #(.width(width)) rd_st7_803  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[803]), .rdlo_in(a7_wr[807]),  .coef_in(coef[384]), .rdup_out(a8_wr[803]), .rdlo_out(a8_wr[807]));
			radix2 #(.width(width)) rd_st7_808  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[808]), .rdlo_in(a7_wr[812]),  .coef_in(coef[0]), .rdup_out(a8_wr[808]), .rdlo_out(a8_wr[812]));
			radix2 #(.width(width)) rd_st7_809  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[809]), .rdlo_in(a7_wr[813]),  .coef_in(coef[128]), .rdup_out(a8_wr[809]), .rdlo_out(a8_wr[813]));
			radix2 #(.width(width)) rd_st7_810  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[810]), .rdlo_in(a7_wr[814]),  .coef_in(coef[256]), .rdup_out(a8_wr[810]), .rdlo_out(a8_wr[814]));
			radix2 #(.width(width)) rd_st7_811  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[811]), .rdlo_in(a7_wr[815]),  .coef_in(coef[384]), .rdup_out(a8_wr[811]), .rdlo_out(a8_wr[815]));
			radix2 #(.width(width)) rd_st7_816  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[816]), .rdlo_in(a7_wr[820]),  .coef_in(coef[0]), .rdup_out(a8_wr[816]), .rdlo_out(a8_wr[820]));
			radix2 #(.width(width)) rd_st7_817  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[817]), .rdlo_in(a7_wr[821]),  .coef_in(coef[128]), .rdup_out(a8_wr[817]), .rdlo_out(a8_wr[821]));
			radix2 #(.width(width)) rd_st7_818  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[818]), .rdlo_in(a7_wr[822]),  .coef_in(coef[256]), .rdup_out(a8_wr[818]), .rdlo_out(a8_wr[822]));
			radix2 #(.width(width)) rd_st7_819  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[819]), .rdlo_in(a7_wr[823]),  .coef_in(coef[384]), .rdup_out(a8_wr[819]), .rdlo_out(a8_wr[823]));
			radix2 #(.width(width)) rd_st7_824  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[824]), .rdlo_in(a7_wr[828]),  .coef_in(coef[0]), .rdup_out(a8_wr[824]), .rdlo_out(a8_wr[828]));
			radix2 #(.width(width)) rd_st7_825  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[825]), .rdlo_in(a7_wr[829]),  .coef_in(coef[128]), .rdup_out(a8_wr[825]), .rdlo_out(a8_wr[829]));
			radix2 #(.width(width)) rd_st7_826  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[826]), .rdlo_in(a7_wr[830]),  .coef_in(coef[256]), .rdup_out(a8_wr[826]), .rdlo_out(a8_wr[830]));
			radix2 #(.width(width)) rd_st7_827  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[827]), .rdlo_in(a7_wr[831]),  .coef_in(coef[384]), .rdup_out(a8_wr[827]), .rdlo_out(a8_wr[831]));
			radix2 #(.width(width)) rd_st7_832  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[832]), .rdlo_in(a7_wr[836]),  .coef_in(coef[0]), .rdup_out(a8_wr[832]), .rdlo_out(a8_wr[836]));
			radix2 #(.width(width)) rd_st7_833  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[833]), .rdlo_in(a7_wr[837]),  .coef_in(coef[128]), .rdup_out(a8_wr[833]), .rdlo_out(a8_wr[837]));
			radix2 #(.width(width)) rd_st7_834  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[834]), .rdlo_in(a7_wr[838]),  .coef_in(coef[256]), .rdup_out(a8_wr[834]), .rdlo_out(a8_wr[838]));
			radix2 #(.width(width)) rd_st7_835  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[835]), .rdlo_in(a7_wr[839]),  .coef_in(coef[384]), .rdup_out(a8_wr[835]), .rdlo_out(a8_wr[839]));
			radix2 #(.width(width)) rd_st7_840  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[840]), .rdlo_in(a7_wr[844]),  .coef_in(coef[0]), .rdup_out(a8_wr[840]), .rdlo_out(a8_wr[844]));
			radix2 #(.width(width)) rd_st7_841  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[841]), .rdlo_in(a7_wr[845]),  .coef_in(coef[128]), .rdup_out(a8_wr[841]), .rdlo_out(a8_wr[845]));
			radix2 #(.width(width)) rd_st7_842  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[842]), .rdlo_in(a7_wr[846]),  .coef_in(coef[256]), .rdup_out(a8_wr[842]), .rdlo_out(a8_wr[846]));
			radix2 #(.width(width)) rd_st7_843  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[843]), .rdlo_in(a7_wr[847]),  .coef_in(coef[384]), .rdup_out(a8_wr[843]), .rdlo_out(a8_wr[847]));
			radix2 #(.width(width)) rd_st7_848  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[848]), .rdlo_in(a7_wr[852]),  .coef_in(coef[0]), .rdup_out(a8_wr[848]), .rdlo_out(a8_wr[852]));
			radix2 #(.width(width)) rd_st7_849  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[849]), .rdlo_in(a7_wr[853]),  .coef_in(coef[128]), .rdup_out(a8_wr[849]), .rdlo_out(a8_wr[853]));
			radix2 #(.width(width)) rd_st7_850  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[850]), .rdlo_in(a7_wr[854]),  .coef_in(coef[256]), .rdup_out(a8_wr[850]), .rdlo_out(a8_wr[854]));
			radix2 #(.width(width)) rd_st7_851  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[851]), .rdlo_in(a7_wr[855]),  .coef_in(coef[384]), .rdup_out(a8_wr[851]), .rdlo_out(a8_wr[855]));
			radix2 #(.width(width)) rd_st7_856  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[856]), .rdlo_in(a7_wr[860]),  .coef_in(coef[0]), .rdup_out(a8_wr[856]), .rdlo_out(a8_wr[860]));
			radix2 #(.width(width)) rd_st7_857  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[857]), .rdlo_in(a7_wr[861]),  .coef_in(coef[128]), .rdup_out(a8_wr[857]), .rdlo_out(a8_wr[861]));
			radix2 #(.width(width)) rd_st7_858  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[858]), .rdlo_in(a7_wr[862]),  .coef_in(coef[256]), .rdup_out(a8_wr[858]), .rdlo_out(a8_wr[862]));
			radix2 #(.width(width)) rd_st7_859  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[859]), .rdlo_in(a7_wr[863]),  .coef_in(coef[384]), .rdup_out(a8_wr[859]), .rdlo_out(a8_wr[863]));
			radix2 #(.width(width)) rd_st7_864  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[864]), .rdlo_in(a7_wr[868]),  .coef_in(coef[0]), .rdup_out(a8_wr[864]), .rdlo_out(a8_wr[868]));
			radix2 #(.width(width)) rd_st7_865  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[865]), .rdlo_in(a7_wr[869]),  .coef_in(coef[128]), .rdup_out(a8_wr[865]), .rdlo_out(a8_wr[869]));
			radix2 #(.width(width)) rd_st7_866  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[866]), .rdlo_in(a7_wr[870]),  .coef_in(coef[256]), .rdup_out(a8_wr[866]), .rdlo_out(a8_wr[870]));
			radix2 #(.width(width)) rd_st7_867  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[867]), .rdlo_in(a7_wr[871]),  .coef_in(coef[384]), .rdup_out(a8_wr[867]), .rdlo_out(a8_wr[871]));
			radix2 #(.width(width)) rd_st7_872  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[872]), .rdlo_in(a7_wr[876]),  .coef_in(coef[0]), .rdup_out(a8_wr[872]), .rdlo_out(a8_wr[876]));
			radix2 #(.width(width)) rd_st7_873  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[873]), .rdlo_in(a7_wr[877]),  .coef_in(coef[128]), .rdup_out(a8_wr[873]), .rdlo_out(a8_wr[877]));
			radix2 #(.width(width)) rd_st7_874  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[874]), .rdlo_in(a7_wr[878]),  .coef_in(coef[256]), .rdup_out(a8_wr[874]), .rdlo_out(a8_wr[878]));
			radix2 #(.width(width)) rd_st7_875  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[875]), .rdlo_in(a7_wr[879]),  .coef_in(coef[384]), .rdup_out(a8_wr[875]), .rdlo_out(a8_wr[879]));
			radix2 #(.width(width)) rd_st7_880  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[880]), .rdlo_in(a7_wr[884]),  .coef_in(coef[0]), .rdup_out(a8_wr[880]), .rdlo_out(a8_wr[884]));
			radix2 #(.width(width)) rd_st7_881  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[881]), .rdlo_in(a7_wr[885]),  .coef_in(coef[128]), .rdup_out(a8_wr[881]), .rdlo_out(a8_wr[885]));
			radix2 #(.width(width)) rd_st7_882  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[882]), .rdlo_in(a7_wr[886]),  .coef_in(coef[256]), .rdup_out(a8_wr[882]), .rdlo_out(a8_wr[886]));
			radix2 #(.width(width)) rd_st7_883  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[883]), .rdlo_in(a7_wr[887]),  .coef_in(coef[384]), .rdup_out(a8_wr[883]), .rdlo_out(a8_wr[887]));
			radix2 #(.width(width)) rd_st7_888  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[888]), .rdlo_in(a7_wr[892]),  .coef_in(coef[0]), .rdup_out(a8_wr[888]), .rdlo_out(a8_wr[892]));
			radix2 #(.width(width)) rd_st7_889  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[889]), .rdlo_in(a7_wr[893]),  .coef_in(coef[128]), .rdup_out(a8_wr[889]), .rdlo_out(a8_wr[893]));
			radix2 #(.width(width)) rd_st7_890  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[890]), .rdlo_in(a7_wr[894]),  .coef_in(coef[256]), .rdup_out(a8_wr[890]), .rdlo_out(a8_wr[894]));
			radix2 #(.width(width)) rd_st7_891  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[891]), .rdlo_in(a7_wr[895]),  .coef_in(coef[384]), .rdup_out(a8_wr[891]), .rdlo_out(a8_wr[895]));
			radix2 #(.width(width)) rd_st7_896  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[896]), .rdlo_in(a7_wr[900]),  .coef_in(coef[0]), .rdup_out(a8_wr[896]), .rdlo_out(a8_wr[900]));
			radix2 #(.width(width)) rd_st7_897  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[897]), .rdlo_in(a7_wr[901]),  .coef_in(coef[128]), .rdup_out(a8_wr[897]), .rdlo_out(a8_wr[901]));
			radix2 #(.width(width)) rd_st7_898  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[898]), .rdlo_in(a7_wr[902]),  .coef_in(coef[256]), .rdup_out(a8_wr[898]), .rdlo_out(a8_wr[902]));
			radix2 #(.width(width)) rd_st7_899  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[899]), .rdlo_in(a7_wr[903]),  .coef_in(coef[384]), .rdup_out(a8_wr[899]), .rdlo_out(a8_wr[903]));
			radix2 #(.width(width)) rd_st7_904  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[904]), .rdlo_in(a7_wr[908]),  .coef_in(coef[0]), .rdup_out(a8_wr[904]), .rdlo_out(a8_wr[908]));
			radix2 #(.width(width)) rd_st7_905  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[905]), .rdlo_in(a7_wr[909]),  .coef_in(coef[128]), .rdup_out(a8_wr[905]), .rdlo_out(a8_wr[909]));
			radix2 #(.width(width)) rd_st7_906  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[906]), .rdlo_in(a7_wr[910]),  .coef_in(coef[256]), .rdup_out(a8_wr[906]), .rdlo_out(a8_wr[910]));
			radix2 #(.width(width)) rd_st7_907  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[907]), .rdlo_in(a7_wr[911]),  .coef_in(coef[384]), .rdup_out(a8_wr[907]), .rdlo_out(a8_wr[911]));
			radix2 #(.width(width)) rd_st7_912  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[912]), .rdlo_in(a7_wr[916]),  .coef_in(coef[0]), .rdup_out(a8_wr[912]), .rdlo_out(a8_wr[916]));
			radix2 #(.width(width)) rd_st7_913  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[913]), .rdlo_in(a7_wr[917]),  .coef_in(coef[128]), .rdup_out(a8_wr[913]), .rdlo_out(a8_wr[917]));
			radix2 #(.width(width)) rd_st7_914  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[914]), .rdlo_in(a7_wr[918]),  .coef_in(coef[256]), .rdup_out(a8_wr[914]), .rdlo_out(a8_wr[918]));
			radix2 #(.width(width)) rd_st7_915  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[915]), .rdlo_in(a7_wr[919]),  .coef_in(coef[384]), .rdup_out(a8_wr[915]), .rdlo_out(a8_wr[919]));
			radix2 #(.width(width)) rd_st7_920  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[920]), .rdlo_in(a7_wr[924]),  .coef_in(coef[0]), .rdup_out(a8_wr[920]), .rdlo_out(a8_wr[924]));
			radix2 #(.width(width)) rd_st7_921  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[921]), .rdlo_in(a7_wr[925]),  .coef_in(coef[128]), .rdup_out(a8_wr[921]), .rdlo_out(a8_wr[925]));
			radix2 #(.width(width)) rd_st7_922  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[922]), .rdlo_in(a7_wr[926]),  .coef_in(coef[256]), .rdup_out(a8_wr[922]), .rdlo_out(a8_wr[926]));
			radix2 #(.width(width)) rd_st7_923  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[923]), .rdlo_in(a7_wr[927]),  .coef_in(coef[384]), .rdup_out(a8_wr[923]), .rdlo_out(a8_wr[927]));
			radix2 #(.width(width)) rd_st7_928  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[928]), .rdlo_in(a7_wr[932]),  .coef_in(coef[0]), .rdup_out(a8_wr[928]), .rdlo_out(a8_wr[932]));
			radix2 #(.width(width)) rd_st7_929  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[929]), .rdlo_in(a7_wr[933]),  .coef_in(coef[128]), .rdup_out(a8_wr[929]), .rdlo_out(a8_wr[933]));
			radix2 #(.width(width)) rd_st7_930  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[930]), .rdlo_in(a7_wr[934]),  .coef_in(coef[256]), .rdup_out(a8_wr[930]), .rdlo_out(a8_wr[934]));
			radix2 #(.width(width)) rd_st7_931  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[931]), .rdlo_in(a7_wr[935]),  .coef_in(coef[384]), .rdup_out(a8_wr[931]), .rdlo_out(a8_wr[935]));
			radix2 #(.width(width)) rd_st7_936  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[936]), .rdlo_in(a7_wr[940]),  .coef_in(coef[0]), .rdup_out(a8_wr[936]), .rdlo_out(a8_wr[940]));
			radix2 #(.width(width)) rd_st7_937  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[937]), .rdlo_in(a7_wr[941]),  .coef_in(coef[128]), .rdup_out(a8_wr[937]), .rdlo_out(a8_wr[941]));
			radix2 #(.width(width)) rd_st7_938  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[938]), .rdlo_in(a7_wr[942]),  .coef_in(coef[256]), .rdup_out(a8_wr[938]), .rdlo_out(a8_wr[942]));
			radix2 #(.width(width)) rd_st7_939  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[939]), .rdlo_in(a7_wr[943]),  .coef_in(coef[384]), .rdup_out(a8_wr[939]), .rdlo_out(a8_wr[943]));
			radix2 #(.width(width)) rd_st7_944  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[944]), .rdlo_in(a7_wr[948]),  .coef_in(coef[0]), .rdup_out(a8_wr[944]), .rdlo_out(a8_wr[948]));
			radix2 #(.width(width)) rd_st7_945  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[945]), .rdlo_in(a7_wr[949]),  .coef_in(coef[128]), .rdup_out(a8_wr[945]), .rdlo_out(a8_wr[949]));
			radix2 #(.width(width)) rd_st7_946  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[946]), .rdlo_in(a7_wr[950]),  .coef_in(coef[256]), .rdup_out(a8_wr[946]), .rdlo_out(a8_wr[950]));
			radix2 #(.width(width)) rd_st7_947  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[947]), .rdlo_in(a7_wr[951]),  .coef_in(coef[384]), .rdup_out(a8_wr[947]), .rdlo_out(a8_wr[951]));
			radix2 #(.width(width)) rd_st7_952  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[952]), .rdlo_in(a7_wr[956]),  .coef_in(coef[0]), .rdup_out(a8_wr[952]), .rdlo_out(a8_wr[956]));
			radix2 #(.width(width)) rd_st7_953  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[953]), .rdlo_in(a7_wr[957]),  .coef_in(coef[128]), .rdup_out(a8_wr[953]), .rdlo_out(a8_wr[957]));
			radix2 #(.width(width)) rd_st7_954  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[954]), .rdlo_in(a7_wr[958]),  .coef_in(coef[256]), .rdup_out(a8_wr[954]), .rdlo_out(a8_wr[958]));
			radix2 #(.width(width)) rd_st7_955  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[955]), .rdlo_in(a7_wr[959]),  .coef_in(coef[384]), .rdup_out(a8_wr[955]), .rdlo_out(a8_wr[959]));
			radix2 #(.width(width)) rd_st7_960  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[960]), .rdlo_in(a7_wr[964]),  .coef_in(coef[0]), .rdup_out(a8_wr[960]), .rdlo_out(a8_wr[964]));
			radix2 #(.width(width)) rd_st7_961  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[961]), .rdlo_in(a7_wr[965]),  .coef_in(coef[128]), .rdup_out(a8_wr[961]), .rdlo_out(a8_wr[965]));
			radix2 #(.width(width)) rd_st7_962  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[962]), .rdlo_in(a7_wr[966]),  .coef_in(coef[256]), .rdup_out(a8_wr[962]), .rdlo_out(a8_wr[966]));
			radix2 #(.width(width)) rd_st7_963  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[963]), .rdlo_in(a7_wr[967]),  .coef_in(coef[384]), .rdup_out(a8_wr[963]), .rdlo_out(a8_wr[967]));
			radix2 #(.width(width)) rd_st7_968  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[968]), .rdlo_in(a7_wr[972]),  .coef_in(coef[0]), .rdup_out(a8_wr[968]), .rdlo_out(a8_wr[972]));
			radix2 #(.width(width)) rd_st7_969  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[969]), .rdlo_in(a7_wr[973]),  .coef_in(coef[128]), .rdup_out(a8_wr[969]), .rdlo_out(a8_wr[973]));
			radix2 #(.width(width)) rd_st7_970  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[970]), .rdlo_in(a7_wr[974]),  .coef_in(coef[256]), .rdup_out(a8_wr[970]), .rdlo_out(a8_wr[974]));
			radix2 #(.width(width)) rd_st7_971  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[971]), .rdlo_in(a7_wr[975]),  .coef_in(coef[384]), .rdup_out(a8_wr[971]), .rdlo_out(a8_wr[975]));
			radix2 #(.width(width)) rd_st7_976  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[976]), .rdlo_in(a7_wr[980]),  .coef_in(coef[0]), .rdup_out(a8_wr[976]), .rdlo_out(a8_wr[980]));
			radix2 #(.width(width)) rd_st7_977  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[977]), .rdlo_in(a7_wr[981]),  .coef_in(coef[128]), .rdup_out(a8_wr[977]), .rdlo_out(a8_wr[981]));
			radix2 #(.width(width)) rd_st7_978  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[978]), .rdlo_in(a7_wr[982]),  .coef_in(coef[256]), .rdup_out(a8_wr[978]), .rdlo_out(a8_wr[982]));
			radix2 #(.width(width)) rd_st7_979  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[979]), .rdlo_in(a7_wr[983]),  .coef_in(coef[384]), .rdup_out(a8_wr[979]), .rdlo_out(a8_wr[983]));
			radix2 #(.width(width)) rd_st7_984  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[984]), .rdlo_in(a7_wr[988]),  .coef_in(coef[0]), .rdup_out(a8_wr[984]), .rdlo_out(a8_wr[988]));
			radix2 #(.width(width)) rd_st7_985  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[985]), .rdlo_in(a7_wr[989]),  .coef_in(coef[128]), .rdup_out(a8_wr[985]), .rdlo_out(a8_wr[989]));
			radix2 #(.width(width)) rd_st7_986  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[986]), .rdlo_in(a7_wr[990]),  .coef_in(coef[256]), .rdup_out(a8_wr[986]), .rdlo_out(a8_wr[990]));
			radix2 #(.width(width)) rd_st7_987  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[987]), .rdlo_in(a7_wr[991]),  .coef_in(coef[384]), .rdup_out(a8_wr[987]), .rdlo_out(a8_wr[991]));
			radix2 #(.width(width)) rd_st7_992  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[992]), .rdlo_in(a7_wr[996]),  .coef_in(coef[0]), .rdup_out(a8_wr[992]), .rdlo_out(a8_wr[996]));
			radix2 #(.width(width)) rd_st7_993  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[993]), .rdlo_in(a7_wr[997]),  .coef_in(coef[128]), .rdup_out(a8_wr[993]), .rdlo_out(a8_wr[997]));
			radix2 #(.width(width)) rd_st7_994  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[994]), .rdlo_in(a7_wr[998]),  .coef_in(coef[256]), .rdup_out(a8_wr[994]), .rdlo_out(a8_wr[998]));
			radix2 #(.width(width)) rd_st7_995  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[995]), .rdlo_in(a7_wr[999]),  .coef_in(coef[384]), .rdup_out(a8_wr[995]), .rdlo_out(a8_wr[999]));
			radix2 #(.width(width)) rd_st7_1000  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1000]), .rdlo_in(a7_wr[1004]),  .coef_in(coef[0]), .rdup_out(a8_wr[1000]), .rdlo_out(a8_wr[1004]));
			radix2 #(.width(width)) rd_st7_1001  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1001]), .rdlo_in(a7_wr[1005]),  .coef_in(coef[128]), .rdup_out(a8_wr[1001]), .rdlo_out(a8_wr[1005]));
			radix2 #(.width(width)) rd_st7_1002  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1002]), .rdlo_in(a7_wr[1006]),  .coef_in(coef[256]), .rdup_out(a8_wr[1002]), .rdlo_out(a8_wr[1006]));
			radix2 #(.width(width)) rd_st7_1003  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1003]), .rdlo_in(a7_wr[1007]),  .coef_in(coef[384]), .rdup_out(a8_wr[1003]), .rdlo_out(a8_wr[1007]));
			radix2 #(.width(width)) rd_st7_1008  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1008]), .rdlo_in(a7_wr[1012]),  .coef_in(coef[0]), .rdup_out(a8_wr[1008]), .rdlo_out(a8_wr[1012]));
			radix2 #(.width(width)) rd_st7_1009  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1009]), .rdlo_in(a7_wr[1013]),  .coef_in(coef[128]), .rdup_out(a8_wr[1009]), .rdlo_out(a8_wr[1013]));
			radix2 #(.width(width)) rd_st7_1010  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1010]), .rdlo_in(a7_wr[1014]),  .coef_in(coef[256]), .rdup_out(a8_wr[1010]), .rdlo_out(a8_wr[1014]));
			radix2 #(.width(width)) rd_st7_1011  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1011]), .rdlo_in(a7_wr[1015]),  .coef_in(coef[384]), .rdup_out(a8_wr[1011]), .rdlo_out(a8_wr[1015]));
			radix2 #(.width(width)) rd_st7_1016  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1016]), .rdlo_in(a7_wr[1020]),  .coef_in(coef[0]), .rdup_out(a8_wr[1016]), .rdlo_out(a8_wr[1020]));
			radix2 #(.width(width)) rd_st7_1017  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1017]), .rdlo_in(a7_wr[1021]),  .coef_in(coef[128]), .rdup_out(a8_wr[1017]), .rdlo_out(a8_wr[1021]));
			radix2 #(.width(width)) rd_st7_1018  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1018]), .rdlo_in(a7_wr[1022]),  .coef_in(coef[256]), .rdup_out(a8_wr[1018]), .rdlo_out(a8_wr[1022]));
			radix2 #(.width(width)) rd_st7_1019  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1019]), .rdlo_in(a7_wr[1023]),  .coef_in(coef[384]), .rdup_out(a8_wr[1019]), .rdlo_out(a8_wr[1023]));

		//--- radix stage 8
			radix2 #(.width(width)) rd_st8_0   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[0]), .rdlo_in(a8_wr[2]),  .coef_in(coef[0]), .rdup_out(a9_wr[0]), .rdlo_out(a9_wr[2]));
			radix2 #(.width(width)) rd_st8_1   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1]), .rdlo_in(a8_wr[3]),  .coef_in(coef[256]), .rdup_out(a9_wr[1]), .rdlo_out(a9_wr[3]));
			radix2 #(.width(width)) rd_st8_4   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[4]), .rdlo_in(a8_wr[6]),  .coef_in(coef[0]), .rdup_out(a9_wr[4]), .rdlo_out(a9_wr[6]));
			radix2 #(.width(width)) rd_st8_5   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[5]), .rdlo_in(a8_wr[7]),  .coef_in(coef[256]), .rdup_out(a9_wr[5]), .rdlo_out(a9_wr[7]));
			radix2 #(.width(width)) rd_st8_8   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[8]), .rdlo_in(a8_wr[10]),  .coef_in(coef[0]), .rdup_out(a9_wr[8]), .rdlo_out(a9_wr[10]));
			radix2 #(.width(width)) rd_st8_9   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[9]), .rdlo_in(a8_wr[11]),  .coef_in(coef[256]), .rdup_out(a9_wr[9]), .rdlo_out(a9_wr[11]));
			radix2 #(.width(width)) rd_st8_12  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[12]), .rdlo_in(a8_wr[14]),  .coef_in(coef[0]), .rdup_out(a9_wr[12]), .rdlo_out(a9_wr[14]));
			radix2 #(.width(width)) rd_st8_13  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[13]), .rdlo_in(a8_wr[15]),  .coef_in(coef[256]), .rdup_out(a9_wr[13]), .rdlo_out(a9_wr[15]));
			radix2 #(.width(width)) rd_st8_16  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[16]), .rdlo_in(a8_wr[18]),  .coef_in(coef[0]), .rdup_out(a9_wr[16]), .rdlo_out(a9_wr[18]));
			radix2 #(.width(width)) rd_st8_17  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[17]), .rdlo_in(a8_wr[19]),  .coef_in(coef[256]), .rdup_out(a9_wr[17]), .rdlo_out(a9_wr[19]));
			radix2 #(.width(width)) rd_st8_20  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[20]), .rdlo_in(a8_wr[22]),  .coef_in(coef[0]), .rdup_out(a9_wr[20]), .rdlo_out(a9_wr[22]));
			radix2 #(.width(width)) rd_st8_21  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[21]), .rdlo_in(a8_wr[23]),  .coef_in(coef[256]), .rdup_out(a9_wr[21]), .rdlo_out(a9_wr[23]));
			radix2 #(.width(width)) rd_st8_24  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[24]), .rdlo_in(a8_wr[26]),  .coef_in(coef[0]), .rdup_out(a9_wr[24]), .rdlo_out(a9_wr[26]));
			radix2 #(.width(width)) rd_st8_25  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[25]), .rdlo_in(a8_wr[27]),  .coef_in(coef[256]), .rdup_out(a9_wr[25]), .rdlo_out(a9_wr[27]));
			radix2 #(.width(width)) rd_st8_28  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[28]), .rdlo_in(a8_wr[30]),  .coef_in(coef[0]), .rdup_out(a9_wr[28]), .rdlo_out(a9_wr[30]));
			radix2 #(.width(width)) rd_st8_29  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[29]), .rdlo_in(a8_wr[31]),  .coef_in(coef[256]), .rdup_out(a9_wr[29]), .rdlo_out(a9_wr[31]));
			radix2 #(.width(width)) rd_st8_32  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[32]), .rdlo_in(a8_wr[34]),  .coef_in(coef[0]), .rdup_out(a9_wr[32]), .rdlo_out(a9_wr[34]));
			radix2 #(.width(width)) rd_st8_33  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[33]), .rdlo_in(a8_wr[35]),  .coef_in(coef[256]), .rdup_out(a9_wr[33]), .rdlo_out(a9_wr[35]));
			radix2 #(.width(width)) rd_st8_36  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[36]), .rdlo_in(a8_wr[38]),  .coef_in(coef[0]), .rdup_out(a9_wr[36]), .rdlo_out(a9_wr[38]));
			radix2 #(.width(width)) rd_st8_37  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[37]), .rdlo_in(a8_wr[39]),  .coef_in(coef[256]), .rdup_out(a9_wr[37]), .rdlo_out(a9_wr[39]));
			radix2 #(.width(width)) rd_st8_40  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[40]), .rdlo_in(a8_wr[42]),  .coef_in(coef[0]), .rdup_out(a9_wr[40]), .rdlo_out(a9_wr[42]));
			radix2 #(.width(width)) rd_st8_41  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[41]), .rdlo_in(a8_wr[43]),  .coef_in(coef[256]), .rdup_out(a9_wr[41]), .rdlo_out(a9_wr[43]));
			radix2 #(.width(width)) rd_st8_44  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[44]), .rdlo_in(a8_wr[46]),  .coef_in(coef[0]), .rdup_out(a9_wr[44]), .rdlo_out(a9_wr[46]));
			radix2 #(.width(width)) rd_st8_45  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[45]), .rdlo_in(a8_wr[47]),  .coef_in(coef[256]), .rdup_out(a9_wr[45]), .rdlo_out(a9_wr[47]));
			radix2 #(.width(width)) rd_st8_48  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[48]), .rdlo_in(a8_wr[50]),  .coef_in(coef[0]), .rdup_out(a9_wr[48]), .rdlo_out(a9_wr[50]));
			radix2 #(.width(width)) rd_st8_49  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[49]), .rdlo_in(a8_wr[51]),  .coef_in(coef[256]), .rdup_out(a9_wr[49]), .rdlo_out(a9_wr[51]));
			radix2 #(.width(width)) rd_st8_52  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[52]), .rdlo_in(a8_wr[54]),  .coef_in(coef[0]), .rdup_out(a9_wr[52]), .rdlo_out(a9_wr[54]));
			radix2 #(.width(width)) rd_st8_53  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[53]), .rdlo_in(a8_wr[55]),  .coef_in(coef[256]), .rdup_out(a9_wr[53]), .rdlo_out(a9_wr[55]));
			radix2 #(.width(width)) rd_st8_56  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[56]), .rdlo_in(a8_wr[58]),  .coef_in(coef[0]), .rdup_out(a9_wr[56]), .rdlo_out(a9_wr[58]));
			radix2 #(.width(width)) rd_st8_57  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[57]), .rdlo_in(a8_wr[59]),  .coef_in(coef[256]), .rdup_out(a9_wr[57]), .rdlo_out(a9_wr[59]));
			radix2 #(.width(width)) rd_st8_60  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[60]), .rdlo_in(a8_wr[62]),  .coef_in(coef[0]), .rdup_out(a9_wr[60]), .rdlo_out(a9_wr[62]));
			radix2 #(.width(width)) rd_st8_61  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[61]), .rdlo_in(a8_wr[63]),  .coef_in(coef[256]), .rdup_out(a9_wr[61]), .rdlo_out(a9_wr[63]));
			radix2 #(.width(width)) rd_st8_64  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[64]), .rdlo_in(a8_wr[66]),  .coef_in(coef[0]), .rdup_out(a9_wr[64]), .rdlo_out(a9_wr[66]));
			radix2 #(.width(width)) rd_st8_65  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[65]), .rdlo_in(a8_wr[67]),  .coef_in(coef[256]), .rdup_out(a9_wr[65]), .rdlo_out(a9_wr[67]));
			radix2 #(.width(width)) rd_st8_68  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[68]), .rdlo_in(a8_wr[70]),  .coef_in(coef[0]), .rdup_out(a9_wr[68]), .rdlo_out(a9_wr[70]));
			radix2 #(.width(width)) rd_st8_69  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[69]), .rdlo_in(a8_wr[71]),  .coef_in(coef[256]), .rdup_out(a9_wr[69]), .rdlo_out(a9_wr[71]));
			radix2 #(.width(width)) rd_st8_72  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[72]), .rdlo_in(a8_wr[74]),  .coef_in(coef[0]), .rdup_out(a9_wr[72]), .rdlo_out(a9_wr[74]));
			radix2 #(.width(width)) rd_st8_73  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[73]), .rdlo_in(a8_wr[75]),  .coef_in(coef[256]), .rdup_out(a9_wr[73]), .rdlo_out(a9_wr[75]));
			radix2 #(.width(width)) rd_st8_76  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[76]), .rdlo_in(a8_wr[78]),  .coef_in(coef[0]), .rdup_out(a9_wr[76]), .rdlo_out(a9_wr[78]));
			radix2 #(.width(width)) rd_st8_77  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[77]), .rdlo_in(a8_wr[79]),  .coef_in(coef[256]), .rdup_out(a9_wr[77]), .rdlo_out(a9_wr[79]));
			radix2 #(.width(width)) rd_st8_80  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[80]), .rdlo_in(a8_wr[82]),  .coef_in(coef[0]), .rdup_out(a9_wr[80]), .rdlo_out(a9_wr[82]));
			radix2 #(.width(width)) rd_st8_81  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[81]), .rdlo_in(a8_wr[83]),  .coef_in(coef[256]), .rdup_out(a9_wr[81]), .rdlo_out(a9_wr[83]));
			radix2 #(.width(width)) rd_st8_84  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[84]), .rdlo_in(a8_wr[86]),  .coef_in(coef[0]), .rdup_out(a9_wr[84]), .rdlo_out(a9_wr[86]));
			radix2 #(.width(width)) rd_st8_85  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[85]), .rdlo_in(a8_wr[87]),  .coef_in(coef[256]), .rdup_out(a9_wr[85]), .rdlo_out(a9_wr[87]));
			radix2 #(.width(width)) rd_st8_88  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[88]), .rdlo_in(a8_wr[90]),  .coef_in(coef[0]), .rdup_out(a9_wr[88]), .rdlo_out(a9_wr[90]));
			radix2 #(.width(width)) rd_st8_89  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[89]), .rdlo_in(a8_wr[91]),  .coef_in(coef[256]), .rdup_out(a9_wr[89]), .rdlo_out(a9_wr[91]));
			radix2 #(.width(width)) rd_st8_92  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[92]), .rdlo_in(a8_wr[94]),  .coef_in(coef[0]), .rdup_out(a9_wr[92]), .rdlo_out(a9_wr[94]));
			radix2 #(.width(width)) rd_st8_93  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[93]), .rdlo_in(a8_wr[95]),  .coef_in(coef[256]), .rdup_out(a9_wr[93]), .rdlo_out(a9_wr[95]));
			radix2 #(.width(width)) rd_st8_96  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[96]), .rdlo_in(a8_wr[98]),  .coef_in(coef[0]), .rdup_out(a9_wr[96]), .rdlo_out(a9_wr[98]));
			radix2 #(.width(width)) rd_st8_97  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[97]), .rdlo_in(a8_wr[99]),  .coef_in(coef[256]), .rdup_out(a9_wr[97]), .rdlo_out(a9_wr[99]));
			radix2 #(.width(width)) rd_st8_100  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[100]), .rdlo_in(a8_wr[102]),  .coef_in(coef[0]), .rdup_out(a9_wr[100]), .rdlo_out(a9_wr[102]));
			radix2 #(.width(width)) rd_st8_101  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[101]), .rdlo_in(a8_wr[103]),  .coef_in(coef[256]), .rdup_out(a9_wr[101]), .rdlo_out(a9_wr[103]));
			radix2 #(.width(width)) rd_st8_104  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[104]), .rdlo_in(a8_wr[106]),  .coef_in(coef[0]), .rdup_out(a9_wr[104]), .rdlo_out(a9_wr[106]));
			radix2 #(.width(width)) rd_st8_105  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[105]), .rdlo_in(a8_wr[107]),  .coef_in(coef[256]), .rdup_out(a9_wr[105]), .rdlo_out(a9_wr[107]));
			radix2 #(.width(width)) rd_st8_108  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[108]), .rdlo_in(a8_wr[110]),  .coef_in(coef[0]), .rdup_out(a9_wr[108]), .rdlo_out(a9_wr[110]));
			radix2 #(.width(width)) rd_st8_109  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[109]), .rdlo_in(a8_wr[111]),  .coef_in(coef[256]), .rdup_out(a9_wr[109]), .rdlo_out(a9_wr[111]));
			radix2 #(.width(width)) rd_st8_112  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[112]), .rdlo_in(a8_wr[114]),  .coef_in(coef[0]), .rdup_out(a9_wr[112]), .rdlo_out(a9_wr[114]));
			radix2 #(.width(width)) rd_st8_113  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[113]), .rdlo_in(a8_wr[115]),  .coef_in(coef[256]), .rdup_out(a9_wr[113]), .rdlo_out(a9_wr[115]));
			radix2 #(.width(width)) rd_st8_116  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[116]), .rdlo_in(a8_wr[118]),  .coef_in(coef[0]), .rdup_out(a9_wr[116]), .rdlo_out(a9_wr[118]));
			radix2 #(.width(width)) rd_st8_117  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[117]), .rdlo_in(a8_wr[119]),  .coef_in(coef[256]), .rdup_out(a9_wr[117]), .rdlo_out(a9_wr[119]));
			radix2 #(.width(width)) rd_st8_120  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[120]), .rdlo_in(a8_wr[122]),  .coef_in(coef[0]), .rdup_out(a9_wr[120]), .rdlo_out(a9_wr[122]));
			radix2 #(.width(width)) rd_st8_121  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[121]), .rdlo_in(a8_wr[123]),  .coef_in(coef[256]), .rdup_out(a9_wr[121]), .rdlo_out(a9_wr[123]));
			radix2 #(.width(width)) rd_st8_124  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[124]), .rdlo_in(a8_wr[126]),  .coef_in(coef[0]), .rdup_out(a9_wr[124]), .rdlo_out(a9_wr[126]));
			radix2 #(.width(width)) rd_st8_125  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[125]), .rdlo_in(a8_wr[127]),  .coef_in(coef[256]), .rdup_out(a9_wr[125]), .rdlo_out(a9_wr[127]));
			radix2 #(.width(width)) rd_st8_128  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[128]), .rdlo_in(a8_wr[130]),  .coef_in(coef[0]), .rdup_out(a9_wr[128]), .rdlo_out(a9_wr[130]));
			radix2 #(.width(width)) rd_st8_129  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[129]), .rdlo_in(a8_wr[131]),  .coef_in(coef[256]), .rdup_out(a9_wr[129]), .rdlo_out(a9_wr[131]));
			radix2 #(.width(width)) rd_st8_132  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[132]), .rdlo_in(a8_wr[134]),  .coef_in(coef[0]), .rdup_out(a9_wr[132]), .rdlo_out(a9_wr[134]));
			radix2 #(.width(width)) rd_st8_133  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[133]), .rdlo_in(a8_wr[135]),  .coef_in(coef[256]), .rdup_out(a9_wr[133]), .rdlo_out(a9_wr[135]));
			radix2 #(.width(width)) rd_st8_136  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[136]), .rdlo_in(a8_wr[138]),  .coef_in(coef[0]), .rdup_out(a9_wr[136]), .rdlo_out(a9_wr[138]));
			radix2 #(.width(width)) rd_st8_137  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[137]), .rdlo_in(a8_wr[139]),  .coef_in(coef[256]), .rdup_out(a9_wr[137]), .rdlo_out(a9_wr[139]));
			radix2 #(.width(width)) rd_st8_140  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[140]), .rdlo_in(a8_wr[142]),  .coef_in(coef[0]), .rdup_out(a9_wr[140]), .rdlo_out(a9_wr[142]));
			radix2 #(.width(width)) rd_st8_141  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[141]), .rdlo_in(a8_wr[143]),  .coef_in(coef[256]), .rdup_out(a9_wr[141]), .rdlo_out(a9_wr[143]));
			radix2 #(.width(width)) rd_st8_144  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[144]), .rdlo_in(a8_wr[146]),  .coef_in(coef[0]), .rdup_out(a9_wr[144]), .rdlo_out(a9_wr[146]));
			radix2 #(.width(width)) rd_st8_145  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[145]), .rdlo_in(a8_wr[147]),  .coef_in(coef[256]), .rdup_out(a9_wr[145]), .rdlo_out(a9_wr[147]));
			radix2 #(.width(width)) rd_st8_148  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[148]), .rdlo_in(a8_wr[150]),  .coef_in(coef[0]), .rdup_out(a9_wr[148]), .rdlo_out(a9_wr[150]));
			radix2 #(.width(width)) rd_st8_149  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[149]), .rdlo_in(a8_wr[151]),  .coef_in(coef[256]), .rdup_out(a9_wr[149]), .rdlo_out(a9_wr[151]));
			radix2 #(.width(width)) rd_st8_152  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[152]), .rdlo_in(a8_wr[154]),  .coef_in(coef[0]), .rdup_out(a9_wr[152]), .rdlo_out(a9_wr[154]));
			radix2 #(.width(width)) rd_st8_153  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[153]), .rdlo_in(a8_wr[155]),  .coef_in(coef[256]), .rdup_out(a9_wr[153]), .rdlo_out(a9_wr[155]));
			radix2 #(.width(width)) rd_st8_156  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[156]), .rdlo_in(a8_wr[158]),  .coef_in(coef[0]), .rdup_out(a9_wr[156]), .rdlo_out(a9_wr[158]));
			radix2 #(.width(width)) rd_st8_157  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[157]), .rdlo_in(a8_wr[159]),  .coef_in(coef[256]), .rdup_out(a9_wr[157]), .rdlo_out(a9_wr[159]));
			radix2 #(.width(width)) rd_st8_160  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[160]), .rdlo_in(a8_wr[162]),  .coef_in(coef[0]), .rdup_out(a9_wr[160]), .rdlo_out(a9_wr[162]));
			radix2 #(.width(width)) rd_st8_161  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[161]), .rdlo_in(a8_wr[163]),  .coef_in(coef[256]), .rdup_out(a9_wr[161]), .rdlo_out(a9_wr[163]));
			radix2 #(.width(width)) rd_st8_164  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[164]), .rdlo_in(a8_wr[166]),  .coef_in(coef[0]), .rdup_out(a9_wr[164]), .rdlo_out(a9_wr[166]));
			radix2 #(.width(width)) rd_st8_165  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[165]), .rdlo_in(a8_wr[167]),  .coef_in(coef[256]), .rdup_out(a9_wr[165]), .rdlo_out(a9_wr[167]));
			radix2 #(.width(width)) rd_st8_168  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[168]), .rdlo_in(a8_wr[170]),  .coef_in(coef[0]), .rdup_out(a9_wr[168]), .rdlo_out(a9_wr[170]));
			radix2 #(.width(width)) rd_st8_169  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[169]), .rdlo_in(a8_wr[171]),  .coef_in(coef[256]), .rdup_out(a9_wr[169]), .rdlo_out(a9_wr[171]));
			radix2 #(.width(width)) rd_st8_172  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[172]), .rdlo_in(a8_wr[174]),  .coef_in(coef[0]), .rdup_out(a9_wr[172]), .rdlo_out(a9_wr[174]));
			radix2 #(.width(width)) rd_st8_173  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[173]), .rdlo_in(a8_wr[175]),  .coef_in(coef[256]), .rdup_out(a9_wr[173]), .rdlo_out(a9_wr[175]));
			radix2 #(.width(width)) rd_st8_176  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[176]), .rdlo_in(a8_wr[178]),  .coef_in(coef[0]), .rdup_out(a9_wr[176]), .rdlo_out(a9_wr[178]));
			radix2 #(.width(width)) rd_st8_177  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[177]), .rdlo_in(a8_wr[179]),  .coef_in(coef[256]), .rdup_out(a9_wr[177]), .rdlo_out(a9_wr[179]));
			radix2 #(.width(width)) rd_st8_180  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[180]), .rdlo_in(a8_wr[182]),  .coef_in(coef[0]), .rdup_out(a9_wr[180]), .rdlo_out(a9_wr[182]));
			radix2 #(.width(width)) rd_st8_181  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[181]), .rdlo_in(a8_wr[183]),  .coef_in(coef[256]), .rdup_out(a9_wr[181]), .rdlo_out(a9_wr[183]));
			radix2 #(.width(width)) rd_st8_184  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[184]), .rdlo_in(a8_wr[186]),  .coef_in(coef[0]), .rdup_out(a9_wr[184]), .rdlo_out(a9_wr[186]));
			radix2 #(.width(width)) rd_st8_185  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[185]), .rdlo_in(a8_wr[187]),  .coef_in(coef[256]), .rdup_out(a9_wr[185]), .rdlo_out(a9_wr[187]));
			radix2 #(.width(width)) rd_st8_188  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[188]), .rdlo_in(a8_wr[190]),  .coef_in(coef[0]), .rdup_out(a9_wr[188]), .rdlo_out(a9_wr[190]));
			radix2 #(.width(width)) rd_st8_189  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[189]), .rdlo_in(a8_wr[191]),  .coef_in(coef[256]), .rdup_out(a9_wr[189]), .rdlo_out(a9_wr[191]));
			radix2 #(.width(width)) rd_st8_192  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[192]), .rdlo_in(a8_wr[194]),  .coef_in(coef[0]), .rdup_out(a9_wr[192]), .rdlo_out(a9_wr[194]));
			radix2 #(.width(width)) rd_st8_193  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[193]), .rdlo_in(a8_wr[195]),  .coef_in(coef[256]), .rdup_out(a9_wr[193]), .rdlo_out(a9_wr[195]));
			radix2 #(.width(width)) rd_st8_196  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[196]), .rdlo_in(a8_wr[198]),  .coef_in(coef[0]), .rdup_out(a9_wr[196]), .rdlo_out(a9_wr[198]));
			radix2 #(.width(width)) rd_st8_197  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[197]), .rdlo_in(a8_wr[199]),  .coef_in(coef[256]), .rdup_out(a9_wr[197]), .rdlo_out(a9_wr[199]));
			radix2 #(.width(width)) rd_st8_200  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[200]), .rdlo_in(a8_wr[202]),  .coef_in(coef[0]), .rdup_out(a9_wr[200]), .rdlo_out(a9_wr[202]));
			radix2 #(.width(width)) rd_st8_201  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[201]), .rdlo_in(a8_wr[203]),  .coef_in(coef[256]), .rdup_out(a9_wr[201]), .rdlo_out(a9_wr[203]));
			radix2 #(.width(width)) rd_st8_204  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[204]), .rdlo_in(a8_wr[206]),  .coef_in(coef[0]), .rdup_out(a9_wr[204]), .rdlo_out(a9_wr[206]));
			radix2 #(.width(width)) rd_st8_205  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[205]), .rdlo_in(a8_wr[207]),  .coef_in(coef[256]), .rdup_out(a9_wr[205]), .rdlo_out(a9_wr[207]));
			radix2 #(.width(width)) rd_st8_208  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[208]), .rdlo_in(a8_wr[210]),  .coef_in(coef[0]), .rdup_out(a9_wr[208]), .rdlo_out(a9_wr[210]));
			radix2 #(.width(width)) rd_st8_209  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[209]), .rdlo_in(a8_wr[211]),  .coef_in(coef[256]), .rdup_out(a9_wr[209]), .rdlo_out(a9_wr[211]));
			radix2 #(.width(width)) rd_st8_212  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[212]), .rdlo_in(a8_wr[214]),  .coef_in(coef[0]), .rdup_out(a9_wr[212]), .rdlo_out(a9_wr[214]));
			radix2 #(.width(width)) rd_st8_213  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[213]), .rdlo_in(a8_wr[215]),  .coef_in(coef[256]), .rdup_out(a9_wr[213]), .rdlo_out(a9_wr[215]));
			radix2 #(.width(width)) rd_st8_216  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[216]), .rdlo_in(a8_wr[218]),  .coef_in(coef[0]), .rdup_out(a9_wr[216]), .rdlo_out(a9_wr[218]));
			radix2 #(.width(width)) rd_st8_217  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[217]), .rdlo_in(a8_wr[219]),  .coef_in(coef[256]), .rdup_out(a9_wr[217]), .rdlo_out(a9_wr[219]));
			radix2 #(.width(width)) rd_st8_220  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[220]), .rdlo_in(a8_wr[222]),  .coef_in(coef[0]), .rdup_out(a9_wr[220]), .rdlo_out(a9_wr[222]));
			radix2 #(.width(width)) rd_st8_221  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[221]), .rdlo_in(a8_wr[223]),  .coef_in(coef[256]), .rdup_out(a9_wr[221]), .rdlo_out(a9_wr[223]));
			radix2 #(.width(width)) rd_st8_224  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[224]), .rdlo_in(a8_wr[226]),  .coef_in(coef[0]), .rdup_out(a9_wr[224]), .rdlo_out(a9_wr[226]));
			radix2 #(.width(width)) rd_st8_225  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[225]), .rdlo_in(a8_wr[227]),  .coef_in(coef[256]), .rdup_out(a9_wr[225]), .rdlo_out(a9_wr[227]));
			radix2 #(.width(width)) rd_st8_228  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[228]), .rdlo_in(a8_wr[230]),  .coef_in(coef[0]), .rdup_out(a9_wr[228]), .rdlo_out(a9_wr[230]));
			radix2 #(.width(width)) rd_st8_229  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[229]), .rdlo_in(a8_wr[231]),  .coef_in(coef[256]), .rdup_out(a9_wr[229]), .rdlo_out(a9_wr[231]));
			radix2 #(.width(width)) rd_st8_232  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[232]), .rdlo_in(a8_wr[234]),  .coef_in(coef[0]), .rdup_out(a9_wr[232]), .rdlo_out(a9_wr[234]));
			radix2 #(.width(width)) rd_st8_233  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[233]), .rdlo_in(a8_wr[235]),  .coef_in(coef[256]), .rdup_out(a9_wr[233]), .rdlo_out(a9_wr[235]));
			radix2 #(.width(width)) rd_st8_236  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[236]), .rdlo_in(a8_wr[238]),  .coef_in(coef[0]), .rdup_out(a9_wr[236]), .rdlo_out(a9_wr[238]));
			radix2 #(.width(width)) rd_st8_237  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[237]), .rdlo_in(a8_wr[239]),  .coef_in(coef[256]), .rdup_out(a9_wr[237]), .rdlo_out(a9_wr[239]));
			radix2 #(.width(width)) rd_st8_240  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[240]), .rdlo_in(a8_wr[242]),  .coef_in(coef[0]), .rdup_out(a9_wr[240]), .rdlo_out(a9_wr[242]));
			radix2 #(.width(width)) rd_st8_241  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[241]), .rdlo_in(a8_wr[243]),  .coef_in(coef[256]), .rdup_out(a9_wr[241]), .rdlo_out(a9_wr[243]));
			radix2 #(.width(width)) rd_st8_244  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[244]), .rdlo_in(a8_wr[246]),  .coef_in(coef[0]), .rdup_out(a9_wr[244]), .rdlo_out(a9_wr[246]));
			radix2 #(.width(width)) rd_st8_245  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[245]), .rdlo_in(a8_wr[247]),  .coef_in(coef[256]), .rdup_out(a9_wr[245]), .rdlo_out(a9_wr[247]));
			radix2 #(.width(width)) rd_st8_248  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[248]), .rdlo_in(a8_wr[250]),  .coef_in(coef[0]), .rdup_out(a9_wr[248]), .rdlo_out(a9_wr[250]));
			radix2 #(.width(width)) rd_st8_249  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[249]), .rdlo_in(a8_wr[251]),  .coef_in(coef[256]), .rdup_out(a9_wr[249]), .rdlo_out(a9_wr[251]));
			radix2 #(.width(width)) rd_st8_252  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[252]), .rdlo_in(a8_wr[254]),  .coef_in(coef[0]), .rdup_out(a9_wr[252]), .rdlo_out(a9_wr[254]));
			radix2 #(.width(width)) rd_st8_253  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[253]), .rdlo_in(a8_wr[255]),  .coef_in(coef[256]), .rdup_out(a9_wr[253]), .rdlo_out(a9_wr[255]));
			radix2 #(.width(width)) rd_st8_256  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[256]), .rdlo_in(a8_wr[258]),  .coef_in(coef[0]), .rdup_out(a9_wr[256]), .rdlo_out(a9_wr[258]));
			radix2 #(.width(width)) rd_st8_257  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[257]), .rdlo_in(a8_wr[259]),  .coef_in(coef[256]), .rdup_out(a9_wr[257]), .rdlo_out(a9_wr[259]));
			radix2 #(.width(width)) rd_st8_260  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[260]), .rdlo_in(a8_wr[262]),  .coef_in(coef[0]), .rdup_out(a9_wr[260]), .rdlo_out(a9_wr[262]));
			radix2 #(.width(width)) rd_st8_261  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[261]), .rdlo_in(a8_wr[263]),  .coef_in(coef[256]), .rdup_out(a9_wr[261]), .rdlo_out(a9_wr[263]));
			radix2 #(.width(width)) rd_st8_264  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[264]), .rdlo_in(a8_wr[266]),  .coef_in(coef[0]), .rdup_out(a9_wr[264]), .rdlo_out(a9_wr[266]));
			radix2 #(.width(width)) rd_st8_265  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[265]), .rdlo_in(a8_wr[267]),  .coef_in(coef[256]), .rdup_out(a9_wr[265]), .rdlo_out(a9_wr[267]));
			radix2 #(.width(width)) rd_st8_268  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[268]), .rdlo_in(a8_wr[270]),  .coef_in(coef[0]), .rdup_out(a9_wr[268]), .rdlo_out(a9_wr[270]));
			radix2 #(.width(width)) rd_st8_269  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[269]), .rdlo_in(a8_wr[271]),  .coef_in(coef[256]), .rdup_out(a9_wr[269]), .rdlo_out(a9_wr[271]));
			radix2 #(.width(width)) rd_st8_272  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[272]), .rdlo_in(a8_wr[274]),  .coef_in(coef[0]), .rdup_out(a9_wr[272]), .rdlo_out(a9_wr[274]));
			radix2 #(.width(width)) rd_st8_273  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[273]), .rdlo_in(a8_wr[275]),  .coef_in(coef[256]), .rdup_out(a9_wr[273]), .rdlo_out(a9_wr[275]));
			radix2 #(.width(width)) rd_st8_276  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[276]), .rdlo_in(a8_wr[278]),  .coef_in(coef[0]), .rdup_out(a9_wr[276]), .rdlo_out(a9_wr[278]));
			radix2 #(.width(width)) rd_st8_277  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[277]), .rdlo_in(a8_wr[279]),  .coef_in(coef[256]), .rdup_out(a9_wr[277]), .rdlo_out(a9_wr[279]));
			radix2 #(.width(width)) rd_st8_280  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[280]), .rdlo_in(a8_wr[282]),  .coef_in(coef[0]), .rdup_out(a9_wr[280]), .rdlo_out(a9_wr[282]));
			radix2 #(.width(width)) rd_st8_281  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[281]), .rdlo_in(a8_wr[283]),  .coef_in(coef[256]), .rdup_out(a9_wr[281]), .rdlo_out(a9_wr[283]));
			radix2 #(.width(width)) rd_st8_284  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[284]), .rdlo_in(a8_wr[286]),  .coef_in(coef[0]), .rdup_out(a9_wr[284]), .rdlo_out(a9_wr[286]));
			radix2 #(.width(width)) rd_st8_285  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[285]), .rdlo_in(a8_wr[287]),  .coef_in(coef[256]), .rdup_out(a9_wr[285]), .rdlo_out(a9_wr[287]));
			radix2 #(.width(width)) rd_st8_288  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[288]), .rdlo_in(a8_wr[290]),  .coef_in(coef[0]), .rdup_out(a9_wr[288]), .rdlo_out(a9_wr[290]));
			radix2 #(.width(width)) rd_st8_289  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[289]), .rdlo_in(a8_wr[291]),  .coef_in(coef[256]), .rdup_out(a9_wr[289]), .rdlo_out(a9_wr[291]));
			radix2 #(.width(width)) rd_st8_292  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[292]), .rdlo_in(a8_wr[294]),  .coef_in(coef[0]), .rdup_out(a9_wr[292]), .rdlo_out(a9_wr[294]));
			radix2 #(.width(width)) rd_st8_293  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[293]), .rdlo_in(a8_wr[295]),  .coef_in(coef[256]), .rdup_out(a9_wr[293]), .rdlo_out(a9_wr[295]));
			radix2 #(.width(width)) rd_st8_296  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[296]), .rdlo_in(a8_wr[298]),  .coef_in(coef[0]), .rdup_out(a9_wr[296]), .rdlo_out(a9_wr[298]));
			radix2 #(.width(width)) rd_st8_297  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[297]), .rdlo_in(a8_wr[299]),  .coef_in(coef[256]), .rdup_out(a9_wr[297]), .rdlo_out(a9_wr[299]));
			radix2 #(.width(width)) rd_st8_300  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[300]), .rdlo_in(a8_wr[302]),  .coef_in(coef[0]), .rdup_out(a9_wr[300]), .rdlo_out(a9_wr[302]));
			radix2 #(.width(width)) rd_st8_301  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[301]), .rdlo_in(a8_wr[303]),  .coef_in(coef[256]), .rdup_out(a9_wr[301]), .rdlo_out(a9_wr[303]));
			radix2 #(.width(width)) rd_st8_304  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[304]), .rdlo_in(a8_wr[306]),  .coef_in(coef[0]), .rdup_out(a9_wr[304]), .rdlo_out(a9_wr[306]));
			radix2 #(.width(width)) rd_st8_305  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[305]), .rdlo_in(a8_wr[307]),  .coef_in(coef[256]), .rdup_out(a9_wr[305]), .rdlo_out(a9_wr[307]));
			radix2 #(.width(width)) rd_st8_308  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[308]), .rdlo_in(a8_wr[310]),  .coef_in(coef[0]), .rdup_out(a9_wr[308]), .rdlo_out(a9_wr[310]));
			radix2 #(.width(width)) rd_st8_309  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[309]), .rdlo_in(a8_wr[311]),  .coef_in(coef[256]), .rdup_out(a9_wr[309]), .rdlo_out(a9_wr[311]));
			radix2 #(.width(width)) rd_st8_312  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[312]), .rdlo_in(a8_wr[314]),  .coef_in(coef[0]), .rdup_out(a9_wr[312]), .rdlo_out(a9_wr[314]));
			radix2 #(.width(width)) rd_st8_313  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[313]), .rdlo_in(a8_wr[315]),  .coef_in(coef[256]), .rdup_out(a9_wr[313]), .rdlo_out(a9_wr[315]));
			radix2 #(.width(width)) rd_st8_316  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[316]), .rdlo_in(a8_wr[318]),  .coef_in(coef[0]), .rdup_out(a9_wr[316]), .rdlo_out(a9_wr[318]));
			radix2 #(.width(width)) rd_st8_317  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[317]), .rdlo_in(a8_wr[319]),  .coef_in(coef[256]), .rdup_out(a9_wr[317]), .rdlo_out(a9_wr[319]));
			radix2 #(.width(width)) rd_st8_320  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[320]), .rdlo_in(a8_wr[322]),  .coef_in(coef[0]), .rdup_out(a9_wr[320]), .rdlo_out(a9_wr[322]));
			radix2 #(.width(width)) rd_st8_321  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[321]), .rdlo_in(a8_wr[323]),  .coef_in(coef[256]), .rdup_out(a9_wr[321]), .rdlo_out(a9_wr[323]));
			radix2 #(.width(width)) rd_st8_324  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[324]), .rdlo_in(a8_wr[326]),  .coef_in(coef[0]), .rdup_out(a9_wr[324]), .rdlo_out(a9_wr[326]));
			radix2 #(.width(width)) rd_st8_325  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[325]), .rdlo_in(a8_wr[327]),  .coef_in(coef[256]), .rdup_out(a9_wr[325]), .rdlo_out(a9_wr[327]));
			radix2 #(.width(width)) rd_st8_328  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[328]), .rdlo_in(a8_wr[330]),  .coef_in(coef[0]), .rdup_out(a9_wr[328]), .rdlo_out(a9_wr[330]));
			radix2 #(.width(width)) rd_st8_329  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[329]), .rdlo_in(a8_wr[331]),  .coef_in(coef[256]), .rdup_out(a9_wr[329]), .rdlo_out(a9_wr[331]));
			radix2 #(.width(width)) rd_st8_332  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[332]), .rdlo_in(a8_wr[334]),  .coef_in(coef[0]), .rdup_out(a9_wr[332]), .rdlo_out(a9_wr[334]));
			radix2 #(.width(width)) rd_st8_333  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[333]), .rdlo_in(a8_wr[335]),  .coef_in(coef[256]), .rdup_out(a9_wr[333]), .rdlo_out(a9_wr[335]));
			radix2 #(.width(width)) rd_st8_336  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[336]), .rdlo_in(a8_wr[338]),  .coef_in(coef[0]), .rdup_out(a9_wr[336]), .rdlo_out(a9_wr[338]));
			radix2 #(.width(width)) rd_st8_337  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[337]), .rdlo_in(a8_wr[339]),  .coef_in(coef[256]), .rdup_out(a9_wr[337]), .rdlo_out(a9_wr[339]));
			radix2 #(.width(width)) rd_st8_340  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[340]), .rdlo_in(a8_wr[342]),  .coef_in(coef[0]), .rdup_out(a9_wr[340]), .rdlo_out(a9_wr[342]));
			radix2 #(.width(width)) rd_st8_341  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[341]), .rdlo_in(a8_wr[343]),  .coef_in(coef[256]), .rdup_out(a9_wr[341]), .rdlo_out(a9_wr[343]));
			radix2 #(.width(width)) rd_st8_344  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[344]), .rdlo_in(a8_wr[346]),  .coef_in(coef[0]), .rdup_out(a9_wr[344]), .rdlo_out(a9_wr[346]));
			radix2 #(.width(width)) rd_st8_345  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[345]), .rdlo_in(a8_wr[347]),  .coef_in(coef[256]), .rdup_out(a9_wr[345]), .rdlo_out(a9_wr[347]));
			radix2 #(.width(width)) rd_st8_348  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[348]), .rdlo_in(a8_wr[350]),  .coef_in(coef[0]), .rdup_out(a9_wr[348]), .rdlo_out(a9_wr[350]));
			radix2 #(.width(width)) rd_st8_349  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[349]), .rdlo_in(a8_wr[351]),  .coef_in(coef[256]), .rdup_out(a9_wr[349]), .rdlo_out(a9_wr[351]));
			radix2 #(.width(width)) rd_st8_352  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[352]), .rdlo_in(a8_wr[354]),  .coef_in(coef[0]), .rdup_out(a9_wr[352]), .rdlo_out(a9_wr[354]));
			radix2 #(.width(width)) rd_st8_353  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[353]), .rdlo_in(a8_wr[355]),  .coef_in(coef[256]), .rdup_out(a9_wr[353]), .rdlo_out(a9_wr[355]));
			radix2 #(.width(width)) rd_st8_356  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[356]), .rdlo_in(a8_wr[358]),  .coef_in(coef[0]), .rdup_out(a9_wr[356]), .rdlo_out(a9_wr[358]));
			radix2 #(.width(width)) rd_st8_357  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[357]), .rdlo_in(a8_wr[359]),  .coef_in(coef[256]), .rdup_out(a9_wr[357]), .rdlo_out(a9_wr[359]));
			radix2 #(.width(width)) rd_st8_360  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[360]), .rdlo_in(a8_wr[362]),  .coef_in(coef[0]), .rdup_out(a9_wr[360]), .rdlo_out(a9_wr[362]));
			radix2 #(.width(width)) rd_st8_361  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[361]), .rdlo_in(a8_wr[363]),  .coef_in(coef[256]), .rdup_out(a9_wr[361]), .rdlo_out(a9_wr[363]));
			radix2 #(.width(width)) rd_st8_364  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[364]), .rdlo_in(a8_wr[366]),  .coef_in(coef[0]), .rdup_out(a9_wr[364]), .rdlo_out(a9_wr[366]));
			radix2 #(.width(width)) rd_st8_365  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[365]), .rdlo_in(a8_wr[367]),  .coef_in(coef[256]), .rdup_out(a9_wr[365]), .rdlo_out(a9_wr[367]));
			radix2 #(.width(width)) rd_st8_368  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[368]), .rdlo_in(a8_wr[370]),  .coef_in(coef[0]), .rdup_out(a9_wr[368]), .rdlo_out(a9_wr[370]));
			radix2 #(.width(width)) rd_st8_369  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[369]), .rdlo_in(a8_wr[371]),  .coef_in(coef[256]), .rdup_out(a9_wr[369]), .rdlo_out(a9_wr[371]));
			radix2 #(.width(width)) rd_st8_372  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[372]), .rdlo_in(a8_wr[374]),  .coef_in(coef[0]), .rdup_out(a9_wr[372]), .rdlo_out(a9_wr[374]));
			radix2 #(.width(width)) rd_st8_373  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[373]), .rdlo_in(a8_wr[375]),  .coef_in(coef[256]), .rdup_out(a9_wr[373]), .rdlo_out(a9_wr[375]));
			radix2 #(.width(width)) rd_st8_376  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[376]), .rdlo_in(a8_wr[378]),  .coef_in(coef[0]), .rdup_out(a9_wr[376]), .rdlo_out(a9_wr[378]));
			radix2 #(.width(width)) rd_st8_377  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[377]), .rdlo_in(a8_wr[379]),  .coef_in(coef[256]), .rdup_out(a9_wr[377]), .rdlo_out(a9_wr[379]));
			radix2 #(.width(width)) rd_st8_380  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[380]), .rdlo_in(a8_wr[382]),  .coef_in(coef[0]), .rdup_out(a9_wr[380]), .rdlo_out(a9_wr[382]));
			radix2 #(.width(width)) rd_st8_381  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[381]), .rdlo_in(a8_wr[383]),  .coef_in(coef[256]), .rdup_out(a9_wr[381]), .rdlo_out(a9_wr[383]));
			radix2 #(.width(width)) rd_st8_384  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[384]), .rdlo_in(a8_wr[386]),  .coef_in(coef[0]), .rdup_out(a9_wr[384]), .rdlo_out(a9_wr[386]));
			radix2 #(.width(width)) rd_st8_385  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[385]), .rdlo_in(a8_wr[387]),  .coef_in(coef[256]), .rdup_out(a9_wr[385]), .rdlo_out(a9_wr[387]));
			radix2 #(.width(width)) rd_st8_388  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[388]), .rdlo_in(a8_wr[390]),  .coef_in(coef[0]), .rdup_out(a9_wr[388]), .rdlo_out(a9_wr[390]));
			radix2 #(.width(width)) rd_st8_389  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[389]), .rdlo_in(a8_wr[391]),  .coef_in(coef[256]), .rdup_out(a9_wr[389]), .rdlo_out(a9_wr[391]));
			radix2 #(.width(width)) rd_st8_392  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[392]), .rdlo_in(a8_wr[394]),  .coef_in(coef[0]), .rdup_out(a9_wr[392]), .rdlo_out(a9_wr[394]));
			radix2 #(.width(width)) rd_st8_393  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[393]), .rdlo_in(a8_wr[395]),  .coef_in(coef[256]), .rdup_out(a9_wr[393]), .rdlo_out(a9_wr[395]));
			radix2 #(.width(width)) rd_st8_396  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[396]), .rdlo_in(a8_wr[398]),  .coef_in(coef[0]), .rdup_out(a9_wr[396]), .rdlo_out(a9_wr[398]));
			radix2 #(.width(width)) rd_st8_397  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[397]), .rdlo_in(a8_wr[399]),  .coef_in(coef[256]), .rdup_out(a9_wr[397]), .rdlo_out(a9_wr[399]));
			radix2 #(.width(width)) rd_st8_400  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[400]), .rdlo_in(a8_wr[402]),  .coef_in(coef[0]), .rdup_out(a9_wr[400]), .rdlo_out(a9_wr[402]));
			radix2 #(.width(width)) rd_st8_401  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[401]), .rdlo_in(a8_wr[403]),  .coef_in(coef[256]), .rdup_out(a9_wr[401]), .rdlo_out(a9_wr[403]));
			radix2 #(.width(width)) rd_st8_404  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[404]), .rdlo_in(a8_wr[406]),  .coef_in(coef[0]), .rdup_out(a9_wr[404]), .rdlo_out(a9_wr[406]));
			radix2 #(.width(width)) rd_st8_405  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[405]), .rdlo_in(a8_wr[407]),  .coef_in(coef[256]), .rdup_out(a9_wr[405]), .rdlo_out(a9_wr[407]));
			radix2 #(.width(width)) rd_st8_408  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[408]), .rdlo_in(a8_wr[410]),  .coef_in(coef[0]), .rdup_out(a9_wr[408]), .rdlo_out(a9_wr[410]));
			radix2 #(.width(width)) rd_st8_409  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[409]), .rdlo_in(a8_wr[411]),  .coef_in(coef[256]), .rdup_out(a9_wr[409]), .rdlo_out(a9_wr[411]));
			radix2 #(.width(width)) rd_st8_412  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[412]), .rdlo_in(a8_wr[414]),  .coef_in(coef[0]), .rdup_out(a9_wr[412]), .rdlo_out(a9_wr[414]));
			radix2 #(.width(width)) rd_st8_413  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[413]), .rdlo_in(a8_wr[415]),  .coef_in(coef[256]), .rdup_out(a9_wr[413]), .rdlo_out(a9_wr[415]));
			radix2 #(.width(width)) rd_st8_416  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[416]), .rdlo_in(a8_wr[418]),  .coef_in(coef[0]), .rdup_out(a9_wr[416]), .rdlo_out(a9_wr[418]));
			radix2 #(.width(width)) rd_st8_417  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[417]), .rdlo_in(a8_wr[419]),  .coef_in(coef[256]), .rdup_out(a9_wr[417]), .rdlo_out(a9_wr[419]));
			radix2 #(.width(width)) rd_st8_420  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[420]), .rdlo_in(a8_wr[422]),  .coef_in(coef[0]), .rdup_out(a9_wr[420]), .rdlo_out(a9_wr[422]));
			radix2 #(.width(width)) rd_st8_421  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[421]), .rdlo_in(a8_wr[423]),  .coef_in(coef[256]), .rdup_out(a9_wr[421]), .rdlo_out(a9_wr[423]));
			radix2 #(.width(width)) rd_st8_424  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[424]), .rdlo_in(a8_wr[426]),  .coef_in(coef[0]), .rdup_out(a9_wr[424]), .rdlo_out(a9_wr[426]));
			radix2 #(.width(width)) rd_st8_425  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[425]), .rdlo_in(a8_wr[427]),  .coef_in(coef[256]), .rdup_out(a9_wr[425]), .rdlo_out(a9_wr[427]));
			radix2 #(.width(width)) rd_st8_428  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[428]), .rdlo_in(a8_wr[430]),  .coef_in(coef[0]), .rdup_out(a9_wr[428]), .rdlo_out(a9_wr[430]));
			radix2 #(.width(width)) rd_st8_429  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[429]), .rdlo_in(a8_wr[431]),  .coef_in(coef[256]), .rdup_out(a9_wr[429]), .rdlo_out(a9_wr[431]));
			radix2 #(.width(width)) rd_st8_432  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[432]), .rdlo_in(a8_wr[434]),  .coef_in(coef[0]), .rdup_out(a9_wr[432]), .rdlo_out(a9_wr[434]));
			radix2 #(.width(width)) rd_st8_433  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[433]), .rdlo_in(a8_wr[435]),  .coef_in(coef[256]), .rdup_out(a9_wr[433]), .rdlo_out(a9_wr[435]));
			radix2 #(.width(width)) rd_st8_436  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[436]), .rdlo_in(a8_wr[438]),  .coef_in(coef[0]), .rdup_out(a9_wr[436]), .rdlo_out(a9_wr[438]));
			radix2 #(.width(width)) rd_st8_437  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[437]), .rdlo_in(a8_wr[439]),  .coef_in(coef[256]), .rdup_out(a9_wr[437]), .rdlo_out(a9_wr[439]));
			radix2 #(.width(width)) rd_st8_440  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[440]), .rdlo_in(a8_wr[442]),  .coef_in(coef[0]), .rdup_out(a9_wr[440]), .rdlo_out(a9_wr[442]));
			radix2 #(.width(width)) rd_st8_441  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[441]), .rdlo_in(a8_wr[443]),  .coef_in(coef[256]), .rdup_out(a9_wr[441]), .rdlo_out(a9_wr[443]));
			radix2 #(.width(width)) rd_st8_444  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[444]), .rdlo_in(a8_wr[446]),  .coef_in(coef[0]), .rdup_out(a9_wr[444]), .rdlo_out(a9_wr[446]));
			radix2 #(.width(width)) rd_st8_445  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[445]), .rdlo_in(a8_wr[447]),  .coef_in(coef[256]), .rdup_out(a9_wr[445]), .rdlo_out(a9_wr[447]));
			radix2 #(.width(width)) rd_st8_448  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[448]), .rdlo_in(a8_wr[450]),  .coef_in(coef[0]), .rdup_out(a9_wr[448]), .rdlo_out(a9_wr[450]));
			radix2 #(.width(width)) rd_st8_449  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[449]), .rdlo_in(a8_wr[451]),  .coef_in(coef[256]), .rdup_out(a9_wr[449]), .rdlo_out(a9_wr[451]));
			radix2 #(.width(width)) rd_st8_452  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[452]), .rdlo_in(a8_wr[454]),  .coef_in(coef[0]), .rdup_out(a9_wr[452]), .rdlo_out(a9_wr[454]));
			radix2 #(.width(width)) rd_st8_453  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[453]), .rdlo_in(a8_wr[455]),  .coef_in(coef[256]), .rdup_out(a9_wr[453]), .rdlo_out(a9_wr[455]));
			radix2 #(.width(width)) rd_st8_456  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[456]), .rdlo_in(a8_wr[458]),  .coef_in(coef[0]), .rdup_out(a9_wr[456]), .rdlo_out(a9_wr[458]));
			radix2 #(.width(width)) rd_st8_457  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[457]), .rdlo_in(a8_wr[459]),  .coef_in(coef[256]), .rdup_out(a9_wr[457]), .rdlo_out(a9_wr[459]));
			radix2 #(.width(width)) rd_st8_460  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[460]), .rdlo_in(a8_wr[462]),  .coef_in(coef[0]), .rdup_out(a9_wr[460]), .rdlo_out(a9_wr[462]));
			radix2 #(.width(width)) rd_st8_461  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[461]), .rdlo_in(a8_wr[463]),  .coef_in(coef[256]), .rdup_out(a9_wr[461]), .rdlo_out(a9_wr[463]));
			radix2 #(.width(width)) rd_st8_464  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[464]), .rdlo_in(a8_wr[466]),  .coef_in(coef[0]), .rdup_out(a9_wr[464]), .rdlo_out(a9_wr[466]));
			radix2 #(.width(width)) rd_st8_465  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[465]), .rdlo_in(a8_wr[467]),  .coef_in(coef[256]), .rdup_out(a9_wr[465]), .rdlo_out(a9_wr[467]));
			radix2 #(.width(width)) rd_st8_468  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[468]), .rdlo_in(a8_wr[470]),  .coef_in(coef[0]), .rdup_out(a9_wr[468]), .rdlo_out(a9_wr[470]));
			radix2 #(.width(width)) rd_st8_469  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[469]), .rdlo_in(a8_wr[471]),  .coef_in(coef[256]), .rdup_out(a9_wr[469]), .rdlo_out(a9_wr[471]));
			radix2 #(.width(width)) rd_st8_472  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[472]), .rdlo_in(a8_wr[474]),  .coef_in(coef[0]), .rdup_out(a9_wr[472]), .rdlo_out(a9_wr[474]));
			radix2 #(.width(width)) rd_st8_473  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[473]), .rdlo_in(a8_wr[475]),  .coef_in(coef[256]), .rdup_out(a9_wr[473]), .rdlo_out(a9_wr[475]));
			radix2 #(.width(width)) rd_st8_476  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[476]), .rdlo_in(a8_wr[478]),  .coef_in(coef[0]), .rdup_out(a9_wr[476]), .rdlo_out(a9_wr[478]));
			radix2 #(.width(width)) rd_st8_477  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[477]), .rdlo_in(a8_wr[479]),  .coef_in(coef[256]), .rdup_out(a9_wr[477]), .rdlo_out(a9_wr[479]));
			radix2 #(.width(width)) rd_st8_480  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[480]), .rdlo_in(a8_wr[482]),  .coef_in(coef[0]), .rdup_out(a9_wr[480]), .rdlo_out(a9_wr[482]));
			radix2 #(.width(width)) rd_st8_481  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[481]), .rdlo_in(a8_wr[483]),  .coef_in(coef[256]), .rdup_out(a9_wr[481]), .rdlo_out(a9_wr[483]));
			radix2 #(.width(width)) rd_st8_484  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[484]), .rdlo_in(a8_wr[486]),  .coef_in(coef[0]), .rdup_out(a9_wr[484]), .rdlo_out(a9_wr[486]));
			radix2 #(.width(width)) rd_st8_485  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[485]), .rdlo_in(a8_wr[487]),  .coef_in(coef[256]), .rdup_out(a9_wr[485]), .rdlo_out(a9_wr[487]));
			radix2 #(.width(width)) rd_st8_488  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[488]), .rdlo_in(a8_wr[490]),  .coef_in(coef[0]), .rdup_out(a9_wr[488]), .rdlo_out(a9_wr[490]));
			radix2 #(.width(width)) rd_st8_489  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[489]), .rdlo_in(a8_wr[491]),  .coef_in(coef[256]), .rdup_out(a9_wr[489]), .rdlo_out(a9_wr[491]));
			radix2 #(.width(width)) rd_st8_492  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[492]), .rdlo_in(a8_wr[494]),  .coef_in(coef[0]), .rdup_out(a9_wr[492]), .rdlo_out(a9_wr[494]));
			radix2 #(.width(width)) rd_st8_493  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[493]), .rdlo_in(a8_wr[495]),  .coef_in(coef[256]), .rdup_out(a9_wr[493]), .rdlo_out(a9_wr[495]));
			radix2 #(.width(width)) rd_st8_496  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[496]), .rdlo_in(a8_wr[498]),  .coef_in(coef[0]), .rdup_out(a9_wr[496]), .rdlo_out(a9_wr[498]));
			radix2 #(.width(width)) rd_st8_497  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[497]), .rdlo_in(a8_wr[499]),  .coef_in(coef[256]), .rdup_out(a9_wr[497]), .rdlo_out(a9_wr[499]));
			radix2 #(.width(width)) rd_st8_500  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[500]), .rdlo_in(a8_wr[502]),  .coef_in(coef[0]), .rdup_out(a9_wr[500]), .rdlo_out(a9_wr[502]));
			radix2 #(.width(width)) rd_st8_501  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[501]), .rdlo_in(a8_wr[503]),  .coef_in(coef[256]), .rdup_out(a9_wr[501]), .rdlo_out(a9_wr[503]));
			radix2 #(.width(width)) rd_st8_504  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[504]), .rdlo_in(a8_wr[506]),  .coef_in(coef[0]), .rdup_out(a9_wr[504]), .rdlo_out(a9_wr[506]));
			radix2 #(.width(width)) rd_st8_505  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[505]), .rdlo_in(a8_wr[507]),  .coef_in(coef[256]), .rdup_out(a9_wr[505]), .rdlo_out(a9_wr[507]));
			radix2 #(.width(width)) rd_st8_508  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[508]), .rdlo_in(a8_wr[510]),  .coef_in(coef[0]), .rdup_out(a9_wr[508]), .rdlo_out(a9_wr[510]));
			radix2 #(.width(width)) rd_st8_509  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[509]), .rdlo_in(a8_wr[511]),  .coef_in(coef[256]), .rdup_out(a9_wr[509]), .rdlo_out(a9_wr[511]));
			radix2 #(.width(width)) rd_st8_512  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[512]), .rdlo_in(a8_wr[514]),  .coef_in(coef[0]), .rdup_out(a9_wr[512]), .rdlo_out(a9_wr[514]));
			radix2 #(.width(width)) rd_st8_513  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[513]), .rdlo_in(a8_wr[515]),  .coef_in(coef[256]), .rdup_out(a9_wr[513]), .rdlo_out(a9_wr[515]));
			radix2 #(.width(width)) rd_st8_516  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[516]), .rdlo_in(a8_wr[518]),  .coef_in(coef[0]), .rdup_out(a9_wr[516]), .rdlo_out(a9_wr[518]));
			radix2 #(.width(width)) rd_st8_517  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[517]), .rdlo_in(a8_wr[519]),  .coef_in(coef[256]), .rdup_out(a9_wr[517]), .rdlo_out(a9_wr[519]));
			radix2 #(.width(width)) rd_st8_520  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[520]), .rdlo_in(a8_wr[522]),  .coef_in(coef[0]), .rdup_out(a9_wr[520]), .rdlo_out(a9_wr[522]));
			radix2 #(.width(width)) rd_st8_521  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[521]), .rdlo_in(a8_wr[523]),  .coef_in(coef[256]), .rdup_out(a9_wr[521]), .rdlo_out(a9_wr[523]));
			radix2 #(.width(width)) rd_st8_524  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[524]), .rdlo_in(a8_wr[526]),  .coef_in(coef[0]), .rdup_out(a9_wr[524]), .rdlo_out(a9_wr[526]));
			radix2 #(.width(width)) rd_st8_525  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[525]), .rdlo_in(a8_wr[527]),  .coef_in(coef[256]), .rdup_out(a9_wr[525]), .rdlo_out(a9_wr[527]));
			radix2 #(.width(width)) rd_st8_528  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[528]), .rdlo_in(a8_wr[530]),  .coef_in(coef[0]), .rdup_out(a9_wr[528]), .rdlo_out(a9_wr[530]));
			radix2 #(.width(width)) rd_st8_529  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[529]), .rdlo_in(a8_wr[531]),  .coef_in(coef[256]), .rdup_out(a9_wr[529]), .rdlo_out(a9_wr[531]));
			radix2 #(.width(width)) rd_st8_532  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[532]), .rdlo_in(a8_wr[534]),  .coef_in(coef[0]), .rdup_out(a9_wr[532]), .rdlo_out(a9_wr[534]));
			radix2 #(.width(width)) rd_st8_533  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[533]), .rdlo_in(a8_wr[535]),  .coef_in(coef[256]), .rdup_out(a9_wr[533]), .rdlo_out(a9_wr[535]));
			radix2 #(.width(width)) rd_st8_536  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[536]), .rdlo_in(a8_wr[538]),  .coef_in(coef[0]), .rdup_out(a9_wr[536]), .rdlo_out(a9_wr[538]));
			radix2 #(.width(width)) rd_st8_537  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[537]), .rdlo_in(a8_wr[539]),  .coef_in(coef[256]), .rdup_out(a9_wr[537]), .rdlo_out(a9_wr[539]));
			radix2 #(.width(width)) rd_st8_540  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[540]), .rdlo_in(a8_wr[542]),  .coef_in(coef[0]), .rdup_out(a9_wr[540]), .rdlo_out(a9_wr[542]));
			radix2 #(.width(width)) rd_st8_541  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[541]), .rdlo_in(a8_wr[543]),  .coef_in(coef[256]), .rdup_out(a9_wr[541]), .rdlo_out(a9_wr[543]));
			radix2 #(.width(width)) rd_st8_544  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[544]), .rdlo_in(a8_wr[546]),  .coef_in(coef[0]), .rdup_out(a9_wr[544]), .rdlo_out(a9_wr[546]));
			radix2 #(.width(width)) rd_st8_545  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[545]), .rdlo_in(a8_wr[547]),  .coef_in(coef[256]), .rdup_out(a9_wr[545]), .rdlo_out(a9_wr[547]));
			radix2 #(.width(width)) rd_st8_548  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[548]), .rdlo_in(a8_wr[550]),  .coef_in(coef[0]), .rdup_out(a9_wr[548]), .rdlo_out(a9_wr[550]));
			radix2 #(.width(width)) rd_st8_549  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[549]), .rdlo_in(a8_wr[551]),  .coef_in(coef[256]), .rdup_out(a9_wr[549]), .rdlo_out(a9_wr[551]));
			radix2 #(.width(width)) rd_st8_552  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[552]), .rdlo_in(a8_wr[554]),  .coef_in(coef[0]), .rdup_out(a9_wr[552]), .rdlo_out(a9_wr[554]));
			radix2 #(.width(width)) rd_st8_553  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[553]), .rdlo_in(a8_wr[555]),  .coef_in(coef[256]), .rdup_out(a9_wr[553]), .rdlo_out(a9_wr[555]));
			radix2 #(.width(width)) rd_st8_556  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[556]), .rdlo_in(a8_wr[558]),  .coef_in(coef[0]), .rdup_out(a9_wr[556]), .rdlo_out(a9_wr[558]));
			radix2 #(.width(width)) rd_st8_557  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[557]), .rdlo_in(a8_wr[559]),  .coef_in(coef[256]), .rdup_out(a9_wr[557]), .rdlo_out(a9_wr[559]));
			radix2 #(.width(width)) rd_st8_560  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[560]), .rdlo_in(a8_wr[562]),  .coef_in(coef[0]), .rdup_out(a9_wr[560]), .rdlo_out(a9_wr[562]));
			radix2 #(.width(width)) rd_st8_561  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[561]), .rdlo_in(a8_wr[563]),  .coef_in(coef[256]), .rdup_out(a9_wr[561]), .rdlo_out(a9_wr[563]));
			radix2 #(.width(width)) rd_st8_564  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[564]), .rdlo_in(a8_wr[566]),  .coef_in(coef[0]), .rdup_out(a9_wr[564]), .rdlo_out(a9_wr[566]));
			radix2 #(.width(width)) rd_st8_565  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[565]), .rdlo_in(a8_wr[567]),  .coef_in(coef[256]), .rdup_out(a9_wr[565]), .rdlo_out(a9_wr[567]));
			radix2 #(.width(width)) rd_st8_568  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[568]), .rdlo_in(a8_wr[570]),  .coef_in(coef[0]), .rdup_out(a9_wr[568]), .rdlo_out(a9_wr[570]));
			radix2 #(.width(width)) rd_st8_569  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[569]), .rdlo_in(a8_wr[571]),  .coef_in(coef[256]), .rdup_out(a9_wr[569]), .rdlo_out(a9_wr[571]));
			radix2 #(.width(width)) rd_st8_572  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[572]), .rdlo_in(a8_wr[574]),  .coef_in(coef[0]), .rdup_out(a9_wr[572]), .rdlo_out(a9_wr[574]));
			radix2 #(.width(width)) rd_st8_573  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[573]), .rdlo_in(a8_wr[575]),  .coef_in(coef[256]), .rdup_out(a9_wr[573]), .rdlo_out(a9_wr[575]));
			radix2 #(.width(width)) rd_st8_576  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[576]), .rdlo_in(a8_wr[578]),  .coef_in(coef[0]), .rdup_out(a9_wr[576]), .rdlo_out(a9_wr[578]));
			radix2 #(.width(width)) rd_st8_577  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[577]), .rdlo_in(a8_wr[579]),  .coef_in(coef[256]), .rdup_out(a9_wr[577]), .rdlo_out(a9_wr[579]));
			radix2 #(.width(width)) rd_st8_580  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[580]), .rdlo_in(a8_wr[582]),  .coef_in(coef[0]), .rdup_out(a9_wr[580]), .rdlo_out(a9_wr[582]));
			radix2 #(.width(width)) rd_st8_581  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[581]), .rdlo_in(a8_wr[583]),  .coef_in(coef[256]), .rdup_out(a9_wr[581]), .rdlo_out(a9_wr[583]));
			radix2 #(.width(width)) rd_st8_584  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[584]), .rdlo_in(a8_wr[586]),  .coef_in(coef[0]), .rdup_out(a9_wr[584]), .rdlo_out(a9_wr[586]));
			radix2 #(.width(width)) rd_st8_585  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[585]), .rdlo_in(a8_wr[587]),  .coef_in(coef[256]), .rdup_out(a9_wr[585]), .rdlo_out(a9_wr[587]));
			radix2 #(.width(width)) rd_st8_588  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[588]), .rdlo_in(a8_wr[590]),  .coef_in(coef[0]), .rdup_out(a9_wr[588]), .rdlo_out(a9_wr[590]));
			radix2 #(.width(width)) rd_st8_589  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[589]), .rdlo_in(a8_wr[591]),  .coef_in(coef[256]), .rdup_out(a9_wr[589]), .rdlo_out(a9_wr[591]));
			radix2 #(.width(width)) rd_st8_592  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[592]), .rdlo_in(a8_wr[594]),  .coef_in(coef[0]), .rdup_out(a9_wr[592]), .rdlo_out(a9_wr[594]));
			radix2 #(.width(width)) rd_st8_593  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[593]), .rdlo_in(a8_wr[595]),  .coef_in(coef[256]), .rdup_out(a9_wr[593]), .rdlo_out(a9_wr[595]));
			radix2 #(.width(width)) rd_st8_596  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[596]), .rdlo_in(a8_wr[598]),  .coef_in(coef[0]), .rdup_out(a9_wr[596]), .rdlo_out(a9_wr[598]));
			radix2 #(.width(width)) rd_st8_597  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[597]), .rdlo_in(a8_wr[599]),  .coef_in(coef[256]), .rdup_out(a9_wr[597]), .rdlo_out(a9_wr[599]));
			radix2 #(.width(width)) rd_st8_600  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[600]), .rdlo_in(a8_wr[602]),  .coef_in(coef[0]), .rdup_out(a9_wr[600]), .rdlo_out(a9_wr[602]));
			radix2 #(.width(width)) rd_st8_601  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[601]), .rdlo_in(a8_wr[603]),  .coef_in(coef[256]), .rdup_out(a9_wr[601]), .rdlo_out(a9_wr[603]));
			radix2 #(.width(width)) rd_st8_604  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[604]), .rdlo_in(a8_wr[606]),  .coef_in(coef[0]), .rdup_out(a9_wr[604]), .rdlo_out(a9_wr[606]));
			radix2 #(.width(width)) rd_st8_605  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[605]), .rdlo_in(a8_wr[607]),  .coef_in(coef[256]), .rdup_out(a9_wr[605]), .rdlo_out(a9_wr[607]));
			radix2 #(.width(width)) rd_st8_608  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[608]), .rdlo_in(a8_wr[610]),  .coef_in(coef[0]), .rdup_out(a9_wr[608]), .rdlo_out(a9_wr[610]));
			radix2 #(.width(width)) rd_st8_609  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[609]), .rdlo_in(a8_wr[611]),  .coef_in(coef[256]), .rdup_out(a9_wr[609]), .rdlo_out(a9_wr[611]));
			radix2 #(.width(width)) rd_st8_612  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[612]), .rdlo_in(a8_wr[614]),  .coef_in(coef[0]), .rdup_out(a9_wr[612]), .rdlo_out(a9_wr[614]));
			radix2 #(.width(width)) rd_st8_613  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[613]), .rdlo_in(a8_wr[615]),  .coef_in(coef[256]), .rdup_out(a9_wr[613]), .rdlo_out(a9_wr[615]));
			radix2 #(.width(width)) rd_st8_616  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[616]), .rdlo_in(a8_wr[618]),  .coef_in(coef[0]), .rdup_out(a9_wr[616]), .rdlo_out(a9_wr[618]));
			radix2 #(.width(width)) rd_st8_617  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[617]), .rdlo_in(a8_wr[619]),  .coef_in(coef[256]), .rdup_out(a9_wr[617]), .rdlo_out(a9_wr[619]));
			radix2 #(.width(width)) rd_st8_620  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[620]), .rdlo_in(a8_wr[622]),  .coef_in(coef[0]), .rdup_out(a9_wr[620]), .rdlo_out(a9_wr[622]));
			radix2 #(.width(width)) rd_st8_621  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[621]), .rdlo_in(a8_wr[623]),  .coef_in(coef[256]), .rdup_out(a9_wr[621]), .rdlo_out(a9_wr[623]));
			radix2 #(.width(width)) rd_st8_624  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[624]), .rdlo_in(a8_wr[626]),  .coef_in(coef[0]), .rdup_out(a9_wr[624]), .rdlo_out(a9_wr[626]));
			radix2 #(.width(width)) rd_st8_625  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[625]), .rdlo_in(a8_wr[627]),  .coef_in(coef[256]), .rdup_out(a9_wr[625]), .rdlo_out(a9_wr[627]));
			radix2 #(.width(width)) rd_st8_628  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[628]), .rdlo_in(a8_wr[630]),  .coef_in(coef[0]), .rdup_out(a9_wr[628]), .rdlo_out(a9_wr[630]));
			radix2 #(.width(width)) rd_st8_629  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[629]), .rdlo_in(a8_wr[631]),  .coef_in(coef[256]), .rdup_out(a9_wr[629]), .rdlo_out(a9_wr[631]));
			radix2 #(.width(width)) rd_st8_632  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[632]), .rdlo_in(a8_wr[634]),  .coef_in(coef[0]), .rdup_out(a9_wr[632]), .rdlo_out(a9_wr[634]));
			radix2 #(.width(width)) rd_st8_633  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[633]), .rdlo_in(a8_wr[635]),  .coef_in(coef[256]), .rdup_out(a9_wr[633]), .rdlo_out(a9_wr[635]));
			radix2 #(.width(width)) rd_st8_636  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[636]), .rdlo_in(a8_wr[638]),  .coef_in(coef[0]), .rdup_out(a9_wr[636]), .rdlo_out(a9_wr[638]));
			radix2 #(.width(width)) rd_st8_637  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[637]), .rdlo_in(a8_wr[639]),  .coef_in(coef[256]), .rdup_out(a9_wr[637]), .rdlo_out(a9_wr[639]));
			radix2 #(.width(width)) rd_st8_640  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[640]), .rdlo_in(a8_wr[642]),  .coef_in(coef[0]), .rdup_out(a9_wr[640]), .rdlo_out(a9_wr[642]));
			radix2 #(.width(width)) rd_st8_641  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[641]), .rdlo_in(a8_wr[643]),  .coef_in(coef[256]), .rdup_out(a9_wr[641]), .rdlo_out(a9_wr[643]));
			radix2 #(.width(width)) rd_st8_644  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[644]), .rdlo_in(a8_wr[646]),  .coef_in(coef[0]), .rdup_out(a9_wr[644]), .rdlo_out(a9_wr[646]));
			radix2 #(.width(width)) rd_st8_645  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[645]), .rdlo_in(a8_wr[647]),  .coef_in(coef[256]), .rdup_out(a9_wr[645]), .rdlo_out(a9_wr[647]));
			radix2 #(.width(width)) rd_st8_648  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[648]), .rdlo_in(a8_wr[650]),  .coef_in(coef[0]), .rdup_out(a9_wr[648]), .rdlo_out(a9_wr[650]));
			radix2 #(.width(width)) rd_st8_649  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[649]), .rdlo_in(a8_wr[651]),  .coef_in(coef[256]), .rdup_out(a9_wr[649]), .rdlo_out(a9_wr[651]));
			radix2 #(.width(width)) rd_st8_652  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[652]), .rdlo_in(a8_wr[654]),  .coef_in(coef[0]), .rdup_out(a9_wr[652]), .rdlo_out(a9_wr[654]));
			radix2 #(.width(width)) rd_st8_653  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[653]), .rdlo_in(a8_wr[655]),  .coef_in(coef[256]), .rdup_out(a9_wr[653]), .rdlo_out(a9_wr[655]));
			radix2 #(.width(width)) rd_st8_656  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[656]), .rdlo_in(a8_wr[658]),  .coef_in(coef[0]), .rdup_out(a9_wr[656]), .rdlo_out(a9_wr[658]));
			radix2 #(.width(width)) rd_st8_657  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[657]), .rdlo_in(a8_wr[659]),  .coef_in(coef[256]), .rdup_out(a9_wr[657]), .rdlo_out(a9_wr[659]));
			radix2 #(.width(width)) rd_st8_660  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[660]), .rdlo_in(a8_wr[662]),  .coef_in(coef[0]), .rdup_out(a9_wr[660]), .rdlo_out(a9_wr[662]));
			radix2 #(.width(width)) rd_st8_661  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[661]), .rdlo_in(a8_wr[663]),  .coef_in(coef[256]), .rdup_out(a9_wr[661]), .rdlo_out(a9_wr[663]));
			radix2 #(.width(width)) rd_st8_664  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[664]), .rdlo_in(a8_wr[666]),  .coef_in(coef[0]), .rdup_out(a9_wr[664]), .rdlo_out(a9_wr[666]));
			radix2 #(.width(width)) rd_st8_665  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[665]), .rdlo_in(a8_wr[667]),  .coef_in(coef[256]), .rdup_out(a9_wr[665]), .rdlo_out(a9_wr[667]));
			radix2 #(.width(width)) rd_st8_668  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[668]), .rdlo_in(a8_wr[670]),  .coef_in(coef[0]), .rdup_out(a9_wr[668]), .rdlo_out(a9_wr[670]));
			radix2 #(.width(width)) rd_st8_669  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[669]), .rdlo_in(a8_wr[671]),  .coef_in(coef[256]), .rdup_out(a9_wr[669]), .rdlo_out(a9_wr[671]));
			radix2 #(.width(width)) rd_st8_672  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[672]), .rdlo_in(a8_wr[674]),  .coef_in(coef[0]), .rdup_out(a9_wr[672]), .rdlo_out(a9_wr[674]));
			radix2 #(.width(width)) rd_st8_673  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[673]), .rdlo_in(a8_wr[675]),  .coef_in(coef[256]), .rdup_out(a9_wr[673]), .rdlo_out(a9_wr[675]));
			radix2 #(.width(width)) rd_st8_676  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[676]), .rdlo_in(a8_wr[678]),  .coef_in(coef[0]), .rdup_out(a9_wr[676]), .rdlo_out(a9_wr[678]));
			radix2 #(.width(width)) rd_st8_677  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[677]), .rdlo_in(a8_wr[679]),  .coef_in(coef[256]), .rdup_out(a9_wr[677]), .rdlo_out(a9_wr[679]));
			radix2 #(.width(width)) rd_st8_680  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[680]), .rdlo_in(a8_wr[682]),  .coef_in(coef[0]), .rdup_out(a9_wr[680]), .rdlo_out(a9_wr[682]));
			radix2 #(.width(width)) rd_st8_681  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[681]), .rdlo_in(a8_wr[683]),  .coef_in(coef[256]), .rdup_out(a9_wr[681]), .rdlo_out(a9_wr[683]));
			radix2 #(.width(width)) rd_st8_684  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[684]), .rdlo_in(a8_wr[686]),  .coef_in(coef[0]), .rdup_out(a9_wr[684]), .rdlo_out(a9_wr[686]));
			radix2 #(.width(width)) rd_st8_685  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[685]), .rdlo_in(a8_wr[687]),  .coef_in(coef[256]), .rdup_out(a9_wr[685]), .rdlo_out(a9_wr[687]));
			radix2 #(.width(width)) rd_st8_688  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[688]), .rdlo_in(a8_wr[690]),  .coef_in(coef[0]), .rdup_out(a9_wr[688]), .rdlo_out(a9_wr[690]));
			radix2 #(.width(width)) rd_st8_689  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[689]), .rdlo_in(a8_wr[691]),  .coef_in(coef[256]), .rdup_out(a9_wr[689]), .rdlo_out(a9_wr[691]));
			radix2 #(.width(width)) rd_st8_692  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[692]), .rdlo_in(a8_wr[694]),  .coef_in(coef[0]), .rdup_out(a9_wr[692]), .rdlo_out(a9_wr[694]));
			radix2 #(.width(width)) rd_st8_693  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[693]), .rdlo_in(a8_wr[695]),  .coef_in(coef[256]), .rdup_out(a9_wr[693]), .rdlo_out(a9_wr[695]));
			radix2 #(.width(width)) rd_st8_696  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[696]), .rdlo_in(a8_wr[698]),  .coef_in(coef[0]), .rdup_out(a9_wr[696]), .rdlo_out(a9_wr[698]));
			radix2 #(.width(width)) rd_st8_697  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[697]), .rdlo_in(a8_wr[699]),  .coef_in(coef[256]), .rdup_out(a9_wr[697]), .rdlo_out(a9_wr[699]));
			radix2 #(.width(width)) rd_st8_700  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[700]), .rdlo_in(a8_wr[702]),  .coef_in(coef[0]), .rdup_out(a9_wr[700]), .rdlo_out(a9_wr[702]));
			radix2 #(.width(width)) rd_st8_701  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[701]), .rdlo_in(a8_wr[703]),  .coef_in(coef[256]), .rdup_out(a9_wr[701]), .rdlo_out(a9_wr[703]));
			radix2 #(.width(width)) rd_st8_704  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[704]), .rdlo_in(a8_wr[706]),  .coef_in(coef[0]), .rdup_out(a9_wr[704]), .rdlo_out(a9_wr[706]));
			radix2 #(.width(width)) rd_st8_705  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[705]), .rdlo_in(a8_wr[707]),  .coef_in(coef[256]), .rdup_out(a9_wr[705]), .rdlo_out(a9_wr[707]));
			radix2 #(.width(width)) rd_st8_708  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[708]), .rdlo_in(a8_wr[710]),  .coef_in(coef[0]), .rdup_out(a9_wr[708]), .rdlo_out(a9_wr[710]));
			radix2 #(.width(width)) rd_st8_709  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[709]), .rdlo_in(a8_wr[711]),  .coef_in(coef[256]), .rdup_out(a9_wr[709]), .rdlo_out(a9_wr[711]));
			radix2 #(.width(width)) rd_st8_712  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[712]), .rdlo_in(a8_wr[714]),  .coef_in(coef[0]), .rdup_out(a9_wr[712]), .rdlo_out(a9_wr[714]));
			radix2 #(.width(width)) rd_st8_713  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[713]), .rdlo_in(a8_wr[715]),  .coef_in(coef[256]), .rdup_out(a9_wr[713]), .rdlo_out(a9_wr[715]));
			radix2 #(.width(width)) rd_st8_716  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[716]), .rdlo_in(a8_wr[718]),  .coef_in(coef[0]), .rdup_out(a9_wr[716]), .rdlo_out(a9_wr[718]));
			radix2 #(.width(width)) rd_st8_717  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[717]), .rdlo_in(a8_wr[719]),  .coef_in(coef[256]), .rdup_out(a9_wr[717]), .rdlo_out(a9_wr[719]));
			radix2 #(.width(width)) rd_st8_720  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[720]), .rdlo_in(a8_wr[722]),  .coef_in(coef[0]), .rdup_out(a9_wr[720]), .rdlo_out(a9_wr[722]));
			radix2 #(.width(width)) rd_st8_721  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[721]), .rdlo_in(a8_wr[723]),  .coef_in(coef[256]), .rdup_out(a9_wr[721]), .rdlo_out(a9_wr[723]));
			radix2 #(.width(width)) rd_st8_724  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[724]), .rdlo_in(a8_wr[726]),  .coef_in(coef[0]), .rdup_out(a9_wr[724]), .rdlo_out(a9_wr[726]));
			radix2 #(.width(width)) rd_st8_725  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[725]), .rdlo_in(a8_wr[727]),  .coef_in(coef[256]), .rdup_out(a9_wr[725]), .rdlo_out(a9_wr[727]));
			radix2 #(.width(width)) rd_st8_728  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[728]), .rdlo_in(a8_wr[730]),  .coef_in(coef[0]), .rdup_out(a9_wr[728]), .rdlo_out(a9_wr[730]));
			radix2 #(.width(width)) rd_st8_729  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[729]), .rdlo_in(a8_wr[731]),  .coef_in(coef[256]), .rdup_out(a9_wr[729]), .rdlo_out(a9_wr[731]));
			radix2 #(.width(width)) rd_st8_732  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[732]), .rdlo_in(a8_wr[734]),  .coef_in(coef[0]), .rdup_out(a9_wr[732]), .rdlo_out(a9_wr[734]));
			radix2 #(.width(width)) rd_st8_733  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[733]), .rdlo_in(a8_wr[735]),  .coef_in(coef[256]), .rdup_out(a9_wr[733]), .rdlo_out(a9_wr[735]));
			radix2 #(.width(width)) rd_st8_736  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[736]), .rdlo_in(a8_wr[738]),  .coef_in(coef[0]), .rdup_out(a9_wr[736]), .rdlo_out(a9_wr[738]));
			radix2 #(.width(width)) rd_st8_737  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[737]), .rdlo_in(a8_wr[739]),  .coef_in(coef[256]), .rdup_out(a9_wr[737]), .rdlo_out(a9_wr[739]));
			radix2 #(.width(width)) rd_st8_740  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[740]), .rdlo_in(a8_wr[742]),  .coef_in(coef[0]), .rdup_out(a9_wr[740]), .rdlo_out(a9_wr[742]));
			radix2 #(.width(width)) rd_st8_741  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[741]), .rdlo_in(a8_wr[743]),  .coef_in(coef[256]), .rdup_out(a9_wr[741]), .rdlo_out(a9_wr[743]));
			radix2 #(.width(width)) rd_st8_744  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[744]), .rdlo_in(a8_wr[746]),  .coef_in(coef[0]), .rdup_out(a9_wr[744]), .rdlo_out(a9_wr[746]));
			radix2 #(.width(width)) rd_st8_745  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[745]), .rdlo_in(a8_wr[747]),  .coef_in(coef[256]), .rdup_out(a9_wr[745]), .rdlo_out(a9_wr[747]));
			radix2 #(.width(width)) rd_st8_748  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[748]), .rdlo_in(a8_wr[750]),  .coef_in(coef[0]), .rdup_out(a9_wr[748]), .rdlo_out(a9_wr[750]));
			radix2 #(.width(width)) rd_st8_749  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[749]), .rdlo_in(a8_wr[751]),  .coef_in(coef[256]), .rdup_out(a9_wr[749]), .rdlo_out(a9_wr[751]));
			radix2 #(.width(width)) rd_st8_752  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[752]), .rdlo_in(a8_wr[754]),  .coef_in(coef[0]), .rdup_out(a9_wr[752]), .rdlo_out(a9_wr[754]));
			radix2 #(.width(width)) rd_st8_753  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[753]), .rdlo_in(a8_wr[755]),  .coef_in(coef[256]), .rdup_out(a9_wr[753]), .rdlo_out(a9_wr[755]));
			radix2 #(.width(width)) rd_st8_756  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[756]), .rdlo_in(a8_wr[758]),  .coef_in(coef[0]), .rdup_out(a9_wr[756]), .rdlo_out(a9_wr[758]));
			radix2 #(.width(width)) rd_st8_757  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[757]), .rdlo_in(a8_wr[759]),  .coef_in(coef[256]), .rdup_out(a9_wr[757]), .rdlo_out(a9_wr[759]));
			radix2 #(.width(width)) rd_st8_760  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[760]), .rdlo_in(a8_wr[762]),  .coef_in(coef[0]), .rdup_out(a9_wr[760]), .rdlo_out(a9_wr[762]));
			radix2 #(.width(width)) rd_st8_761  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[761]), .rdlo_in(a8_wr[763]),  .coef_in(coef[256]), .rdup_out(a9_wr[761]), .rdlo_out(a9_wr[763]));
			radix2 #(.width(width)) rd_st8_764  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[764]), .rdlo_in(a8_wr[766]),  .coef_in(coef[0]), .rdup_out(a9_wr[764]), .rdlo_out(a9_wr[766]));
			radix2 #(.width(width)) rd_st8_765  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[765]), .rdlo_in(a8_wr[767]),  .coef_in(coef[256]), .rdup_out(a9_wr[765]), .rdlo_out(a9_wr[767]));
			radix2 #(.width(width)) rd_st8_768  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[768]), .rdlo_in(a8_wr[770]),  .coef_in(coef[0]), .rdup_out(a9_wr[768]), .rdlo_out(a9_wr[770]));
			radix2 #(.width(width)) rd_st8_769  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[769]), .rdlo_in(a8_wr[771]),  .coef_in(coef[256]), .rdup_out(a9_wr[769]), .rdlo_out(a9_wr[771]));
			radix2 #(.width(width)) rd_st8_772  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[772]), .rdlo_in(a8_wr[774]),  .coef_in(coef[0]), .rdup_out(a9_wr[772]), .rdlo_out(a9_wr[774]));
			radix2 #(.width(width)) rd_st8_773  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[773]), .rdlo_in(a8_wr[775]),  .coef_in(coef[256]), .rdup_out(a9_wr[773]), .rdlo_out(a9_wr[775]));
			radix2 #(.width(width)) rd_st8_776  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[776]), .rdlo_in(a8_wr[778]),  .coef_in(coef[0]), .rdup_out(a9_wr[776]), .rdlo_out(a9_wr[778]));
			radix2 #(.width(width)) rd_st8_777  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[777]), .rdlo_in(a8_wr[779]),  .coef_in(coef[256]), .rdup_out(a9_wr[777]), .rdlo_out(a9_wr[779]));
			radix2 #(.width(width)) rd_st8_780  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[780]), .rdlo_in(a8_wr[782]),  .coef_in(coef[0]), .rdup_out(a9_wr[780]), .rdlo_out(a9_wr[782]));
			radix2 #(.width(width)) rd_st8_781  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[781]), .rdlo_in(a8_wr[783]),  .coef_in(coef[256]), .rdup_out(a9_wr[781]), .rdlo_out(a9_wr[783]));
			radix2 #(.width(width)) rd_st8_784  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[784]), .rdlo_in(a8_wr[786]),  .coef_in(coef[0]), .rdup_out(a9_wr[784]), .rdlo_out(a9_wr[786]));
			radix2 #(.width(width)) rd_st8_785  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[785]), .rdlo_in(a8_wr[787]),  .coef_in(coef[256]), .rdup_out(a9_wr[785]), .rdlo_out(a9_wr[787]));
			radix2 #(.width(width)) rd_st8_788  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[788]), .rdlo_in(a8_wr[790]),  .coef_in(coef[0]), .rdup_out(a9_wr[788]), .rdlo_out(a9_wr[790]));
			radix2 #(.width(width)) rd_st8_789  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[789]), .rdlo_in(a8_wr[791]),  .coef_in(coef[256]), .rdup_out(a9_wr[789]), .rdlo_out(a9_wr[791]));
			radix2 #(.width(width)) rd_st8_792  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[792]), .rdlo_in(a8_wr[794]),  .coef_in(coef[0]), .rdup_out(a9_wr[792]), .rdlo_out(a9_wr[794]));
			radix2 #(.width(width)) rd_st8_793  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[793]), .rdlo_in(a8_wr[795]),  .coef_in(coef[256]), .rdup_out(a9_wr[793]), .rdlo_out(a9_wr[795]));
			radix2 #(.width(width)) rd_st8_796  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[796]), .rdlo_in(a8_wr[798]),  .coef_in(coef[0]), .rdup_out(a9_wr[796]), .rdlo_out(a9_wr[798]));
			radix2 #(.width(width)) rd_st8_797  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[797]), .rdlo_in(a8_wr[799]),  .coef_in(coef[256]), .rdup_out(a9_wr[797]), .rdlo_out(a9_wr[799]));
			radix2 #(.width(width)) rd_st8_800  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[800]), .rdlo_in(a8_wr[802]),  .coef_in(coef[0]), .rdup_out(a9_wr[800]), .rdlo_out(a9_wr[802]));
			radix2 #(.width(width)) rd_st8_801  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[801]), .rdlo_in(a8_wr[803]),  .coef_in(coef[256]), .rdup_out(a9_wr[801]), .rdlo_out(a9_wr[803]));
			radix2 #(.width(width)) rd_st8_804  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[804]), .rdlo_in(a8_wr[806]),  .coef_in(coef[0]), .rdup_out(a9_wr[804]), .rdlo_out(a9_wr[806]));
			radix2 #(.width(width)) rd_st8_805  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[805]), .rdlo_in(a8_wr[807]),  .coef_in(coef[256]), .rdup_out(a9_wr[805]), .rdlo_out(a9_wr[807]));
			radix2 #(.width(width)) rd_st8_808  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[808]), .rdlo_in(a8_wr[810]),  .coef_in(coef[0]), .rdup_out(a9_wr[808]), .rdlo_out(a9_wr[810]));
			radix2 #(.width(width)) rd_st8_809  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[809]), .rdlo_in(a8_wr[811]),  .coef_in(coef[256]), .rdup_out(a9_wr[809]), .rdlo_out(a9_wr[811]));
			radix2 #(.width(width)) rd_st8_812  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[812]), .rdlo_in(a8_wr[814]),  .coef_in(coef[0]), .rdup_out(a9_wr[812]), .rdlo_out(a9_wr[814]));
			radix2 #(.width(width)) rd_st8_813  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[813]), .rdlo_in(a8_wr[815]),  .coef_in(coef[256]), .rdup_out(a9_wr[813]), .rdlo_out(a9_wr[815]));
			radix2 #(.width(width)) rd_st8_816  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[816]), .rdlo_in(a8_wr[818]),  .coef_in(coef[0]), .rdup_out(a9_wr[816]), .rdlo_out(a9_wr[818]));
			radix2 #(.width(width)) rd_st8_817  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[817]), .rdlo_in(a8_wr[819]),  .coef_in(coef[256]), .rdup_out(a9_wr[817]), .rdlo_out(a9_wr[819]));
			radix2 #(.width(width)) rd_st8_820  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[820]), .rdlo_in(a8_wr[822]),  .coef_in(coef[0]), .rdup_out(a9_wr[820]), .rdlo_out(a9_wr[822]));
			radix2 #(.width(width)) rd_st8_821  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[821]), .rdlo_in(a8_wr[823]),  .coef_in(coef[256]), .rdup_out(a9_wr[821]), .rdlo_out(a9_wr[823]));
			radix2 #(.width(width)) rd_st8_824  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[824]), .rdlo_in(a8_wr[826]),  .coef_in(coef[0]), .rdup_out(a9_wr[824]), .rdlo_out(a9_wr[826]));
			radix2 #(.width(width)) rd_st8_825  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[825]), .rdlo_in(a8_wr[827]),  .coef_in(coef[256]), .rdup_out(a9_wr[825]), .rdlo_out(a9_wr[827]));
			radix2 #(.width(width)) rd_st8_828  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[828]), .rdlo_in(a8_wr[830]),  .coef_in(coef[0]), .rdup_out(a9_wr[828]), .rdlo_out(a9_wr[830]));
			radix2 #(.width(width)) rd_st8_829  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[829]), .rdlo_in(a8_wr[831]),  .coef_in(coef[256]), .rdup_out(a9_wr[829]), .rdlo_out(a9_wr[831]));
			radix2 #(.width(width)) rd_st8_832  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[832]), .rdlo_in(a8_wr[834]),  .coef_in(coef[0]), .rdup_out(a9_wr[832]), .rdlo_out(a9_wr[834]));
			radix2 #(.width(width)) rd_st8_833  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[833]), .rdlo_in(a8_wr[835]),  .coef_in(coef[256]), .rdup_out(a9_wr[833]), .rdlo_out(a9_wr[835]));
			radix2 #(.width(width)) rd_st8_836  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[836]), .rdlo_in(a8_wr[838]),  .coef_in(coef[0]), .rdup_out(a9_wr[836]), .rdlo_out(a9_wr[838]));
			radix2 #(.width(width)) rd_st8_837  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[837]), .rdlo_in(a8_wr[839]),  .coef_in(coef[256]), .rdup_out(a9_wr[837]), .rdlo_out(a9_wr[839]));
			radix2 #(.width(width)) rd_st8_840  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[840]), .rdlo_in(a8_wr[842]),  .coef_in(coef[0]), .rdup_out(a9_wr[840]), .rdlo_out(a9_wr[842]));
			radix2 #(.width(width)) rd_st8_841  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[841]), .rdlo_in(a8_wr[843]),  .coef_in(coef[256]), .rdup_out(a9_wr[841]), .rdlo_out(a9_wr[843]));
			radix2 #(.width(width)) rd_st8_844  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[844]), .rdlo_in(a8_wr[846]),  .coef_in(coef[0]), .rdup_out(a9_wr[844]), .rdlo_out(a9_wr[846]));
			radix2 #(.width(width)) rd_st8_845  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[845]), .rdlo_in(a8_wr[847]),  .coef_in(coef[256]), .rdup_out(a9_wr[845]), .rdlo_out(a9_wr[847]));
			radix2 #(.width(width)) rd_st8_848  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[848]), .rdlo_in(a8_wr[850]),  .coef_in(coef[0]), .rdup_out(a9_wr[848]), .rdlo_out(a9_wr[850]));
			radix2 #(.width(width)) rd_st8_849  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[849]), .rdlo_in(a8_wr[851]),  .coef_in(coef[256]), .rdup_out(a9_wr[849]), .rdlo_out(a9_wr[851]));
			radix2 #(.width(width)) rd_st8_852  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[852]), .rdlo_in(a8_wr[854]),  .coef_in(coef[0]), .rdup_out(a9_wr[852]), .rdlo_out(a9_wr[854]));
			radix2 #(.width(width)) rd_st8_853  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[853]), .rdlo_in(a8_wr[855]),  .coef_in(coef[256]), .rdup_out(a9_wr[853]), .rdlo_out(a9_wr[855]));
			radix2 #(.width(width)) rd_st8_856  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[856]), .rdlo_in(a8_wr[858]),  .coef_in(coef[0]), .rdup_out(a9_wr[856]), .rdlo_out(a9_wr[858]));
			radix2 #(.width(width)) rd_st8_857  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[857]), .rdlo_in(a8_wr[859]),  .coef_in(coef[256]), .rdup_out(a9_wr[857]), .rdlo_out(a9_wr[859]));
			radix2 #(.width(width)) rd_st8_860  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[860]), .rdlo_in(a8_wr[862]),  .coef_in(coef[0]), .rdup_out(a9_wr[860]), .rdlo_out(a9_wr[862]));
			radix2 #(.width(width)) rd_st8_861  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[861]), .rdlo_in(a8_wr[863]),  .coef_in(coef[256]), .rdup_out(a9_wr[861]), .rdlo_out(a9_wr[863]));
			radix2 #(.width(width)) rd_st8_864  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[864]), .rdlo_in(a8_wr[866]),  .coef_in(coef[0]), .rdup_out(a9_wr[864]), .rdlo_out(a9_wr[866]));
			radix2 #(.width(width)) rd_st8_865  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[865]), .rdlo_in(a8_wr[867]),  .coef_in(coef[256]), .rdup_out(a9_wr[865]), .rdlo_out(a9_wr[867]));
			radix2 #(.width(width)) rd_st8_868  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[868]), .rdlo_in(a8_wr[870]),  .coef_in(coef[0]), .rdup_out(a9_wr[868]), .rdlo_out(a9_wr[870]));
			radix2 #(.width(width)) rd_st8_869  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[869]), .rdlo_in(a8_wr[871]),  .coef_in(coef[256]), .rdup_out(a9_wr[869]), .rdlo_out(a9_wr[871]));
			radix2 #(.width(width)) rd_st8_872  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[872]), .rdlo_in(a8_wr[874]),  .coef_in(coef[0]), .rdup_out(a9_wr[872]), .rdlo_out(a9_wr[874]));
			radix2 #(.width(width)) rd_st8_873  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[873]), .rdlo_in(a8_wr[875]),  .coef_in(coef[256]), .rdup_out(a9_wr[873]), .rdlo_out(a9_wr[875]));
			radix2 #(.width(width)) rd_st8_876  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[876]), .rdlo_in(a8_wr[878]),  .coef_in(coef[0]), .rdup_out(a9_wr[876]), .rdlo_out(a9_wr[878]));
			radix2 #(.width(width)) rd_st8_877  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[877]), .rdlo_in(a8_wr[879]),  .coef_in(coef[256]), .rdup_out(a9_wr[877]), .rdlo_out(a9_wr[879]));
			radix2 #(.width(width)) rd_st8_880  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[880]), .rdlo_in(a8_wr[882]),  .coef_in(coef[0]), .rdup_out(a9_wr[880]), .rdlo_out(a9_wr[882]));
			radix2 #(.width(width)) rd_st8_881  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[881]), .rdlo_in(a8_wr[883]),  .coef_in(coef[256]), .rdup_out(a9_wr[881]), .rdlo_out(a9_wr[883]));
			radix2 #(.width(width)) rd_st8_884  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[884]), .rdlo_in(a8_wr[886]),  .coef_in(coef[0]), .rdup_out(a9_wr[884]), .rdlo_out(a9_wr[886]));
			radix2 #(.width(width)) rd_st8_885  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[885]), .rdlo_in(a8_wr[887]),  .coef_in(coef[256]), .rdup_out(a9_wr[885]), .rdlo_out(a9_wr[887]));
			radix2 #(.width(width)) rd_st8_888  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[888]), .rdlo_in(a8_wr[890]),  .coef_in(coef[0]), .rdup_out(a9_wr[888]), .rdlo_out(a9_wr[890]));
			radix2 #(.width(width)) rd_st8_889  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[889]), .rdlo_in(a8_wr[891]),  .coef_in(coef[256]), .rdup_out(a9_wr[889]), .rdlo_out(a9_wr[891]));
			radix2 #(.width(width)) rd_st8_892  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[892]), .rdlo_in(a8_wr[894]),  .coef_in(coef[0]), .rdup_out(a9_wr[892]), .rdlo_out(a9_wr[894]));
			radix2 #(.width(width)) rd_st8_893  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[893]), .rdlo_in(a8_wr[895]),  .coef_in(coef[256]), .rdup_out(a9_wr[893]), .rdlo_out(a9_wr[895]));
			radix2 #(.width(width)) rd_st8_896  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[896]), .rdlo_in(a8_wr[898]),  .coef_in(coef[0]), .rdup_out(a9_wr[896]), .rdlo_out(a9_wr[898]));
			radix2 #(.width(width)) rd_st8_897  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[897]), .rdlo_in(a8_wr[899]),  .coef_in(coef[256]), .rdup_out(a9_wr[897]), .rdlo_out(a9_wr[899]));
			radix2 #(.width(width)) rd_st8_900  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[900]), .rdlo_in(a8_wr[902]),  .coef_in(coef[0]), .rdup_out(a9_wr[900]), .rdlo_out(a9_wr[902]));
			radix2 #(.width(width)) rd_st8_901  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[901]), .rdlo_in(a8_wr[903]),  .coef_in(coef[256]), .rdup_out(a9_wr[901]), .rdlo_out(a9_wr[903]));
			radix2 #(.width(width)) rd_st8_904  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[904]), .rdlo_in(a8_wr[906]),  .coef_in(coef[0]), .rdup_out(a9_wr[904]), .rdlo_out(a9_wr[906]));
			radix2 #(.width(width)) rd_st8_905  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[905]), .rdlo_in(a8_wr[907]),  .coef_in(coef[256]), .rdup_out(a9_wr[905]), .rdlo_out(a9_wr[907]));
			radix2 #(.width(width)) rd_st8_908  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[908]), .rdlo_in(a8_wr[910]),  .coef_in(coef[0]), .rdup_out(a9_wr[908]), .rdlo_out(a9_wr[910]));
			radix2 #(.width(width)) rd_st8_909  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[909]), .rdlo_in(a8_wr[911]),  .coef_in(coef[256]), .rdup_out(a9_wr[909]), .rdlo_out(a9_wr[911]));
			radix2 #(.width(width)) rd_st8_912  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[912]), .rdlo_in(a8_wr[914]),  .coef_in(coef[0]), .rdup_out(a9_wr[912]), .rdlo_out(a9_wr[914]));
			radix2 #(.width(width)) rd_st8_913  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[913]), .rdlo_in(a8_wr[915]),  .coef_in(coef[256]), .rdup_out(a9_wr[913]), .rdlo_out(a9_wr[915]));
			radix2 #(.width(width)) rd_st8_916  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[916]), .rdlo_in(a8_wr[918]),  .coef_in(coef[0]), .rdup_out(a9_wr[916]), .rdlo_out(a9_wr[918]));
			radix2 #(.width(width)) rd_st8_917  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[917]), .rdlo_in(a8_wr[919]),  .coef_in(coef[256]), .rdup_out(a9_wr[917]), .rdlo_out(a9_wr[919]));
			radix2 #(.width(width)) rd_st8_920  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[920]), .rdlo_in(a8_wr[922]),  .coef_in(coef[0]), .rdup_out(a9_wr[920]), .rdlo_out(a9_wr[922]));
			radix2 #(.width(width)) rd_st8_921  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[921]), .rdlo_in(a8_wr[923]),  .coef_in(coef[256]), .rdup_out(a9_wr[921]), .rdlo_out(a9_wr[923]));
			radix2 #(.width(width)) rd_st8_924  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[924]), .rdlo_in(a8_wr[926]),  .coef_in(coef[0]), .rdup_out(a9_wr[924]), .rdlo_out(a9_wr[926]));
			radix2 #(.width(width)) rd_st8_925  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[925]), .rdlo_in(a8_wr[927]),  .coef_in(coef[256]), .rdup_out(a9_wr[925]), .rdlo_out(a9_wr[927]));
			radix2 #(.width(width)) rd_st8_928  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[928]), .rdlo_in(a8_wr[930]),  .coef_in(coef[0]), .rdup_out(a9_wr[928]), .rdlo_out(a9_wr[930]));
			radix2 #(.width(width)) rd_st8_929  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[929]), .rdlo_in(a8_wr[931]),  .coef_in(coef[256]), .rdup_out(a9_wr[929]), .rdlo_out(a9_wr[931]));
			radix2 #(.width(width)) rd_st8_932  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[932]), .rdlo_in(a8_wr[934]),  .coef_in(coef[0]), .rdup_out(a9_wr[932]), .rdlo_out(a9_wr[934]));
			radix2 #(.width(width)) rd_st8_933  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[933]), .rdlo_in(a8_wr[935]),  .coef_in(coef[256]), .rdup_out(a9_wr[933]), .rdlo_out(a9_wr[935]));
			radix2 #(.width(width)) rd_st8_936  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[936]), .rdlo_in(a8_wr[938]),  .coef_in(coef[0]), .rdup_out(a9_wr[936]), .rdlo_out(a9_wr[938]));
			radix2 #(.width(width)) rd_st8_937  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[937]), .rdlo_in(a8_wr[939]),  .coef_in(coef[256]), .rdup_out(a9_wr[937]), .rdlo_out(a9_wr[939]));
			radix2 #(.width(width)) rd_st8_940  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[940]), .rdlo_in(a8_wr[942]),  .coef_in(coef[0]), .rdup_out(a9_wr[940]), .rdlo_out(a9_wr[942]));
			radix2 #(.width(width)) rd_st8_941  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[941]), .rdlo_in(a8_wr[943]),  .coef_in(coef[256]), .rdup_out(a9_wr[941]), .rdlo_out(a9_wr[943]));
			radix2 #(.width(width)) rd_st8_944  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[944]), .rdlo_in(a8_wr[946]),  .coef_in(coef[0]), .rdup_out(a9_wr[944]), .rdlo_out(a9_wr[946]));
			radix2 #(.width(width)) rd_st8_945  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[945]), .rdlo_in(a8_wr[947]),  .coef_in(coef[256]), .rdup_out(a9_wr[945]), .rdlo_out(a9_wr[947]));
			radix2 #(.width(width)) rd_st8_948  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[948]), .rdlo_in(a8_wr[950]),  .coef_in(coef[0]), .rdup_out(a9_wr[948]), .rdlo_out(a9_wr[950]));
			radix2 #(.width(width)) rd_st8_949  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[949]), .rdlo_in(a8_wr[951]),  .coef_in(coef[256]), .rdup_out(a9_wr[949]), .rdlo_out(a9_wr[951]));
			radix2 #(.width(width)) rd_st8_952  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[952]), .rdlo_in(a8_wr[954]),  .coef_in(coef[0]), .rdup_out(a9_wr[952]), .rdlo_out(a9_wr[954]));
			radix2 #(.width(width)) rd_st8_953  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[953]), .rdlo_in(a8_wr[955]),  .coef_in(coef[256]), .rdup_out(a9_wr[953]), .rdlo_out(a9_wr[955]));
			radix2 #(.width(width)) rd_st8_956  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[956]), .rdlo_in(a8_wr[958]),  .coef_in(coef[0]), .rdup_out(a9_wr[956]), .rdlo_out(a9_wr[958]));
			radix2 #(.width(width)) rd_st8_957  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[957]), .rdlo_in(a8_wr[959]),  .coef_in(coef[256]), .rdup_out(a9_wr[957]), .rdlo_out(a9_wr[959]));
			radix2 #(.width(width)) rd_st8_960  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[960]), .rdlo_in(a8_wr[962]),  .coef_in(coef[0]), .rdup_out(a9_wr[960]), .rdlo_out(a9_wr[962]));
			radix2 #(.width(width)) rd_st8_961  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[961]), .rdlo_in(a8_wr[963]),  .coef_in(coef[256]), .rdup_out(a9_wr[961]), .rdlo_out(a9_wr[963]));
			radix2 #(.width(width)) rd_st8_964  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[964]), .rdlo_in(a8_wr[966]),  .coef_in(coef[0]), .rdup_out(a9_wr[964]), .rdlo_out(a9_wr[966]));
			radix2 #(.width(width)) rd_st8_965  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[965]), .rdlo_in(a8_wr[967]),  .coef_in(coef[256]), .rdup_out(a9_wr[965]), .rdlo_out(a9_wr[967]));
			radix2 #(.width(width)) rd_st8_968  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[968]), .rdlo_in(a8_wr[970]),  .coef_in(coef[0]), .rdup_out(a9_wr[968]), .rdlo_out(a9_wr[970]));
			radix2 #(.width(width)) rd_st8_969  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[969]), .rdlo_in(a8_wr[971]),  .coef_in(coef[256]), .rdup_out(a9_wr[969]), .rdlo_out(a9_wr[971]));
			radix2 #(.width(width)) rd_st8_972  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[972]), .rdlo_in(a8_wr[974]),  .coef_in(coef[0]), .rdup_out(a9_wr[972]), .rdlo_out(a9_wr[974]));
			radix2 #(.width(width)) rd_st8_973  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[973]), .rdlo_in(a8_wr[975]),  .coef_in(coef[256]), .rdup_out(a9_wr[973]), .rdlo_out(a9_wr[975]));
			radix2 #(.width(width)) rd_st8_976  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[976]), .rdlo_in(a8_wr[978]),  .coef_in(coef[0]), .rdup_out(a9_wr[976]), .rdlo_out(a9_wr[978]));
			radix2 #(.width(width)) rd_st8_977  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[977]), .rdlo_in(a8_wr[979]),  .coef_in(coef[256]), .rdup_out(a9_wr[977]), .rdlo_out(a9_wr[979]));
			radix2 #(.width(width)) rd_st8_980  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[980]), .rdlo_in(a8_wr[982]),  .coef_in(coef[0]), .rdup_out(a9_wr[980]), .rdlo_out(a9_wr[982]));
			radix2 #(.width(width)) rd_st8_981  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[981]), .rdlo_in(a8_wr[983]),  .coef_in(coef[256]), .rdup_out(a9_wr[981]), .rdlo_out(a9_wr[983]));
			radix2 #(.width(width)) rd_st8_984  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[984]), .rdlo_in(a8_wr[986]),  .coef_in(coef[0]), .rdup_out(a9_wr[984]), .rdlo_out(a9_wr[986]));
			radix2 #(.width(width)) rd_st8_985  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[985]), .rdlo_in(a8_wr[987]),  .coef_in(coef[256]), .rdup_out(a9_wr[985]), .rdlo_out(a9_wr[987]));
			radix2 #(.width(width)) rd_st8_988  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[988]), .rdlo_in(a8_wr[990]),  .coef_in(coef[0]), .rdup_out(a9_wr[988]), .rdlo_out(a9_wr[990]));
			radix2 #(.width(width)) rd_st8_989  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[989]), .rdlo_in(a8_wr[991]),  .coef_in(coef[256]), .rdup_out(a9_wr[989]), .rdlo_out(a9_wr[991]));
			radix2 #(.width(width)) rd_st8_992  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[992]), .rdlo_in(a8_wr[994]),  .coef_in(coef[0]), .rdup_out(a9_wr[992]), .rdlo_out(a9_wr[994]));
			radix2 #(.width(width)) rd_st8_993  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[993]), .rdlo_in(a8_wr[995]),  .coef_in(coef[256]), .rdup_out(a9_wr[993]), .rdlo_out(a9_wr[995]));
			radix2 #(.width(width)) rd_st8_996  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[996]), .rdlo_in(a8_wr[998]),  .coef_in(coef[0]), .rdup_out(a9_wr[996]), .rdlo_out(a9_wr[998]));
			radix2 #(.width(width)) rd_st8_997  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[997]), .rdlo_in(a8_wr[999]),  .coef_in(coef[256]), .rdup_out(a9_wr[997]), .rdlo_out(a9_wr[999]));
			radix2 #(.width(width)) rd_st8_1000  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1000]), .rdlo_in(a8_wr[1002]),  .coef_in(coef[0]), .rdup_out(a9_wr[1000]), .rdlo_out(a9_wr[1002]));
			radix2 #(.width(width)) rd_st8_1001  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1001]), .rdlo_in(a8_wr[1003]),  .coef_in(coef[256]), .rdup_out(a9_wr[1001]), .rdlo_out(a9_wr[1003]));
			radix2 #(.width(width)) rd_st8_1004  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1004]), .rdlo_in(a8_wr[1006]),  .coef_in(coef[0]), .rdup_out(a9_wr[1004]), .rdlo_out(a9_wr[1006]));
			radix2 #(.width(width)) rd_st8_1005  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1005]), .rdlo_in(a8_wr[1007]),  .coef_in(coef[256]), .rdup_out(a9_wr[1005]), .rdlo_out(a9_wr[1007]));
			radix2 #(.width(width)) rd_st8_1008  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1008]), .rdlo_in(a8_wr[1010]),  .coef_in(coef[0]), .rdup_out(a9_wr[1008]), .rdlo_out(a9_wr[1010]));
			radix2 #(.width(width)) rd_st8_1009  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1009]), .rdlo_in(a8_wr[1011]),  .coef_in(coef[256]), .rdup_out(a9_wr[1009]), .rdlo_out(a9_wr[1011]));
			radix2 #(.width(width)) rd_st8_1012  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1012]), .rdlo_in(a8_wr[1014]),  .coef_in(coef[0]), .rdup_out(a9_wr[1012]), .rdlo_out(a9_wr[1014]));
			radix2 #(.width(width)) rd_st8_1013  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1013]), .rdlo_in(a8_wr[1015]),  .coef_in(coef[256]), .rdup_out(a9_wr[1013]), .rdlo_out(a9_wr[1015]));
			radix2 #(.width(width)) rd_st8_1016  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1016]), .rdlo_in(a8_wr[1018]),  .coef_in(coef[0]), .rdup_out(a9_wr[1016]), .rdlo_out(a9_wr[1018]));
			radix2 #(.width(width)) rd_st8_1017  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1017]), .rdlo_in(a8_wr[1019]),  .coef_in(coef[256]), .rdup_out(a9_wr[1017]), .rdlo_out(a9_wr[1019]));
			radix2 #(.width(width)) rd_st8_1020  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1020]), .rdlo_in(a8_wr[1022]),  .coef_in(coef[0]), .rdup_out(a9_wr[1020]), .rdlo_out(a9_wr[1022]));
			radix2 #(.width(width)) rd_st8_1021  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1021]), .rdlo_in(a8_wr[1023]),  .coef_in(coef[256]), .rdup_out(a9_wr[1021]), .rdlo_out(a9_wr[1023]));

		//--- radix stage 9
			radix2 #(.width(width)) rd_st9_0   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[0]), .rdlo_in(a9_wr[1]),  .coef_in(coef[0]), .rdup_out(a10_wr[0]), .rdlo_out(a10_wr[1]));
			radix2 #(.width(width)) rd_st9_2   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[2]), .rdlo_in(a9_wr[3]),  .coef_in(coef[0]), .rdup_out(a10_wr[2]), .rdlo_out(a10_wr[3]));
			radix2 #(.width(width)) rd_st9_4   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[4]), .rdlo_in(a9_wr[5]),  .coef_in(coef[0]), .rdup_out(a10_wr[4]), .rdlo_out(a10_wr[5]));
			radix2 #(.width(width)) rd_st9_6   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[6]), .rdlo_in(a9_wr[7]),  .coef_in(coef[0]), .rdup_out(a10_wr[6]), .rdlo_out(a10_wr[7]));
			radix2 #(.width(width)) rd_st9_8   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[8]), .rdlo_in(a9_wr[9]),  .coef_in(coef[0]), .rdup_out(a10_wr[8]), .rdlo_out(a10_wr[9]));
			radix2 #(.width(width)) rd_st9_10  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[10]), .rdlo_in(a9_wr[11]),  .coef_in(coef[0]), .rdup_out(a10_wr[10]), .rdlo_out(a10_wr[11]));
			radix2 #(.width(width)) rd_st9_12  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[12]), .rdlo_in(a9_wr[13]),  .coef_in(coef[0]), .rdup_out(a10_wr[12]), .rdlo_out(a10_wr[13]));
			radix2 #(.width(width)) rd_st9_14  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[14]), .rdlo_in(a9_wr[15]),  .coef_in(coef[0]), .rdup_out(a10_wr[14]), .rdlo_out(a10_wr[15]));
			radix2 #(.width(width)) rd_st9_16  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[16]), .rdlo_in(a9_wr[17]),  .coef_in(coef[0]), .rdup_out(a10_wr[16]), .rdlo_out(a10_wr[17]));
			radix2 #(.width(width)) rd_st9_18  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[18]), .rdlo_in(a9_wr[19]),  .coef_in(coef[0]), .rdup_out(a10_wr[18]), .rdlo_out(a10_wr[19]));
			radix2 #(.width(width)) rd_st9_20  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[20]), .rdlo_in(a9_wr[21]),  .coef_in(coef[0]), .rdup_out(a10_wr[20]), .rdlo_out(a10_wr[21]));
			radix2 #(.width(width)) rd_st9_22  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[22]), .rdlo_in(a9_wr[23]),  .coef_in(coef[0]), .rdup_out(a10_wr[22]), .rdlo_out(a10_wr[23]));
			radix2 #(.width(width)) rd_st9_24  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[24]), .rdlo_in(a9_wr[25]),  .coef_in(coef[0]), .rdup_out(a10_wr[24]), .rdlo_out(a10_wr[25]));
			radix2 #(.width(width)) rd_st9_26  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[26]), .rdlo_in(a9_wr[27]),  .coef_in(coef[0]), .rdup_out(a10_wr[26]), .rdlo_out(a10_wr[27]));
			radix2 #(.width(width)) rd_st9_28  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[28]), .rdlo_in(a9_wr[29]),  .coef_in(coef[0]), .rdup_out(a10_wr[28]), .rdlo_out(a10_wr[29]));
			radix2 #(.width(width)) rd_st9_30  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[30]), .rdlo_in(a9_wr[31]),  .coef_in(coef[0]), .rdup_out(a10_wr[30]), .rdlo_out(a10_wr[31]));
			radix2 #(.width(width)) rd_st9_32  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[32]), .rdlo_in(a9_wr[33]),  .coef_in(coef[0]), .rdup_out(a10_wr[32]), .rdlo_out(a10_wr[33]));
			radix2 #(.width(width)) rd_st9_34  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[34]), .rdlo_in(a9_wr[35]),  .coef_in(coef[0]), .rdup_out(a10_wr[34]), .rdlo_out(a10_wr[35]));
			radix2 #(.width(width)) rd_st9_36  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[36]), .rdlo_in(a9_wr[37]),  .coef_in(coef[0]), .rdup_out(a10_wr[36]), .rdlo_out(a10_wr[37]));
			radix2 #(.width(width)) rd_st9_38  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[38]), .rdlo_in(a9_wr[39]),  .coef_in(coef[0]), .rdup_out(a10_wr[38]), .rdlo_out(a10_wr[39]));
			radix2 #(.width(width)) rd_st9_40  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[40]), .rdlo_in(a9_wr[41]),  .coef_in(coef[0]), .rdup_out(a10_wr[40]), .rdlo_out(a10_wr[41]));
			radix2 #(.width(width)) rd_st9_42  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[42]), .rdlo_in(a9_wr[43]),  .coef_in(coef[0]), .rdup_out(a10_wr[42]), .rdlo_out(a10_wr[43]));
			radix2 #(.width(width)) rd_st9_44  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[44]), .rdlo_in(a9_wr[45]),  .coef_in(coef[0]), .rdup_out(a10_wr[44]), .rdlo_out(a10_wr[45]));
			radix2 #(.width(width)) rd_st9_46  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[46]), .rdlo_in(a9_wr[47]),  .coef_in(coef[0]), .rdup_out(a10_wr[46]), .rdlo_out(a10_wr[47]));
			radix2 #(.width(width)) rd_st9_48  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[48]), .rdlo_in(a9_wr[49]),  .coef_in(coef[0]), .rdup_out(a10_wr[48]), .rdlo_out(a10_wr[49]));
			radix2 #(.width(width)) rd_st9_50  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[50]), .rdlo_in(a9_wr[51]),  .coef_in(coef[0]), .rdup_out(a10_wr[50]), .rdlo_out(a10_wr[51]));
			radix2 #(.width(width)) rd_st9_52  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[52]), .rdlo_in(a9_wr[53]),  .coef_in(coef[0]), .rdup_out(a10_wr[52]), .rdlo_out(a10_wr[53]));
			radix2 #(.width(width)) rd_st9_54  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[54]), .rdlo_in(a9_wr[55]),  .coef_in(coef[0]), .rdup_out(a10_wr[54]), .rdlo_out(a10_wr[55]));
			radix2 #(.width(width)) rd_st9_56  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[56]), .rdlo_in(a9_wr[57]),  .coef_in(coef[0]), .rdup_out(a10_wr[56]), .rdlo_out(a10_wr[57]));
			radix2 #(.width(width)) rd_st9_58  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[58]), .rdlo_in(a9_wr[59]),  .coef_in(coef[0]), .rdup_out(a10_wr[58]), .rdlo_out(a10_wr[59]));
			radix2 #(.width(width)) rd_st9_60  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[60]), .rdlo_in(a9_wr[61]),  .coef_in(coef[0]), .rdup_out(a10_wr[60]), .rdlo_out(a10_wr[61]));
			radix2 #(.width(width)) rd_st9_62  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[62]), .rdlo_in(a9_wr[63]),  .coef_in(coef[0]), .rdup_out(a10_wr[62]), .rdlo_out(a10_wr[63]));
			radix2 #(.width(width)) rd_st9_64  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[64]), .rdlo_in(a9_wr[65]),  .coef_in(coef[0]), .rdup_out(a10_wr[64]), .rdlo_out(a10_wr[65]));
			radix2 #(.width(width)) rd_st9_66  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[66]), .rdlo_in(a9_wr[67]),  .coef_in(coef[0]), .rdup_out(a10_wr[66]), .rdlo_out(a10_wr[67]));
			radix2 #(.width(width)) rd_st9_68  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[68]), .rdlo_in(a9_wr[69]),  .coef_in(coef[0]), .rdup_out(a10_wr[68]), .rdlo_out(a10_wr[69]));
			radix2 #(.width(width)) rd_st9_70  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[70]), .rdlo_in(a9_wr[71]),  .coef_in(coef[0]), .rdup_out(a10_wr[70]), .rdlo_out(a10_wr[71]));
			radix2 #(.width(width)) rd_st9_72  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[72]), .rdlo_in(a9_wr[73]),  .coef_in(coef[0]), .rdup_out(a10_wr[72]), .rdlo_out(a10_wr[73]));
			radix2 #(.width(width)) rd_st9_74  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[74]), .rdlo_in(a9_wr[75]),  .coef_in(coef[0]), .rdup_out(a10_wr[74]), .rdlo_out(a10_wr[75]));
			radix2 #(.width(width)) rd_st9_76  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[76]), .rdlo_in(a9_wr[77]),  .coef_in(coef[0]), .rdup_out(a10_wr[76]), .rdlo_out(a10_wr[77]));
			radix2 #(.width(width)) rd_st9_78  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[78]), .rdlo_in(a9_wr[79]),  .coef_in(coef[0]), .rdup_out(a10_wr[78]), .rdlo_out(a10_wr[79]));
			radix2 #(.width(width)) rd_st9_80  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[80]), .rdlo_in(a9_wr[81]),  .coef_in(coef[0]), .rdup_out(a10_wr[80]), .rdlo_out(a10_wr[81]));
			radix2 #(.width(width)) rd_st9_82  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[82]), .rdlo_in(a9_wr[83]),  .coef_in(coef[0]), .rdup_out(a10_wr[82]), .rdlo_out(a10_wr[83]));
			radix2 #(.width(width)) rd_st9_84  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[84]), .rdlo_in(a9_wr[85]),  .coef_in(coef[0]), .rdup_out(a10_wr[84]), .rdlo_out(a10_wr[85]));
			radix2 #(.width(width)) rd_st9_86  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[86]), .rdlo_in(a9_wr[87]),  .coef_in(coef[0]), .rdup_out(a10_wr[86]), .rdlo_out(a10_wr[87]));
			radix2 #(.width(width)) rd_st9_88  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[88]), .rdlo_in(a9_wr[89]),  .coef_in(coef[0]), .rdup_out(a10_wr[88]), .rdlo_out(a10_wr[89]));
			radix2 #(.width(width)) rd_st9_90  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[90]), .rdlo_in(a9_wr[91]),  .coef_in(coef[0]), .rdup_out(a10_wr[90]), .rdlo_out(a10_wr[91]));
			radix2 #(.width(width)) rd_st9_92  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[92]), .rdlo_in(a9_wr[93]),  .coef_in(coef[0]), .rdup_out(a10_wr[92]), .rdlo_out(a10_wr[93]));
			radix2 #(.width(width)) rd_st9_94  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[94]), .rdlo_in(a9_wr[95]),  .coef_in(coef[0]), .rdup_out(a10_wr[94]), .rdlo_out(a10_wr[95]));
			radix2 #(.width(width)) rd_st9_96  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[96]), .rdlo_in(a9_wr[97]),  .coef_in(coef[0]), .rdup_out(a10_wr[96]), .rdlo_out(a10_wr[97]));
			radix2 #(.width(width)) rd_st9_98  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[98]), .rdlo_in(a9_wr[99]),  .coef_in(coef[0]), .rdup_out(a10_wr[98]), .rdlo_out(a10_wr[99]));
			radix2 #(.width(width)) rd_st9_100  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[100]), .rdlo_in(a9_wr[101]),  .coef_in(coef[0]), .rdup_out(a10_wr[100]), .rdlo_out(a10_wr[101]));
			radix2 #(.width(width)) rd_st9_102  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[102]), .rdlo_in(a9_wr[103]),  .coef_in(coef[0]), .rdup_out(a10_wr[102]), .rdlo_out(a10_wr[103]));
			radix2 #(.width(width)) rd_st9_104  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[104]), .rdlo_in(a9_wr[105]),  .coef_in(coef[0]), .rdup_out(a10_wr[104]), .rdlo_out(a10_wr[105]));
			radix2 #(.width(width)) rd_st9_106  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[106]), .rdlo_in(a9_wr[107]),  .coef_in(coef[0]), .rdup_out(a10_wr[106]), .rdlo_out(a10_wr[107]));
			radix2 #(.width(width)) rd_st9_108  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[108]), .rdlo_in(a9_wr[109]),  .coef_in(coef[0]), .rdup_out(a10_wr[108]), .rdlo_out(a10_wr[109]));
			radix2 #(.width(width)) rd_st9_110  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[110]), .rdlo_in(a9_wr[111]),  .coef_in(coef[0]), .rdup_out(a10_wr[110]), .rdlo_out(a10_wr[111]));
			radix2 #(.width(width)) rd_st9_112  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[112]), .rdlo_in(a9_wr[113]),  .coef_in(coef[0]), .rdup_out(a10_wr[112]), .rdlo_out(a10_wr[113]));
			radix2 #(.width(width)) rd_st9_114  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[114]), .rdlo_in(a9_wr[115]),  .coef_in(coef[0]), .rdup_out(a10_wr[114]), .rdlo_out(a10_wr[115]));
			radix2 #(.width(width)) rd_st9_116  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[116]), .rdlo_in(a9_wr[117]),  .coef_in(coef[0]), .rdup_out(a10_wr[116]), .rdlo_out(a10_wr[117]));
			radix2 #(.width(width)) rd_st9_118  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[118]), .rdlo_in(a9_wr[119]),  .coef_in(coef[0]), .rdup_out(a10_wr[118]), .rdlo_out(a10_wr[119]));
			radix2 #(.width(width)) rd_st9_120  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[120]), .rdlo_in(a9_wr[121]),  .coef_in(coef[0]), .rdup_out(a10_wr[120]), .rdlo_out(a10_wr[121]));
			radix2 #(.width(width)) rd_st9_122  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[122]), .rdlo_in(a9_wr[123]),  .coef_in(coef[0]), .rdup_out(a10_wr[122]), .rdlo_out(a10_wr[123]));
			radix2 #(.width(width)) rd_st9_124  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[124]), .rdlo_in(a9_wr[125]),  .coef_in(coef[0]), .rdup_out(a10_wr[124]), .rdlo_out(a10_wr[125]));
			radix2 #(.width(width)) rd_st9_126  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[126]), .rdlo_in(a9_wr[127]),  .coef_in(coef[0]), .rdup_out(a10_wr[126]), .rdlo_out(a10_wr[127]));
			radix2 #(.width(width)) rd_st9_128  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[128]), .rdlo_in(a9_wr[129]),  .coef_in(coef[0]), .rdup_out(a10_wr[128]), .rdlo_out(a10_wr[129]));
			radix2 #(.width(width)) rd_st9_130  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[130]), .rdlo_in(a9_wr[131]),  .coef_in(coef[0]), .rdup_out(a10_wr[130]), .rdlo_out(a10_wr[131]));
			radix2 #(.width(width)) rd_st9_132  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[132]), .rdlo_in(a9_wr[133]),  .coef_in(coef[0]), .rdup_out(a10_wr[132]), .rdlo_out(a10_wr[133]));
			radix2 #(.width(width)) rd_st9_134  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[134]), .rdlo_in(a9_wr[135]),  .coef_in(coef[0]), .rdup_out(a10_wr[134]), .rdlo_out(a10_wr[135]));
			radix2 #(.width(width)) rd_st9_136  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[136]), .rdlo_in(a9_wr[137]),  .coef_in(coef[0]), .rdup_out(a10_wr[136]), .rdlo_out(a10_wr[137]));
			radix2 #(.width(width)) rd_st9_138  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[138]), .rdlo_in(a9_wr[139]),  .coef_in(coef[0]), .rdup_out(a10_wr[138]), .rdlo_out(a10_wr[139]));
			radix2 #(.width(width)) rd_st9_140  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[140]), .rdlo_in(a9_wr[141]),  .coef_in(coef[0]), .rdup_out(a10_wr[140]), .rdlo_out(a10_wr[141]));
			radix2 #(.width(width)) rd_st9_142  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[142]), .rdlo_in(a9_wr[143]),  .coef_in(coef[0]), .rdup_out(a10_wr[142]), .rdlo_out(a10_wr[143]));
			radix2 #(.width(width)) rd_st9_144  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[144]), .rdlo_in(a9_wr[145]),  .coef_in(coef[0]), .rdup_out(a10_wr[144]), .rdlo_out(a10_wr[145]));
			radix2 #(.width(width)) rd_st9_146  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[146]), .rdlo_in(a9_wr[147]),  .coef_in(coef[0]), .rdup_out(a10_wr[146]), .rdlo_out(a10_wr[147]));
			radix2 #(.width(width)) rd_st9_148  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[148]), .rdlo_in(a9_wr[149]),  .coef_in(coef[0]), .rdup_out(a10_wr[148]), .rdlo_out(a10_wr[149]));
			radix2 #(.width(width)) rd_st9_150  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[150]), .rdlo_in(a9_wr[151]),  .coef_in(coef[0]), .rdup_out(a10_wr[150]), .rdlo_out(a10_wr[151]));
			radix2 #(.width(width)) rd_st9_152  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[152]), .rdlo_in(a9_wr[153]),  .coef_in(coef[0]), .rdup_out(a10_wr[152]), .rdlo_out(a10_wr[153]));
			radix2 #(.width(width)) rd_st9_154  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[154]), .rdlo_in(a9_wr[155]),  .coef_in(coef[0]), .rdup_out(a10_wr[154]), .rdlo_out(a10_wr[155]));
			radix2 #(.width(width)) rd_st9_156  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[156]), .rdlo_in(a9_wr[157]),  .coef_in(coef[0]), .rdup_out(a10_wr[156]), .rdlo_out(a10_wr[157]));
			radix2 #(.width(width)) rd_st9_158  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[158]), .rdlo_in(a9_wr[159]),  .coef_in(coef[0]), .rdup_out(a10_wr[158]), .rdlo_out(a10_wr[159]));
			radix2 #(.width(width)) rd_st9_160  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[160]), .rdlo_in(a9_wr[161]),  .coef_in(coef[0]), .rdup_out(a10_wr[160]), .rdlo_out(a10_wr[161]));
			radix2 #(.width(width)) rd_st9_162  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[162]), .rdlo_in(a9_wr[163]),  .coef_in(coef[0]), .rdup_out(a10_wr[162]), .rdlo_out(a10_wr[163]));
			radix2 #(.width(width)) rd_st9_164  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[164]), .rdlo_in(a9_wr[165]),  .coef_in(coef[0]), .rdup_out(a10_wr[164]), .rdlo_out(a10_wr[165]));
			radix2 #(.width(width)) rd_st9_166  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[166]), .rdlo_in(a9_wr[167]),  .coef_in(coef[0]), .rdup_out(a10_wr[166]), .rdlo_out(a10_wr[167]));
			radix2 #(.width(width)) rd_st9_168  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[168]), .rdlo_in(a9_wr[169]),  .coef_in(coef[0]), .rdup_out(a10_wr[168]), .rdlo_out(a10_wr[169]));
			radix2 #(.width(width)) rd_st9_170  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[170]), .rdlo_in(a9_wr[171]),  .coef_in(coef[0]), .rdup_out(a10_wr[170]), .rdlo_out(a10_wr[171]));
			radix2 #(.width(width)) rd_st9_172  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[172]), .rdlo_in(a9_wr[173]),  .coef_in(coef[0]), .rdup_out(a10_wr[172]), .rdlo_out(a10_wr[173]));
			radix2 #(.width(width)) rd_st9_174  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[174]), .rdlo_in(a9_wr[175]),  .coef_in(coef[0]), .rdup_out(a10_wr[174]), .rdlo_out(a10_wr[175]));
			radix2 #(.width(width)) rd_st9_176  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[176]), .rdlo_in(a9_wr[177]),  .coef_in(coef[0]), .rdup_out(a10_wr[176]), .rdlo_out(a10_wr[177]));
			radix2 #(.width(width)) rd_st9_178  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[178]), .rdlo_in(a9_wr[179]),  .coef_in(coef[0]), .rdup_out(a10_wr[178]), .rdlo_out(a10_wr[179]));
			radix2 #(.width(width)) rd_st9_180  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[180]), .rdlo_in(a9_wr[181]),  .coef_in(coef[0]), .rdup_out(a10_wr[180]), .rdlo_out(a10_wr[181]));
			radix2 #(.width(width)) rd_st9_182  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[182]), .rdlo_in(a9_wr[183]),  .coef_in(coef[0]), .rdup_out(a10_wr[182]), .rdlo_out(a10_wr[183]));
			radix2 #(.width(width)) rd_st9_184  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[184]), .rdlo_in(a9_wr[185]),  .coef_in(coef[0]), .rdup_out(a10_wr[184]), .rdlo_out(a10_wr[185]));
			radix2 #(.width(width)) rd_st9_186  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[186]), .rdlo_in(a9_wr[187]),  .coef_in(coef[0]), .rdup_out(a10_wr[186]), .rdlo_out(a10_wr[187]));
			radix2 #(.width(width)) rd_st9_188  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[188]), .rdlo_in(a9_wr[189]),  .coef_in(coef[0]), .rdup_out(a10_wr[188]), .rdlo_out(a10_wr[189]));
			radix2 #(.width(width)) rd_st9_190  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[190]), .rdlo_in(a9_wr[191]),  .coef_in(coef[0]), .rdup_out(a10_wr[190]), .rdlo_out(a10_wr[191]));
			radix2 #(.width(width)) rd_st9_192  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[192]), .rdlo_in(a9_wr[193]),  .coef_in(coef[0]), .rdup_out(a10_wr[192]), .rdlo_out(a10_wr[193]));
			radix2 #(.width(width)) rd_st9_194  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[194]), .rdlo_in(a9_wr[195]),  .coef_in(coef[0]), .rdup_out(a10_wr[194]), .rdlo_out(a10_wr[195]));
			radix2 #(.width(width)) rd_st9_196  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[196]), .rdlo_in(a9_wr[197]),  .coef_in(coef[0]), .rdup_out(a10_wr[196]), .rdlo_out(a10_wr[197]));
			radix2 #(.width(width)) rd_st9_198  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[198]), .rdlo_in(a9_wr[199]),  .coef_in(coef[0]), .rdup_out(a10_wr[198]), .rdlo_out(a10_wr[199]));
			radix2 #(.width(width)) rd_st9_200  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[200]), .rdlo_in(a9_wr[201]),  .coef_in(coef[0]), .rdup_out(a10_wr[200]), .rdlo_out(a10_wr[201]));
			radix2 #(.width(width)) rd_st9_202  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[202]), .rdlo_in(a9_wr[203]),  .coef_in(coef[0]), .rdup_out(a10_wr[202]), .rdlo_out(a10_wr[203]));
			radix2 #(.width(width)) rd_st9_204  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[204]), .rdlo_in(a9_wr[205]),  .coef_in(coef[0]), .rdup_out(a10_wr[204]), .rdlo_out(a10_wr[205]));
			radix2 #(.width(width)) rd_st9_206  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[206]), .rdlo_in(a9_wr[207]),  .coef_in(coef[0]), .rdup_out(a10_wr[206]), .rdlo_out(a10_wr[207]));
			radix2 #(.width(width)) rd_st9_208  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[208]), .rdlo_in(a9_wr[209]),  .coef_in(coef[0]), .rdup_out(a10_wr[208]), .rdlo_out(a10_wr[209]));
			radix2 #(.width(width)) rd_st9_210  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[210]), .rdlo_in(a9_wr[211]),  .coef_in(coef[0]), .rdup_out(a10_wr[210]), .rdlo_out(a10_wr[211]));
			radix2 #(.width(width)) rd_st9_212  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[212]), .rdlo_in(a9_wr[213]),  .coef_in(coef[0]), .rdup_out(a10_wr[212]), .rdlo_out(a10_wr[213]));
			radix2 #(.width(width)) rd_st9_214  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[214]), .rdlo_in(a9_wr[215]),  .coef_in(coef[0]), .rdup_out(a10_wr[214]), .rdlo_out(a10_wr[215]));
			radix2 #(.width(width)) rd_st9_216  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[216]), .rdlo_in(a9_wr[217]),  .coef_in(coef[0]), .rdup_out(a10_wr[216]), .rdlo_out(a10_wr[217]));
			radix2 #(.width(width)) rd_st9_218  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[218]), .rdlo_in(a9_wr[219]),  .coef_in(coef[0]), .rdup_out(a10_wr[218]), .rdlo_out(a10_wr[219]));
			radix2 #(.width(width)) rd_st9_220  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[220]), .rdlo_in(a9_wr[221]),  .coef_in(coef[0]), .rdup_out(a10_wr[220]), .rdlo_out(a10_wr[221]));
			radix2 #(.width(width)) rd_st9_222  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[222]), .rdlo_in(a9_wr[223]),  .coef_in(coef[0]), .rdup_out(a10_wr[222]), .rdlo_out(a10_wr[223]));
			radix2 #(.width(width)) rd_st9_224  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[224]), .rdlo_in(a9_wr[225]),  .coef_in(coef[0]), .rdup_out(a10_wr[224]), .rdlo_out(a10_wr[225]));
			radix2 #(.width(width)) rd_st9_226  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[226]), .rdlo_in(a9_wr[227]),  .coef_in(coef[0]), .rdup_out(a10_wr[226]), .rdlo_out(a10_wr[227]));
			radix2 #(.width(width)) rd_st9_228  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[228]), .rdlo_in(a9_wr[229]),  .coef_in(coef[0]), .rdup_out(a10_wr[228]), .rdlo_out(a10_wr[229]));
			radix2 #(.width(width)) rd_st9_230  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[230]), .rdlo_in(a9_wr[231]),  .coef_in(coef[0]), .rdup_out(a10_wr[230]), .rdlo_out(a10_wr[231]));
			radix2 #(.width(width)) rd_st9_232  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[232]), .rdlo_in(a9_wr[233]),  .coef_in(coef[0]), .rdup_out(a10_wr[232]), .rdlo_out(a10_wr[233]));
			radix2 #(.width(width)) rd_st9_234  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[234]), .rdlo_in(a9_wr[235]),  .coef_in(coef[0]), .rdup_out(a10_wr[234]), .rdlo_out(a10_wr[235]));
			radix2 #(.width(width)) rd_st9_236  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[236]), .rdlo_in(a9_wr[237]),  .coef_in(coef[0]), .rdup_out(a10_wr[236]), .rdlo_out(a10_wr[237]));
			radix2 #(.width(width)) rd_st9_238  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[238]), .rdlo_in(a9_wr[239]),  .coef_in(coef[0]), .rdup_out(a10_wr[238]), .rdlo_out(a10_wr[239]));
			radix2 #(.width(width)) rd_st9_240  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[240]), .rdlo_in(a9_wr[241]),  .coef_in(coef[0]), .rdup_out(a10_wr[240]), .rdlo_out(a10_wr[241]));
			radix2 #(.width(width)) rd_st9_242  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[242]), .rdlo_in(a9_wr[243]),  .coef_in(coef[0]), .rdup_out(a10_wr[242]), .rdlo_out(a10_wr[243]));
			radix2 #(.width(width)) rd_st9_244  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[244]), .rdlo_in(a9_wr[245]),  .coef_in(coef[0]), .rdup_out(a10_wr[244]), .rdlo_out(a10_wr[245]));
			radix2 #(.width(width)) rd_st9_246  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[246]), .rdlo_in(a9_wr[247]),  .coef_in(coef[0]), .rdup_out(a10_wr[246]), .rdlo_out(a10_wr[247]));
			radix2 #(.width(width)) rd_st9_248  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[248]), .rdlo_in(a9_wr[249]),  .coef_in(coef[0]), .rdup_out(a10_wr[248]), .rdlo_out(a10_wr[249]));
			radix2 #(.width(width)) rd_st9_250  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[250]), .rdlo_in(a9_wr[251]),  .coef_in(coef[0]), .rdup_out(a10_wr[250]), .rdlo_out(a10_wr[251]));
			radix2 #(.width(width)) rd_st9_252  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[252]), .rdlo_in(a9_wr[253]),  .coef_in(coef[0]), .rdup_out(a10_wr[252]), .rdlo_out(a10_wr[253]));
			radix2 #(.width(width)) rd_st9_254  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[254]), .rdlo_in(a9_wr[255]),  .coef_in(coef[0]), .rdup_out(a10_wr[254]), .rdlo_out(a10_wr[255]));
			radix2 #(.width(width)) rd_st9_256  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[256]), .rdlo_in(a9_wr[257]),  .coef_in(coef[0]), .rdup_out(a10_wr[256]), .rdlo_out(a10_wr[257]));
			radix2 #(.width(width)) rd_st9_258  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[258]), .rdlo_in(a9_wr[259]),  .coef_in(coef[0]), .rdup_out(a10_wr[258]), .rdlo_out(a10_wr[259]));
			radix2 #(.width(width)) rd_st9_260  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[260]), .rdlo_in(a9_wr[261]),  .coef_in(coef[0]), .rdup_out(a10_wr[260]), .rdlo_out(a10_wr[261]));
			radix2 #(.width(width)) rd_st9_262  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[262]), .rdlo_in(a9_wr[263]),  .coef_in(coef[0]), .rdup_out(a10_wr[262]), .rdlo_out(a10_wr[263]));
			radix2 #(.width(width)) rd_st9_264  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[264]), .rdlo_in(a9_wr[265]),  .coef_in(coef[0]), .rdup_out(a10_wr[264]), .rdlo_out(a10_wr[265]));
			radix2 #(.width(width)) rd_st9_266  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[266]), .rdlo_in(a9_wr[267]),  .coef_in(coef[0]), .rdup_out(a10_wr[266]), .rdlo_out(a10_wr[267]));
			radix2 #(.width(width)) rd_st9_268  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[268]), .rdlo_in(a9_wr[269]),  .coef_in(coef[0]), .rdup_out(a10_wr[268]), .rdlo_out(a10_wr[269]));
			radix2 #(.width(width)) rd_st9_270  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[270]), .rdlo_in(a9_wr[271]),  .coef_in(coef[0]), .rdup_out(a10_wr[270]), .rdlo_out(a10_wr[271]));
			radix2 #(.width(width)) rd_st9_272  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[272]), .rdlo_in(a9_wr[273]),  .coef_in(coef[0]), .rdup_out(a10_wr[272]), .rdlo_out(a10_wr[273]));
			radix2 #(.width(width)) rd_st9_274  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[274]), .rdlo_in(a9_wr[275]),  .coef_in(coef[0]), .rdup_out(a10_wr[274]), .rdlo_out(a10_wr[275]));
			radix2 #(.width(width)) rd_st9_276  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[276]), .rdlo_in(a9_wr[277]),  .coef_in(coef[0]), .rdup_out(a10_wr[276]), .rdlo_out(a10_wr[277]));
			radix2 #(.width(width)) rd_st9_278  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[278]), .rdlo_in(a9_wr[279]),  .coef_in(coef[0]), .rdup_out(a10_wr[278]), .rdlo_out(a10_wr[279]));
			radix2 #(.width(width)) rd_st9_280  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[280]), .rdlo_in(a9_wr[281]),  .coef_in(coef[0]), .rdup_out(a10_wr[280]), .rdlo_out(a10_wr[281]));
			radix2 #(.width(width)) rd_st9_282  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[282]), .rdlo_in(a9_wr[283]),  .coef_in(coef[0]), .rdup_out(a10_wr[282]), .rdlo_out(a10_wr[283]));
			radix2 #(.width(width)) rd_st9_284  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[284]), .rdlo_in(a9_wr[285]),  .coef_in(coef[0]), .rdup_out(a10_wr[284]), .rdlo_out(a10_wr[285]));
			radix2 #(.width(width)) rd_st9_286  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[286]), .rdlo_in(a9_wr[287]),  .coef_in(coef[0]), .rdup_out(a10_wr[286]), .rdlo_out(a10_wr[287]));
			radix2 #(.width(width)) rd_st9_288  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[288]), .rdlo_in(a9_wr[289]),  .coef_in(coef[0]), .rdup_out(a10_wr[288]), .rdlo_out(a10_wr[289]));
			radix2 #(.width(width)) rd_st9_290  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[290]), .rdlo_in(a9_wr[291]),  .coef_in(coef[0]), .rdup_out(a10_wr[290]), .rdlo_out(a10_wr[291]));
			radix2 #(.width(width)) rd_st9_292  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[292]), .rdlo_in(a9_wr[293]),  .coef_in(coef[0]), .rdup_out(a10_wr[292]), .rdlo_out(a10_wr[293]));
			radix2 #(.width(width)) rd_st9_294  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[294]), .rdlo_in(a9_wr[295]),  .coef_in(coef[0]), .rdup_out(a10_wr[294]), .rdlo_out(a10_wr[295]));
			radix2 #(.width(width)) rd_st9_296  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[296]), .rdlo_in(a9_wr[297]),  .coef_in(coef[0]), .rdup_out(a10_wr[296]), .rdlo_out(a10_wr[297]));
			radix2 #(.width(width)) rd_st9_298  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[298]), .rdlo_in(a9_wr[299]),  .coef_in(coef[0]), .rdup_out(a10_wr[298]), .rdlo_out(a10_wr[299]));
			radix2 #(.width(width)) rd_st9_300  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[300]), .rdlo_in(a9_wr[301]),  .coef_in(coef[0]), .rdup_out(a10_wr[300]), .rdlo_out(a10_wr[301]));
			radix2 #(.width(width)) rd_st9_302  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[302]), .rdlo_in(a9_wr[303]),  .coef_in(coef[0]), .rdup_out(a10_wr[302]), .rdlo_out(a10_wr[303]));
			radix2 #(.width(width)) rd_st9_304  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[304]), .rdlo_in(a9_wr[305]),  .coef_in(coef[0]), .rdup_out(a10_wr[304]), .rdlo_out(a10_wr[305]));
			radix2 #(.width(width)) rd_st9_306  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[306]), .rdlo_in(a9_wr[307]),  .coef_in(coef[0]), .rdup_out(a10_wr[306]), .rdlo_out(a10_wr[307]));
			radix2 #(.width(width)) rd_st9_308  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[308]), .rdlo_in(a9_wr[309]),  .coef_in(coef[0]), .rdup_out(a10_wr[308]), .rdlo_out(a10_wr[309]));
			radix2 #(.width(width)) rd_st9_310  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[310]), .rdlo_in(a9_wr[311]),  .coef_in(coef[0]), .rdup_out(a10_wr[310]), .rdlo_out(a10_wr[311]));
			radix2 #(.width(width)) rd_st9_312  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[312]), .rdlo_in(a9_wr[313]),  .coef_in(coef[0]), .rdup_out(a10_wr[312]), .rdlo_out(a10_wr[313]));
			radix2 #(.width(width)) rd_st9_314  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[314]), .rdlo_in(a9_wr[315]),  .coef_in(coef[0]), .rdup_out(a10_wr[314]), .rdlo_out(a10_wr[315]));
			radix2 #(.width(width)) rd_st9_316  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[316]), .rdlo_in(a9_wr[317]),  .coef_in(coef[0]), .rdup_out(a10_wr[316]), .rdlo_out(a10_wr[317]));
			radix2 #(.width(width)) rd_st9_318  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[318]), .rdlo_in(a9_wr[319]),  .coef_in(coef[0]), .rdup_out(a10_wr[318]), .rdlo_out(a10_wr[319]));
			radix2 #(.width(width)) rd_st9_320  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[320]), .rdlo_in(a9_wr[321]),  .coef_in(coef[0]), .rdup_out(a10_wr[320]), .rdlo_out(a10_wr[321]));
			radix2 #(.width(width)) rd_st9_322  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[322]), .rdlo_in(a9_wr[323]),  .coef_in(coef[0]), .rdup_out(a10_wr[322]), .rdlo_out(a10_wr[323]));
			radix2 #(.width(width)) rd_st9_324  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[324]), .rdlo_in(a9_wr[325]),  .coef_in(coef[0]), .rdup_out(a10_wr[324]), .rdlo_out(a10_wr[325]));
			radix2 #(.width(width)) rd_st9_326  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[326]), .rdlo_in(a9_wr[327]),  .coef_in(coef[0]), .rdup_out(a10_wr[326]), .rdlo_out(a10_wr[327]));
			radix2 #(.width(width)) rd_st9_328  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[328]), .rdlo_in(a9_wr[329]),  .coef_in(coef[0]), .rdup_out(a10_wr[328]), .rdlo_out(a10_wr[329]));
			radix2 #(.width(width)) rd_st9_330  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[330]), .rdlo_in(a9_wr[331]),  .coef_in(coef[0]), .rdup_out(a10_wr[330]), .rdlo_out(a10_wr[331]));
			radix2 #(.width(width)) rd_st9_332  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[332]), .rdlo_in(a9_wr[333]),  .coef_in(coef[0]), .rdup_out(a10_wr[332]), .rdlo_out(a10_wr[333]));
			radix2 #(.width(width)) rd_st9_334  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[334]), .rdlo_in(a9_wr[335]),  .coef_in(coef[0]), .rdup_out(a10_wr[334]), .rdlo_out(a10_wr[335]));
			radix2 #(.width(width)) rd_st9_336  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[336]), .rdlo_in(a9_wr[337]),  .coef_in(coef[0]), .rdup_out(a10_wr[336]), .rdlo_out(a10_wr[337]));
			radix2 #(.width(width)) rd_st9_338  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[338]), .rdlo_in(a9_wr[339]),  .coef_in(coef[0]), .rdup_out(a10_wr[338]), .rdlo_out(a10_wr[339]));
			radix2 #(.width(width)) rd_st9_340  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[340]), .rdlo_in(a9_wr[341]),  .coef_in(coef[0]), .rdup_out(a10_wr[340]), .rdlo_out(a10_wr[341]));
			radix2 #(.width(width)) rd_st9_342  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[342]), .rdlo_in(a9_wr[343]),  .coef_in(coef[0]), .rdup_out(a10_wr[342]), .rdlo_out(a10_wr[343]));
			radix2 #(.width(width)) rd_st9_344  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[344]), .rdlo_in(a9_wr[345]),  .coef_in(coef[0]), .rdup_out(a10_wr[344]), .rdlo_out(a10_wr[345]));
			radix2 #(.width(width)) rd_st9_346  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[346]), .rdlo_in(a9_wr[347]),  .coef_in(coef[0]), .rdup_out(a10_wr[346]), .rdlo_out(a10_wr[347]));
			radix2 #(.width(width)) rd_st9_348  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[348]), .rdlo_in(a9_wr[349]),  .coef_in(coef[0]), .rdup_out(a10_wr[348]), .rdlo_out(a10_wr[349]));
			radix2 #(.width(width)) rd_st9_350  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[350]), .rdlo_in(a9_wr[351]),  .coef_in(coef[0]), .rdup_out(a10_wr[350]), .rdlo_out(a10_wr[351]));
			radix2 #(.width(width)) rd_st9_352  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[352]), .rdlo_in(a9_wr[353]),  .coef_in(coef[0]), .rdup_out(a10_wr[352]), .rdlo_out(a10_wr[353]));
			radix2 #(.width(width)) rd_st9_354  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[354]), .rdlo_in(a9_wr[355]),  .coef_in(coef[0]), .rdup_out(a10_wr[354]), .rdlo_out(a10_wr[355]));
			radix2 #(.width(width)) rd_st9_356  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[356]), .rdlo_in(a9_wr[357]),  .coef_in(coef[0]), .rdup_out(a10_wr[356]), .rdlo_out(a10_wr[357]));
			radix2 #(.width(width)) rd_st9_358  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[358]), .rdlo_in(a9_wr[359]),  .coef_in(coef[0]), .rdup_out(a10_wr[358]), .rdlo_out(a10_wr[359]));
			radix2 #(.width(width)) rd_st9_360  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[360]), .rdlo_in(a9_wr[361]),  .coef_in(coef[0]), .rdup_out(a10_wr[360]), .rdlo_out(a10_wr[361]));
			radix2 #(.width(width)) rd_st9_362  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[362]), .rdlo_in(a9_wr[363]),  .coef_in(coef[0]), .rdup_out(a10_wr[362]), .rdlo_out(a10_wr[363]));
			radix2 #(.width(width)) rd_st9_364  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[364]), .rdlo_in(a9_wr[365]),  .coef_in(coef[0]), .rdup_out(a10_wr[364]), .rdlo_out(a10_wr[365]));
			radix2 #(.width(width)) rd_st9_366  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[366]), .rdlo_in(a9_wr[367]),  .coef_in(coef[0]), .rdup_out(a10_wr[366]), .rdlo_out(a10_wr[367]));
			radix2 #(.width(width)) rd_st9_368  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[368]), .rdlo_in(a9_wr[369]),  .coef_in(coef[0]), .rdup_out(a10_wr[368]), .rdlo_out(a10_wr[369]));
			radix2 #(.width(width)) rd_st9_370  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[370]), .rdlo_in(a9_wr[371]),  .coef_in(coef[0]), .rdup_out(a10_wr[370]), .rdlo_out(a10_wr[371]));
			radix2 #(.width(width)) rd_st9_372  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[372]), .rdlo_in(a9_wr[373]),  .coef_in(coef[0]), .rdup_out(a10_wr[372]), .rdlo_out(a10_wr[373]));
			radix2 #(.width(width)) rd_st9_374  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[374]), .rdlo_in(a9_wr[375]),  .coef_in(coef[0]), .rdup_out(a10_wr[374]), .rdlo_out(a10_wr[375]));
			radix2 #(.width(width)) rd_st9_376  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[376]), .rdlo_in(a9_wr[377]),  .coef_in(coef[0]), .rdup_out(a10_wr[376]), .rdlo_out(a10_wr[377]));
			radix2 #(.width(width)) rd_st9_378  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[378]), .rdlo_in(a9_wr[379]),  .coef_in(coef[0]), .rdup_out(a10_wr[378]), .rdlo_out(a10_wr[379]));
			radix2 #(.width(width)) rd_st9_380  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[380]), .rdlo_in(a9_wr[381]),  .coef_in(coef[0]), .rdup_out(a10_wr[380]), .rdlo_out(a10_wr[381]));
			radix2 #(.width(width)) rd_st9_382  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[382]), .rdlo_in(a9_wr[383]),  .coef_in(coef[0]), .rdup_out(a10_wr[382]), .rdlo_out(a10_wr[383]));
			radix2 #(.width(width)) rd_st9_384  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[384]), .rdlo_in(a9_wr[385]),  .coef_in(coef[0]), .rdup_out(a10_wr[384]), .rdlo_out(a10_wr[385]));
			radix2 #(.width(width)) rd_st9_386  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[386]), .rdlo_in(a9_wr[387]),  .coef_in(coef[0]), .rdup_out(a10_wr[386]), .rdlo_out(a10_wr[387]));
			radix2 #(.width(width)) rd_st9_388  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[388]), .rdlo_in(a9_wr[389]),  .coef_in(coef[0]), .rdup_out(a10_wr[388]), .rdlo_out(a10_wr[389]));
			radix2 #(.width(width)) rd_st9_390  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[390]), .rdlo_in(a9_wr[391]),  .coef_in(coef[0]), .rdup_out(a10_wr[390]), .rdlo_out(a10_wr[391]));
			radix2 #(.width(width)) rd_st9_392  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[392]), .rdlo_in(a9_wr[393]),  .coef_in(coef[0]), .rdup_out(a10_wr[392]), .rdlo_out(a10_wr[393]));
			radix2 #(.width(width)) rd_st9_394  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[394]), .rdlo_in(a9_wr[395]),  .coef_in(coef[0]), .rdup_out(a10_wr[394]), .rdlo_out(a10_wr[395]));
			radix2 #(.width(width)) rd_st9_396  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[396]), .rdlo_in(a9_wr[397]),  .coef_in(coef[0]), .rdup_out(a10_wr[396]), .rdlo_out(a10_wr[397]));
			radix2 #(.width(width)) rd_st9_398  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[398]), .rdlo_in(a9_wr[399]),  .coef_in(coef[0]), .rdup_out(a10_wr[398]), .rdlo_out(a10_wr[399]));
			radix2 #(.width(width)) rd_st9_400  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[400]), .rdlo_in(a9_wr[401]),  .coef_in(coef[0]), .rdup_out(a10_wr[400]), .rdlo_out(a10_wr[401]));
			radix2 #(.width(width)) rd_st9_402  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[402]), .rdlo_in(a9_wr[403]),  .coef_in(coef[0]), .rdup_out(a10_wr[402]), .rdlo_out(a10_wr[403]));
			radix2 #(.width(width)) rd_st9_404  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[404]), .rdlo_in(a9_wr[405]),  .coef_in(coef[0]), .rdup_out(a10_wr[404]), .rdlo_out(a10_wr[405]));
			radix2 #(.width(width)) rd_st9_406  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[406]), .rdlo_in(a9_wr[407]),  .coef_in(coef[0]), .rdup_out(a10_wr[406]), .rdlo_out(a10_wr[407]));
			radix2 #(.width(width)) rd_st9_408  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[408]), .rdlo_in(a9_wr[409]),  .coef_in(coef[0]), .rdup_out(a10_wr[408]), .rdlo_out(a10_wr[409]));
			radix2 #(.width(width)) rd_st9_410  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[410]), .rdlo_in(a9_wr[411]),  .coef_in(coef[0]), .rdup_out(a10_wr[410]), .rdlo_out(a10_wr[411]));
			radix2 #(.width(width)) rd_st9_412  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[412]), .rdlo_in(a9_wr[413]),  .coef_in(coef[0]), .rdup_out(a10_wr[412]), .rdlo_out(a10_wr[413]));
			radix2 #(.width(width)) rd_st9_414  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[414]), .rdlo_in(a9_wr[415]),  .coef_in(coef[0]), .rdup_out(a10_wr[414]), .rdlo_out(a10_wr[415]));
			radix2 #(.width(width)) rd_st9_416  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[416]), .rdlo_in(a9_wr[417]),  .coef_in(coef[0]), .rdup_out(a10_wr[416]), .rdlo_out(a10_wr[417]));
			radix2 #(.width(width)) rd_st9_418  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[418]), .rdlo_in(a9_wr[419]),  .coef_in(coef[0]), .rdup_out(a10_wr[418]), .rdlo_out(a10_wr[419]));
			radix2 #(.width(width)) rd_st9_420  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[420]), .rdlo_in(a9_wr[421]),  .coef_in(coef[0]), .rdup_out(a10_wr[420]), .rdlo_out(a10_wr[421]));
			radix2 #(.width(width)) rd_st9_422  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[422]), .rdlo_in(a9_wr[423]),  .coef_in(coef[0]), .rdup_out(a10_wr[422]), .rdlo_out(a10_wr[423]));
			radix2 #(.width(width)) rd_st9_424  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[424]), .rdlo_in(a9_wr[425]),  .coef_in(coef[0]), .rdup_out(a10_wr[424]), .rdlo_out(a10_wr[425]));
			radix2 #(.width(width)) rd_st9_426  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[426]), .rdlo_in(a9_wr[427]),  .coef_in(coef[0]), .rdup_out(a10_wr[426]), .rdlo_out(a10_wr[427]));
			radix2 #(.width(width)) rd_st9_428  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[428]), .rdlo_in(a9_wr[429]),  .coef_in(coef[0]), .rdup_out(a10_wr[428]), .rdlo_out(a10_wr[429]));
			radix2 #(.width(width)) rd_st9_430  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[430]), .rdlo_in(a9_wr[431]),  .coef_in(coef[0]), .rdup_out(a10_wr[430]), .rdlo_out(a10_wr[431]));
			radix2 #(.width(width)) rd_st9_432  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[432]), .rdlo_in(a9_wr[433]),  .coef_in(coef[0]), .rdup_out(a10_wr[432]), .rdlo_out(a10_wr[433]));
			radix2 #(.width(width)) rd_st9_434  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[434]), .rdlo_in(a9_wr[435]),  .coef_in(coef[0]), .rdup_out(a10_wr[434]), .rdlo_out(a10_wr[435]));
			radix2 #(.width(width)) rd_st9_436  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[436]), .rdlo_in(a9_wr[437]),  .coef_in(coef[0]), .rdup_out(a10_wr[436]), .rdlo_out(a10_wr[437]));
			radix2 #(.width(width)) rd_st9_438  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[438]), .rdlo_in(a9_wr[439]),  .coef_in(coef[0]), .rdup_out(a10_wr[438]), .rdlo_out(a10_wr[439]));
			radix2 #(.width(width)) rd_st9_440  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[440]), .rdlo_in(a9_wr[441]),  .coef_in(coef[0]), .rdup_out(a10_wr[440]), .rdlo_out(a10_wr[441]));
			radix2 #(.width(width)) rd_st9_442  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[442]), .rdlo_in(a9_wr[443]),  .coef_in(coef[0]), .rdup_out(a10_wr[442]), .rdlo_out(a10_wr[443]));
			radix2 #(.width(width)) rd_st9_444  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[444]), .rdlo_in(a9_wr[445]),  .coef_in(coef[0]), .rdup_out(a10_wr[444]), .rdlo_out(a10_wr[445]));
			radix2 #(.width(width)) rd_st9_446  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[446]), .rdlo_in(a9_wr[447]),  .coef_in(coef[0]), .rdup_out(a10_wr[446]), .rdlo_out(a10_wr[447]));
			radix2 #(.width(width)) rd_st9_448  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[448]), .rdlo_in(a9_wr[449]),  .coef_in(coef[0]), .rdup_out(a10_wr[448]), .rdlo_out(a10_wr[449]));
			radix2 #(.width(width)) rd_st9_450  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[450]), .rdlo_in(a9_wr[451]),  .coef_in(coef[0]), .rdup_out(a10_wr[450]), .rdlo_out(a10_wr[451]));
			radix2 #(.width(width)) rd_st9_452  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[452]), .rdlo_in(a9_wr[453]),  .coef_in(coef[0]), .rdup_out(a10_wr[452]), .rdlo_out(a10_wr[453]));
			radix2 #(.width(width)) rd_st9_454  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[454]), .rdlo_in(a9_wr[455]),  .coef_in(coef[0]), .rdup_out(a10_wr[454]), .rdlo_out(a10_wr[455]));
			radix2 #(.width(width)) rd_st9_456  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[456]), .rdlo_in(a9_wr[457]),  .coef_in(coef[0]), .rdup_out(a10_wr[456]), .rdlo_out(a10_wr[457]));
			radix2 #(.width(width)) rd_st9_458  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[458]), .rdlo_in(a9_wr[459]),  .coef_in(coef[0]), .rdup_out(a10_wr[458]), .rdlo_out(a10_wr[459]));
			radix2 #(.width(width)) rd_st9_460  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[460]), .rdlo_in(a9_wr[461]),  .coef_in(coef[0]), .rdup_out(a10_wr[460]), .rdlo_out(a10_wr[461]));
			radix2 #(.width(width)) rd_st9_462  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[462]), .rdlo_in(a9_wr[463]),  .coef_in(coef[0]), .rdup_out(a10_wr[462]), .rdlo_out(a10_wr[463]));
			radix2 #(.width(width)) rd_st9_464  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[464]), .rdlo_in(a9_wr[465]),  .coef_in(coef[0]), .rdup_out(a10_wr[464]), .rdlo_out(a10_wr[465]));
			radix2 #(.width(width)) rd_st9_466  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[466]), .rdlo_in(a9_wr[467]),  .coef_in(coef[0]), .rdup_out(a10_wr[466]), .rdlo_out(a10_wr[467]));
			radix2 #(.width(width)) rd_st9_468  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[468]), .rdlo_in(a9_wr[469]),  .coef_in(coef[0]), .rdup_out(a10_wr[468]), .rdlo_out(a10_wr[469]));
			radix2 #(.width(width)) rd_st9_470  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[470]), .rdlo_in(a9_wr[471]),  .coef_in(coef[0]), .rdup_out(a10_wr[470]), .rdlo_out(a10_wr[471]));
			radix2 #(.width(width)) rd_st9_472  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[472]), .rdlo_in(a9_wr[473]),  .coef_in(coef[0]), .rdup_out(a10_wr[472]), .rdlo_out(a10_wr[473]));
			radix2 #(.width(width)) rd_st9_474  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[474]), .rdlo_in(a9_wr[475]),  .coef_in(coef[0]), .rdup_out(a10_wr[474]), .rdlo_out(a10_wr[475]));
			radix2 #(.width(width)) rd_st9_476  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[476]), .rdlo_in(a9_wr[477]),  .coef_in(coef[0]), .rdup_out(a10_wr[476]), .rdlo_out(a10_wr[477]));
			radix2 #(.width(width)) rd_st9_478  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[478]), .rdlo_in(a9_wr[479]),  .coef_in(coef[0]), .rdup_out(a10_wr[478]), .rdlo_out(a10_wr[479]));
			radix2 #(.width(width)) rd_st9_480  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[480]), .rdlo_in(a9_wr[481]),  .coef_in(coef[0]), .rdup_out(a10_wr[480]), .rdlo_out(a10_wr[481]));
			radix2 #(.width(width)) rd_st9_482  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[482]), .rdlo_in(a9_wr[483]),  .coef_in(coef[0]), .rdup_out(a10_wr[482]), .rdlo_out(a10_wr[483]));
			radix2 #(.width(width)) rd_st9_484  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[484]), .rdlo_in(a9_wr[485]),  .coef_in(coef[0]), .rdup_out(a10_wr[484]), .rdlo_out(a10_wr[485]));
			radix2 #(.width(width)) rd_st9_486  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[486]), .rdlo_in(a9_wr[487]),  .coef_in(coef[0]), .rdup_out(a10_wr[486]), .rdlo_out(a10_wr[487]));
			radix2 #(.width(width)) rd_st9_488  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[488]), .rdlo_in(a9_wr[489]),  .coef_in(coef[0]), .rdup_out(a10_wr[488]), .rdlo_out(a10_wr[489]));
			radix2 #(.width(width)) rd_st9_490  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[490]), .rdlo_in(a9_wr[491]),  .coef_in(coef[0]), .rdup_out(a10_wr[490]), .rdlo_out(a10_wr[491]));
			radix2 #(.width(width)) rd_st9_492  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[492]), .rdlo_in(a9_wr[493]),  .coef_in(coef[0]), .rdup_out(a10_wr[492]), .rdlo_out(a10_wr[493]));
			radix2 #(.width(width)) rd_st9_494  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[494]), .rdlo_in(a9_wr[495]),  .coef_in(coef[0]), .rdup_out(a10_wr[494]), .rdlo_out(a10_wr[495]));
			radix2 #(.width(width)) rd_st9_496  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[496]), .rdlo_in(a9_wr[497]),  .coef_in(coef[0]), .rdup_out(a10_wr[496]), .rdlo_out(a10_wr[497]));
			radix2 #(.width(width)) rd_st9_498  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[498]), .rdlo_in(a9_wr[499]),  .coef_in(coef[0]), .rdup_out(a10_wr[498]), .rdlo_out(a10_wr[499]));
			radix2 #(.width(width)) rd_st9_500  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[500]), .rdlo_in(a9_wr[501]),  .coef_in(coef[0]), .rdup_out(a10_wr[500]), .rdlo_out(a10_wr[501]));
			radix2 #(.width(width)) rd_st9_502  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[502]), .rdlo_in(a9_wr[503]),  .coef_in(coef[0]), .rdup_out(a10_wr[502]), .rdlo_out(a10_wr[503]));
			radix2 #(.width(width)) rd_st9_504  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[504]), .rdlo_in(a9_wr[505]),  .coef_in(coef[0]), .rdup_out(a10_wr[504]), .rdlo_out(a10_wr[505]));
			radix2 #(.width(width)) rd_st9_506  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[506]), .rdlo_in(a9_wr[507]),  .coef_in(coef[0]), .rdup_out(a10_wr[506]), .rdlo_out(a10_wr[507]));
			radix2 #(.width(width)) rd_st9_508  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[508]), .rdlo_in(a9_wr[509]),  .coef_in(coef[0]), .rdup_out(a10_wr[508]), .rdlo_out(a10_wr[509]));
			radix2 #(.width(width)) rd_st9_510  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[510]), .rdlo_in(a9_wr[511]),  .coef_in(coef[0]), .rdup_out(a10_wr[510]), .rdlo_out(a10_wr[511]));
			radix2 #(.width(width)) rd_st9_512  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[512]), .rdlo_in(a9_wr[513]),  .coef_in(coef[0]), .rdup_out(a10_wr[512]), .rdlo_out(a10_wr[513]));
			radix2 #(.width(width)) rd_st9_514  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[514]), .rdlo_in(a9_wr[515]),  .coef_in(coef[0]), .rdup_out(a10_wr[514]), .rdlo_out(a10_wr[515]));
			radix2 #(.width(width)) rd_st9_516  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[516]), .rdlo_in(a9_wr[517]),  .coef_in(coef[0]), .rdup_out(a10_wr[516]), .rdlo_out(a10_wr[517]));
			radix2 #(.width(width)) rd_st9_518  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[518]), .rdlo_in(a9_wr[519]),  .coef_in(coef[0]), .rdup_out(a10_wr[518]), .rdlo_out(a10_wr[519]));
			radix2 #(.width(width)) rd_st9_520  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[520]), .rdlo_in(a9_wr[521]),  .coef_in(coef[0]), .rdup_out(a10_wr[520]), .rdlo_out(a10_wr[521]));
			radix2 #(.width(width)) rd_st9_522  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[522]), .rdlo_in(a9_wr[523]),  .coef_in(coef[0]), .rdup_out(a10_wr[522]), .rdlo_out(a10_wr[523]));
			radix2 #(.width(width)) rd_st9_524  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[524]), .rdlo_in(a9_wr[525]),  .coef_in(coef[0]), .rdup_out(a10_wr[524]), .rdlo_out(a10_wr[525]));
			radix2 #(.width(width)) rd_st9_526  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[526]), .rdlo_in(a9_wr[527]),  .coef_in(coef[0]), .rdup_out(a10_wr[526]), .rdlo_out(a10_wr[527]));
			radix2 #(.width(width)) rd_st9_528  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[528]), .rdlo_in(a9_wr[529]),  .coef_in(coef[0]), .rdup_out(a10_wr[528]), .rdlo_out(a10_wr[529]));
			radix2 #(.width(width)) rd_st9_530  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[530]), .rdlo_in(a9_wr[531]),  .coef_in(coef[0]), .rdup_out(a10_wr[530]), .rdlo_out(a10_wr[531]));
			radix2 #(.width(width)) rd_st9_532  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[532]), .rdlo_in(a9_wr[533]),  .coef_in(coef[0]), .rdup_out(a10_wr[532]), .rdlo_out(a10_wr[533]));
			radix2 #(.width(width)) rd_st9_534  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[534]), .rdlo_in(a9_wr[535]),  .coef_in(coef[0]), .rdup_out(a10_wr[534]), .rdlo_out(a10_wr[535]));
			radix2 #(.width(width)) rd_st9_536  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[536]), .rdlo_in(a9_wr[537]),  .coef_in(coef[0]), .rdup_out(a10_wr[536]), .rdlo_out(a10_wr[537]));
			radix2 #(.width(width)) rd_st9_538  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[538]), .rdlo_in(a9_wr[539]),  .coef_in(coef[0]), .rdup_out(a10_wr[538]), .rdlo_out(a10_wr[539]));
			radix2 #(.width(width)) rd_st9_540  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[540]), .rdlo_in(a9_wr[541]),  .coef_in(coef[0]), .rdup_out(a10_wr[540]), .rdlo_out(a10_wr[541]));
			radix2 #(.width(width)) rd_st9_542  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[542]), .rdlo_in(a9_wr[543]),  .coef_in(coef[0]), .rdup_out(a10_wr[542]), .rdlo_out(a10_wr[543]));
			radix2 #(.width(width)) rd_st9_544  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[544]), .rdlo_in(a9_wr[545]),  .coef_in(coef[0]), .rdup_out(a10_wr[544]), .rdlo_out(a10_wr[545]));
			radix2 #(.width(width)) rd_st9_546  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[546]), .rdlo_in(a9_wr[547]),  .coef_in(coef[0]), .rdup_out(a10_wr[546]), .rdlo_out(a10_wr[547]));
			radix2 #(.width(width)) rd_st9_548  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[548]), .rdlo_in(a9_wr[549]),  .coef_in(coef[0]), .rdup_out(a10_wr[548]), .rdlo_out(a10_wr[549]));
			radix2 #(.width(width)) rd_st9_550  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[550]), .rdlo_in(a9_wr[551]),  .coef_in(coef[0]), .rdup_out(a10_wr[550]), .rdlo_out(a10_wr[551]));
			radix2 #(.width(width)) rd_st9_552  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[552]), .rdlo_in(a9_wr[553]),  .coef_in(coef[0]), .rdup_out(a10_wr[552]), .rdlo_out(a10_wr[553]));
			radix2 #(.width(width)) rd_st9_554  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[554]), .rdlo_in(a9_wr[555]),  .coef_in(coef[0]), .rdup_out(a10_wr[554]), .rdlo_out(a10_wr[555]));
			radix2 #(.width(width)) rd_st9_556  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[556]), .rdlo_in(a9_wr[557]),  .coef_in(coef[0]), .rdup_out(a10_wr[556]), .rdlo_out(a10_wr[557]));
			radix2 #(.width(width)) rd_st9_558  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[558]), .rdlo_in(a9_wr[559]),  .coef_in(coef[0]), .rdup_out(a10_wr[558]), .rdlo_out(a10_wr[559]));
			radix2 #(.width(width)) rd_st9_560  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[560]), .rdlo_in(a9_wr[561]),  .coef_in(coef[0]), .rdup_out(a10_wr[560]), .rdlo_out(a10_wr[561]));
			radix2 #(.width(width)) rd_st9_562  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[562]), .rdlo_in(a9_wr[563]),  .coef_in(coef[0]), .rdup_out(a10_wr[562]), .rdlo_out(a10_wr[563]));
			radix2 #(.width(width)) rd_st9_564  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[564]), .rdlo_in(a9_wr[565]),  .coef_in(coef[0]), .rdup_out(a10_wr[564]), .rdlo_out(a10_wr[565]));
			radix2 #(.width(width)) rd_st9_566  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[566]), .rdlo_in(a9_wr[567]),  .coef_in(coef[0]), .rdup_out(a10_wr[566]), .rdlo_out(a10_wr[567]));
			radix2 #(.width(width)) rd_st9_568  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[568]), .rdlo_in(a9_wr[569]),  .coef_in(coef[0]), .rdup_out(a10_wr[568]), .rdlo_out(a10_wr[569]));
			radix2 #(.width(width)) rd_st9_570  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[570]), .rdlo_in(a9_wr[571]),  .coef_in(coef[0]), .rdup_out(a10_wr[570]), .rdlo_out(a10_wr[571]));
			radix2 #(.width(width)) rd_st9_572  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[572]), .rdlo_in(a9_wr[573]),  .coef_in(coef[0]), .rdup_out(a10_wr[572]), .rdlo_out(a10_wr[573]));
			radix2 #(.width(width)) rd_st9_574  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[574]), .rdlo_in(a9_wr[575]),  .coef_in(coef[0]), .rdup_out(a10_wr[574]), .rdlo_out(a10_wr[575]));
			radix2 #(.width(width)) rd_st9_576  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[576]), .rdlo_in(a9_wr[577]),  .coef_in(coef[0]), .rdup_out(a10_wr[576]), .rdlo_out(a10_wr[577]));
			radix2 #(.width(width)) rd_st9_578  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[578]), .rdlo_in(a9_wr[579]),  .coef_in(coef[0]), .rdup_out(a10_wr[578]), .rdlo_out(a10_wr[579]));
			radix2 #(.width(width)) rd_st9_580  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[580]), .rdlo_in(a9_wr[581]),  .coef_in(coef[0]), .rdup_out(a10_wr[580]), .rdlo_out(a10_wr[581]));
			radix2 #(.width(width)) rd_st9_582  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[582]), .rdlo_in(a9_wr[583]),  .coef_in(coef[0]), .rdup_out(a10_wr[582]), .rdlo_out(a10_wr[583]));
			radix2 #(.width(width)) rd_st9_584  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[584]), .rdlo_in(a9_wr[585]),  .coef_in(coef[0]), .rdup_out(a10_wr[584]), .rdlo_out(a10_wr[585]));
			radix2 #(.width(width)) rd_st9_586  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[586]), .rdlo_in(a9_wr[587]),  .coef_in(coef[0]), .rdup_out(a10_wr[586]), .rdlo_out(a10_wr[587]));
			radix2 #(.width(width)) rd_st9_588  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[588]), .rdlo_in(a9_wr[589]),  .coef_in(coef[0]), .rdup_out(a10_wr[588]), .rdlo_out(a10_wr[589]));
			radix2 #(.width(width)) rd_st9_590  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[590]), .rdlo_in(a9_wr[591]),  .coef_in(coef[0]), .rdup_out(a10_wr[590]), .rdlo_out(a10_wr[591]));
			radix2 #(.width(width)) rd_st9_592  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[592]), .rdlo_in(a9_wr[593]),  .coef_in(coef[0]), .rdup_out(a10_wr[592]), .rdlo_out(a10_wr[593]));
			radix2 #(.width(width)) rd_st9_594  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[594]), .rdlo_in(a9_wr[595]),  .coef_in(coef[0]), .rdup_out(a10_wr[594]), .rdlo_out(a10_wr[595]));
			radix2 #(.width(width)) rd_st9_596  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[596]), .rdlo_in(a9_wr[597]),  .coef_in(coef[0]), .rdup_out(a10_wr[596]), .rdlo_out(a10_wr[597]));
			radix2 #(.width(width)) rd_st9_598  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[598]), .rdlo_in(a9_wr[599]),  .coef_in(coef[0]), .rdup_out(a10_wr[598]), .rdlo_out(a10_wr[599]));
			radix2 #(.width(width)) rd_st9_600  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[600]), .rdlo_in(a9_wr[601]),  .coef_in(coef[0]), .rdup_out(a10_wr[600]), .rdlo_out(a10_wr[601]));
			radix2 #(.width(width)) rd_st9_602  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[602]), .rdlo_in(a9_wr[603]),  .coef_in(coef[0]), .rdup_out(a10_wr[602]), .rdlo_out(a10_wr[603]));
			radix2 #(.width(width)) rd_st9_604  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[604]), .rdlo_in(a9_wr[605]),  .coef_in(coef[0]), .rdup_out(a10_wr[604]), .rdlo_out(a10_wr[605]));
			radix2 #(.width(width)) rd_st9_606  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[606]), .rdlo_in(a9_wr[607]),  .coef_in(coef[0]), .rdup_out(a10_wr[606]), .rdlo_out(a10_wr[607]));
			radix2 #(.width(width)) rd_st9_608  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[608]), .rdlo_in(a9_wr[609]),  .coef_in(coef[0]), .rdup_out(a10_wr[608]), .rdlo_out(a10_wr[609]));
			radix2 #(.width(width)) rd_st9_610  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[610]), .rdlo_in(a9_wr[611]),  .coef_in(coef[0]), .rdup_out(a10_wr[610]), .rdlo_out(a10_wr[611]));
			radix2 #(.width(width)) rd_st9_612  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[612]), .rdlo_in(a9_wr[613]),  .coef_in(coef[0]), .rdup_out(a10_wr[612]), .rdlo_out(a10_wr[613]));
			radix2 #(.width(width)) rd_st9_614  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[614]), .rdlo_in(a9_wr[615]),  .coef_in(coef[0]), .rdup_out(a10_wr[614]), .rdlo_out(a10_wr[615]));
			radix2 #(.width(width)) rd_st9_616  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[616]), .rdlo_in(a9_wr[617]),  .coef_in(coef[0]), .rdup_out(a10_wr[616]), .rdlo_out(a10_wr[617]));
			radix2 #(.width(width)) rd_st9_618  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[618]), .rdlo_in(a9_wr[619]),  .coef_in(coef[0]), .rdup_out(a10_wr[618]), .rdlo_out(a10_wr[619]));
			radix2 #(.width(width)) rd_st9_620  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[620]), .rdlo_in(a9_wr[621]),  .coef_in(coef[0]), .rdup_out(a10_wr[620]), .rdlo_out(a10_wr[621]));
			radix2 #(.width(width)) rd_st9_622  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[622]), .rdlo_in(a9_wr[623]),  .coef_in(coef[0]), .rdup_out(a10_wr[622]), .rdlo_out(a10_wr[623]));
			radix2 #(.width(width)) rd_st9_624  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[624]), .rdlo_in(a9_wr[625]),  .coef_in(coef[0]), .rdup_out(a10_wr[624]), .rdlo_out(a10_wr[625]));
			radix2 #(.width(width)) rd_st9_626  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[626]), .rdlo_in(a9_wr[627]),  .coef_in(coef[0]), .rdup_out(a10_wr[626]), .rdlo_out(a10_wr[627]));
			radix2 #(.width(width)) rd_st9_628  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[628]), .rdlo_in(a9_wr[629]),  .coef_in(coef[0]), .rdup_out(a10_wr[628]), .rdlo_out(a10_wr[629]));
			radix2 #(.width(width)) rd_st9_630  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[630]), .rdlo_in(a9_wr[631]),  .coef_in(coef[0]), .rdup_out(a10_wr[630]), .rdlo_out(a10_wr[631]));
			radix2 #(.width(width)) rd_st9_632  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[632]), .rdlo_in(a9_wr[633]),  .coef_in(coef[0]), .rdup_out(a10_wr[632]), .rdlo_out(a10_wr[633]));
			radix2 #(.width(width)) rd_st9_634  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[634]), .rdlo_in(a9_wr[635]),  .coef_in(coef[0]), .rdup_out(a10_wr[634]), .rdlo_out(a10_wr[635]));
			radix2 #(.width(width)) rd_st9_636  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[636]), .rdlo_in(a9_wr[637]),  .coef_in(coef[0]), .rdup_out(a10_wr[636]), .rdlo_out(a10_wr[637]));
			radix2 #(.width(width)) rd_st9_638  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[638]), .rdlo_in(a9_wr[639]),  .coef_in(coef[0]), .rdup_out(a10_wr[638]), .rdlo_out(a10_wr[639]));
			radix2 #(.width(width)) rd_st9_640  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[640]), .rdlo_in(a9_wr[641]),  .coef_in(coef[0]), .rdup_out(a10_wr[640]), .rdlo_out(a10_wr[641]));
			radix2 #(.width(width)) rd_st9_642  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[642]), .rdlo_in(a9_wr[643]),  .coef_in(coef[0]), .rdup_out(a10_wr[642]), .rdlo_out(a10_wr[643]));
			radix2 #(.width(width)) rd_st9_644  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[644]), .rdlo_in(a9_wr[645]),  .coef_in(coef[0]), .rdup_out(a10_wr[644]), .rdlo_out(a10_wr[645]));
			radix2 #(.width(width)) rd_st9_646  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[646]), .rdlo_in(a9_wr[647]),  .coef_in(coef[0]), .rdup_out(a10_wr[646]), .rdlo_out(a10_wr[647]));
			radix2 #(.width(width)) rd_st9_648  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[648]), .rdlo_in(a9_wr[649]),  .coef_in(coef[0]), .rdup_out(a10_wr[648]), .rdlo_out(a10_wr[649]));
			radix2 #(.width(width)) rd_st9_650  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[650]), .rdlo_in(a9_wr[651]),  .coef_in(coef[0]), .rdup_out(a10_wr[650]), .rdlo_out(a10_wr[651]));
			radix2 #(.width(width)) rd_st9_652  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[652]), .rdlo_in(a9_wr[653]),  .coef_in(coef[0]), .rdup_out(a10_wr[652]), .rdlo_out(a10_wr[653]));
			radix2 #(.width(width)) rd_st9_654  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[654]), .rdlo_in(a9_wr[655]),  .coef_in(coef[0]), .rdup_out(a10_wr[654]), .rdlo_out(a10_wr[655]));
			radix2 #(.width(width)) rd_st9_656  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[656]), .rdlo_in(a9_wr[657]),  .coef_in(coef[0]), .rdup_out(a10_wr[656]), .rdlo_out(a10_wr[657]));
			radix2 #(.width(width)) rd_st9_658  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[658]), .rdlo_in(a9_wr[659]),  .coef_in(coef[0]), .rdup_out(a10_wr[658]), .rdlo_out(a10_wr[659]));
			radix2 #(.width(width)) rd_st9_660  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[660]), .rdlo_in(a9_wr[661]),  .coef_in(coef[0]), .rdup_out(a10_wr[660]), .rdlo_out(a10_wr[661]));
			radix2 #(.width(width)) rd_st9_662  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[662]), .rdlo_in(a9_wr[663]),  .coef_in(coef[0]), .rdup_out(a10_wr[662]), .rdlo_out(a10_wr[663]));
			radix2 #(.width(width)) rd_st9_664  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[664]), .rdlo_in(a9_wr[665]),  .coef_in(coef[0]), .rdup_out(a10_wr[664]), .rdlo_out(a10_wr[665]));
			radix2 #(.width(width)) rd_st9_666  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[666]), .rdlo_in(a9_wr[667]),  .coef_in(coef[0]), .rdup_out(a10_wr[666]), .rdlo_out(a10_wr[667]));
			radix2 #(.width(width)) rd_st9_668  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[668]), .rdlo_in(a9_wr[669]),  .coef_in(coef[0]), .rdup_out(a10_wr[668]), .rdlo_out(a10_wr[669]));
			radix2 #(.width(width)) rd_st9_670  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[670]), .rdlo_in(a9_wr[671]),  .coef_in(coef[0]), .rdup_out(a10_wr[670]), .rdlo_out(a10_wr[671]));
			radix2 #(.width(width)) rd_st9_672  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[672]), .rdlo_in(a9_wr[673]),  .coef_in(coef[0]), .rdup_out(a10_wr[672]), .rdlo_out(a10_wr[673]));
			radix2 #(.width(width)) rd_st9_674  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[674]), .rdlo_in(a9_wr[675]),  .coef_in(coef[0]), .rdup_out(a10_wr[674]), .rdlo_out(a10_wr[675]));
			radix2 #(.width(width)) rd_st9_676  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[676]), .rdlo_in(a9_wr[677]),  .coef_in(coef[0]), .rdup_out(a10_wr[676]), .rdlo_out(a10_wr[677]));
			radix2 #(.width(width)) rd_st9_678  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[678]), .rdlo_in(a9_wr[679]),  .coef_in(coef[0]), .rdup_out(a10_wr[678]), .rdlo_out(a10_wr[679]));
			radix2 #(.width(width)) rd_st9_680  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[680]), .rdlo_in(a9_wr[681]),  .coef_in(coef[0]), .rdup_out(a10_wr[680]), .rdlo_out(a10_wr[681]));
			radix2 #(.width(width)) rd_st9_682  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[682]), .rdlo_in(a9_wr[683]),  .coef_in(coef[0]), .rdup_out(a10_wr[682]), .rdlo_out(a10_wr[683]));
			radix2 #(.width(width)) rd_st9_684  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[684]), .rdlo_in(a9_wr[685]),  .coef_in(coef[0]), .rdup_out(a10_wr[684]), .rdlo_out(a10_wr[685]));
			radix2 #(.width(width)) rd_st9_686  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[686]), .rdlo_in(a9_wr[687]),  .coef_in(coef[0]), .rdup_out(a10_wr[686]), .rdlo_out(a10_wr[687]));
			radix2 #(.width(width)) rd_st9_688  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[688]), .rdlo_in(a9_wr[689]),  .coef_in(coef[0]), .rdup_out(a10_wr[688]), .rdlo_out(a10_wr[689]));
			radix2 #(.width(width)) rd_st9_690  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[690]), .rdlo_in(a9_wr[691]),  .coef_in(coef[0]), .rdup_out(a10_wr[690]), .rdlo_out(a10_wr[691]));
			radix2 #(.width(width)) rd_st9_692  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[692]), .rdlo_in(a9_wr[693]),  .coef_in(coef[0]), .rdup_out(a10_wr[692]), .rdlo_out(a10_wr[693]));
			radix2 #(.width(width)) rd_st9_694  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[694]), .rdlo_in(a9_wr[695]),  .coef_in(coef[0]), .rdup_out(a10_wr[694]), .rdlo_out(a10_wr[695]));
			radix2 #(.width(width)) rd_st9_696  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[696]), .rdlo_in(a9_wr[697]),  .coef_in(coef[0]), .rdup_out(a10_wr[696]), .rdlo_out(a10_wr[697]));
			radix2 #(.width(width)) rd_st9_698  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[698]), .rdlo_in(a9_wr[699]),  .coef_in(coef[0]), .rdup_out(a10_wr[698]), .rdlo_out(a10_wr[699]));
			radix2 #(.width(width)) rd_st9_700  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[700]), .rdlo_in(a9_wr[701]),  .coef_in(coef[0]), .rdup_out(a10_wr[700]), .rdlo_out(a10_wr[701]));
			radix2 #(.width(width)) rd_st9_702  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[702]), .rdlo_in(a9_wr[703]),  .coef_in(coef[0]), .rdup_out(a10_wr[702]), .rdlo_out(a10_wr[703]));
			radix2 #(.width(width)) rd_st9_704  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[704]), .rdlo_in(a9_wr[705]),  .coef_in(coef[0]), .rdup_out(a10_wr[704]), .rdlo_out(a10_wr[705]));
			radix2 #(.width(width)) rd_st9_706  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[706]), .rdlo_in(a9_wr[707]),  .coef_in(coef[0]), .rdup_out(a10_wr[706]), .rdlo_out(a10_wr[707]));
			radix2 #(.width(width)) rd_st9_708  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[708]), .rdlo_in(a9_wr[709]),  .coef_in(coef[0]), .rdup_out(a10_wr[708]), .rdlo_out(a10_wr[709]));
			radix2 #(.width(width)) rd_st9_710  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[710]), .rdlo_in(a9_wr[711]),  .coef_in(coef[0]), .rdup_out(a10_wr[710]), .rdlo_out(a10_wr[711]));
			radix2 #(.width(width)) rd_st9_712  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[712]), .rdlo_in(a9_wr[713]),  .coef_in(coef[0]), .rdup_out(a10_wr[712]), .rdlo_out(a10_wr[713]));
			radix2 #(.width(width)) rd_st9_714  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[714]), .rdlo_in(a9_wr[715]),  .coef_in(coef[0]), .rdup_out(a10_wr[714]), .rdlo_out(a10_wr[715]));
			radix2 #(.width(width)) rd_st9_716  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[716]), .rdlo_in(a9_wr[717]),  .coef_in(coef[0]), .rdup_out(a10_wr[716]), .rdlo_out(a10_wr[717]));
			radix2 #(.width(width)) rd_st9_718  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[718]), .rdlo_in(a9_wr[719]),  .coef_in(coef[0]), .rdup_out(a10_wr[718]), .rdlo_out(a10_wr[719]));
			radix2 #(.width(width)) rd_st9_720  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[720]), .rdlo_in(a9_wr[721]),  .coef_in(coef[0]), .rdup_out(a10_wr[720]), .rdlo_out(a10_wr[721]));
			radix2 #(.width(width)) rd_st9_722  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[722]), .rdlo_in(a9_wr[723]),  .coef_in(coef[0]), .rdup_out(a10_wr[722]), .rdlo_out(a10_wr[723]));
			radix2 #(.width(width)) rd_st9_724  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[724]), .rdlo_in(a9_wr[725]),  .coef_in(coef[0]), .rdup_out(a10_wr[724]), .rdlo_out(a10_wr[725]));
			radix2 #(.width(width)) rd_st9_726  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[726]), .rdlo_in(a9_wr[727]),  .coef_in(coef[0]), .rdup_out(a10_wr[726]), .rdlo_out(a10_wr[727]));
			radix2 #(.width(width)) rd_st9_728  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[728]), .rdlo_in(a9_wr[729]),  .coef_in(coef[0]), .rdup_out(a10_wr[728]), .rdlo_out(a10_wr[729]));
			radix2 #(.width(width)) rd_st9_730  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[730]), .rdlo_in(a9_wr[731]),  .coef_in(coef[0]), .rdup_out(a10_wr[730]), .rdlo_out(a10_wr[731]));
			radix2 #(.width(width)) rd_st9_732  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[732]), .rdlo_in(a9_wr[733]),  .coef_in(coef[0]), .rdup_out(a10_wr[732]), .rdlo_out(a10_wr[733]));
			radix2 #(.width(width)) rd_st9_734  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[734]), .rdlo_in(a9_wr[735]),  .coef_in(coef[0]), .rdup_out(a10_wr[734]), .rdlo_out(a10_wr[735]));
			radix2 #(.width(width)) rd_st9_736  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[736]), .rdlo_in(a9_wr[737]),  .coef_in(coef[0]), .rdup_out(a10_wr[736]), .rdlo_out(a10_wr[737]));
			radix2 #(.width(width)) rd_st9_738  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[738]), .rdlo_in(a9_wr[739]),  .coef_in(coef[0]), .rdup_out(a10_wr[738]), .rdlo_out(a10_wr[739]));
			radix2 #(.width(width)) rd_st9_740  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[740]), .rdlo_in(a9_wr[741]),  .coef_in(coef[0]), .rdup_out(a10_wr[740]), .rdlo_out(a10_wr[741]));
			radix2 #(.width(width)) rd_st9_742  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[742]), .rdlo_in(a9_wr[743]),  .coef_in(coef[0]), .rdup_out(a10_wr[742]), .rdlo_out(a10_wr[743]));
			radix2 #(.width(width)) rd_st9_744  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[744]), .rdlo_in(a9_wr[745]),  .coef_in(coef[0]), .rdup_out(a10_wr[744]), .rdlo_out(a10_wr[745]));
			radix2 #(.width(width)) rd_st9_746  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[746]), .rdlo_in(a9_wr[747]),  .coef_in(coef[0]), .rdup_out(a10_wr[746]), .rdlo_out(a10_wr[747]));
			radix2 #(.width(width)) rd_st9_748  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[748]), .rdlo_in(a9_wr[749]),  .coef_in(coef[0]), .rdup_out(a10_wr[748]), .rdlo_out(a10_wr[749]));
			radix2 #(.width(width)) rd_st9_750  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[750]), .rdlo_in(a9_wr[751]),  .coef_in(coef[0]), .rdup_out(a10_wr[750]), .rdlo_out(a10_wr[751]));
			radix2 #(.width(width)) rd_st9_752  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[752]), .rdlo_in(a9_wr[753]),  .coef_in(coef[0]), .rdup_out(a10_wr[752]), .rdlo_out(a10_wr[753]));
			radix2 #(.width(width)) rd_st9_754  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[754]), .rdlo_in(a9_wr[755]),  .coef_in(coef[0]), .rdup_out(a10_wr[754]), .rdlo_out(a10_wr[755]));
			radix2 #(.width(width)) rd_st9_756  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[756]), .rdlo_in(a9_wr[757]),  .coef_in(coef[0]), .rdup_out(a10_wr[756]), .rdlo_out(a10_wr[757]));
			radix2 #(.width(width)) rd_st9_758  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[758]), .rdlo_in(a9_wr[759]),  .coef_in(coef[0]), .rdup_out(a10_wr[758]), .rdlo_out(a10_wr[759]));
			radix2 #(.width(width)) rd_st9_760  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[760]), .rdlo_in(a9_wr[761]),  .coef_in(coef[0]), .rdup_out(a10_wr[760]), .rdlo_out(a10_wr[761]));
			radix2 #(.width(width)) rd_st9_762  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[762]), .rdlo_in(a9_wr[763]),  .coef_in(coef[0]), .rdup_out(a10_wr[762]), .rdlo_out(a10_wr[763]));
			radix2 #(.width(width)) rd_st9_764  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[764]), .rdlo_in(a9_wr[765]),  .coef_in(coef[0]), .rdup_out(a10_wr[764]), .rdlo_out(a10_wr[765]));
			radix2 #(.width(width)) rd_st9_766  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[766]), .rdlo_in(a9_wr[767]),  .coef_in(coef[0]), .rdup_out(a10_wr[766]), .rdlo_out(a10_wr[767]));
			radix2 #(.width(width)) rd_st9_768  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[768]), .rdlo_in(a9_wr[769]),  .coef_in(coef[0]), .rdup_out(a10_wr[768]), .rdlo_out(a10_wr[769]));
			radix2 #(.width(width)) rd_st9_770  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[770]), .rdlo_in(a9_wr[771]),  .coef_in(coef[0]), .rdup_out(a10_wr[770]), .rdlo_out(a10_wr[771]));
			radix2 #(.width(width)) rd_st9_772  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[772]), .rdlo_in(a9_wr[773]),  .coef_in(coef[0]), .rdup_out(a10_wr[772]), .rdlo_out(a10_wr[773]));
			radix2 #(.width(width)) rd_st9_774  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[774]), .rdlo_in(a9_wr[775]),  .coef_in(coef[0]), .rdup_out(a10_wr[774]), .rdlo_out(a10_wr[775]));
			radix2 #(.width(width)) rd_st9_776  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[776]), .rdlo_in(a9_wr[777]),  .coef_in(coef[0]), .rdup_out(a10_wr[776]), .rdlo_out(a10_wr[777]));
			radix2 #(.width(width)) rd_st9_778  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[778]), .rdlo_in(a9_wr[779]),  .coef_in(coef[0]), .rdup_out(a10_wr[778]), .rdlo_out(a10_wr[779]));
			radix2 #(.width(width)) rd_st9_780  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[780]), .rdlo_in(a9_wr[781]),  .coef_in(coef[0]), .rdup_out(a10_wr[780]), .rdlo_out(a10_wr[781]));
			radix2 #(.width(width)) rd_st9_782  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[782]), .rdlo_in(a9_wr[783]),  .coef_in(coef[0]), .rdup_out(a10_wr[782]), .rdlo_out(a10_wr[783]));
			radix2 #(.width(width)) rd_st9_784  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[784]), .rdlo_in(a9_wr[785]),  .coef_in(coef[0]), .rdup_out(a10_wr[784]), .rdlo_out(a10_wr[785]));
			radix2 #(.width(width)) rd_st9_786  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[786]), .rdlo_in(a9_wr[787]),  .coef_in(coef[0]), .rdup_out(a10_wr[786]), .rdlo_out(a10_wr[787]));
			radix2 #(.width(width)) rd_st9_788  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[788]), .rdlo_in(a9_wr[789]),  .coef_in(coef[0]), .rdup_out(a10_wr[788]), .rdlo_out(a10_wr[789]));
			radix2 #(.width(width)) rd_st9_790  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[790]), .rdlo_in(a9_wr[791]),  .coef_in(coef[0]), .rdup_out(a10_wr[790]), .rdlo_out(a10_wr[791]));
			radix2 #(.width(width)) rd_st9_792  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[792]), .rdlo_in(a9_wr[793]),  .coef_in(coef[0]), .rdup_out(a10_wr[792]), .rdlo_out(a10_wr[793]));
			radix2 #(.width(width)) rd_st9_794  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[794]), .rdlo_in(a9_wr[795]),  .coef_in(coef[0]), .rdup_out(a10_wr[794]), .rdlo_out(a10_wr[795]));
			radix2 #(.width(width)) rd_st9_796  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[796]), .rdlo_in(a9_wr[797]),  .coef_in(coef[0]), .rdup_out(a10_wr[796]), .rdlo_out(a10_wr[797]));
			radix2 #(.width(width)) rd_st9_798  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[798]), .rdlo_in(a9_wr[799]),  .coef_in(coef[0]), .rdup_out(a10_wr[798]), .rdlo_out(a10_wr[799]));
			radix2 #(.width(width)) rd_st9_800  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[800]), .rdlo_in(a9_wr[801]),  .coef_in(coef[0]), .rdup_out(a10_wr[800]), .rdlo_out(a10_wr[801]));
			radix2 #(.width(width)) rd_st9_802  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[802]), .rdlo_in(a9_wr[803]),  .coef_in(coef[0]), .rdup_out(a10_wr[802]), .rdlo_out(a10_wr[803]));
			radix2 #(.width(width)) rd_st9_804  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[804]), .rdlo_in(a9_wr[805]),  .coef_in(coef[0]), .rdup_out(a10_wr[804]), .rdlo_out(a10_wr[805]));
			radix2 #(.width(width)) rd_st9_806  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[806]), .rdlo_in(a9_wr[807]),  .coef_in(coef[0]), .rdup_out(a10_wr[806]), .rdlo_out(a10_wr[807]));
			radix2 #(.width(width)) rd_st9_808  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[808]), .rdlo_in(a9_wr[809]),  .coef_in(coef[0]), .rdup_out(a10_wr[808]), .rdlo_out(a10_wr[809]));
			radix2 #(.width(width)) rd_st9_810  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[810]), .rdlo_in(a9_wr[811]),  .coef_in(coef[0]), .rdup_out(a10_wr[810]), .rdlo_out(a10_wr[811]));
			radix2 #(.width(width)) rd_st9_812  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[812]), .rdlo_in(a9_wr[813]),  .coef_in(coef[0]), .rdup_out(a10_wr[812]), .rdlo_out(a10_wr[813]));
			radix2 #(.width(width)) rd_st9_814  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[814]), .rdlo_in(a9_wr[815]),  .coef_in(coef[0]), .rdup_out(a10_wr[814]), .rdlo_out(a10_wr[815]));
			radix2 #(.width(width)) rd_st9_816  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[816]), .rdlo_in(a9_wr[817]),  .coef_in(coef[0]), .rdup_out(a10_wr[816]), .rdlo_out(a10_wr[817]));
			radix2 #(.width(width)) rd_st9_818  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[818]), .rdlo_in(a9_wr[819]),  .coef_in(coef[0]), .rdup_out(a10_wr[818]), .rdlo_out(a10_wr[819]));
			radix2 #(.width(width)) rd_st9_820  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[820]), .rdlo_in(a9_wr[821]),  .coef_in(coef[0]), .rdup_out(a10_wr[820]), .rdlo_out(a10_wr[821]));
			radix2 #(.width(width)) rd_st9_822  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[822]), .rdlo_in(a9_wr[823]),  .coef_in(coef[0]), .rdup_out(a10_wr[822]), .rdlo_out(a10_wr[823]));
			radix2 #(.width(width)) rd_st9_824  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[824]), .rdlo_in(a9_wr[825]),  .coef_in(coef[0]), .rdup_out(a10_wr[824]), .rdlo_out(a10_wr[825]));
			radix2 #(.width(width)) rd_st9_826  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[826]), .rdlo_in(a9_wr[827]),  .coef_in(coef[0]), .rdup_out(a10_wr[826]), .rdlo_out(a10_wr[827]));
			radix2 #(.width(width)) rd_st9_828  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[828]), .rdlo_in(a9_wr[829]),  .coef_in(coef[0]), .rdup_out(a10_wr[828]), .rdlo_out(a10_wr[829]));
			radix2 #(.width(width)) rd_st9_830  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[830]), .rdlo_in(a9_wr[831]),  .coef_in(coef[0]), .rdup_out(a10_wr[830]), .rdlo_out(a10_wr[831]));
			radix2 #(.width(width)) rd_st9_832  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[832]), .rdlo_in(a9_wr[833]),  .coef_in(coef[0]), .rdup_out(a10_wr[832]), .rdlo_out(a10_wr[833]));
			radix2 #(.width(width)) rd_st9_834  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[834]), .rdlo_in(a9_wr[835]),  .coef_in(coef[0]), .rdup_out(a10_wr[834]), .rdlo_out(a10_wr[835]));
			radix2 #(.width(width)) rd_st9_836  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[836]), .rdlo_in(a9_wr[837]),  .coef_in(coef[0]), .rdup_out(a10_wr[836]), .rdlo_out(a10_wr[837]));
			radix2 #(.width(width)) rd_st9_838  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[838]), .rdlo_in(a9_wr[839]),  .coef_in(coef[0]), .rdup_out(a10_wr[838]), .rdlo_out(a10_wr[839]));
			radix2 #(.width(width)) rd_st9_840  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[840]), .rdlo_in(a9_wr[841]),  .coef_in(coef[0]), .rdup_out(a10_wr[840]), .rdlo_out(a10_wr[841]));
			radix2 #(.width(width)) rd_st9_842  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[842]), .rdlo_in(a9_wr[843]),  .coef_in(coef[0]), .rdup_out(a10_wr[842]), .rdlo_out(a10_wr[843]));
			radix2 #(.width(width)) rd_st9_844  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[844]), .rdlo_in(a9_wr[845]),  .coef_in(coef[0]), .rdup_out(a10_wr[844]), .rdlo_out(a10_wr[845]));
			radix2 #(.width(width)) rd_st9_846  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[846]), .rdlo_in(a9_wr[847]),  .coef_in(coef[0]), .rdup_out(a10_wr[846]), .rdlo_out(a10_wr[847]));
			radix2 #(.width(width)) rd_st9_848  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[848]), .rdlo_in(a9_wr[849]),  .coef_in(coef[0]), .rdup_out(a10_wr[848]), .rdlo_out(a10_wr[849]));
			radix2 #(.width(width)) rd_st9_850  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[850]), .rdlo_in(a9_wr[851]),  .coef_in(coef[0]), .rdup_out(a10_wr[850]), .rdlo_out(a10_wr[851]));
			radix2 #(.width(width)) rd_st9_852  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[852]), .rdlo_in(a9_wr[853]),  .coef_in(coef[0]), .rdup_out(a10_wr[852]), .rdlo_out(a10_wr[853]));
			radix2 #(.width(width)) rd_st9_854  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[854]), .rdlo_in(a9_wr[855]),  .coef_in(coef[0]), .rdup_out(a10_wr[854]), .rdlo_out(a10_wr[855]));
			radix2 #(.width(width)) rd_st9_856  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[856]), .rdlo_in(a9_wr[857]),  .coef_in(coef[0]), .rdup_out(a10_wr[856]), .rdlo_out(a10_wr[857]));
			radix2 #(.width(width)) rd_st9_858  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[858]), .rdlo_in(a9_wr[859]),  .coef_in(coef[0]), .rdup_out(a10_wr[858]), .rdlo_out(a10_wr[859]));
			radix2 #(.width(width)) rd_st9_860  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[860]), .rdlo_in(a9_wr[861]),  .coef_in(coef[0]), .rdup_out(a10_wr[860]), .rdlo_out(a10_wr[861]));
			radix2 #(.width(width)) rd_st9_862  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[862]), .rdlo_in(a9_wr[863]),  .coef_in(coef[0]), .rdup_out(a10_wr[862]), .rdlo_out(a10_wr[863]));
			radix2 #(.width(width)) rd_st9_864  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[864]), .rdlo_in(a9_wr[865]),  .coef_in(coef[0]), .rdup_out(a10_wr[864]), .rdlo_out(a10_wr[865]));
			radix2 #(.width(width)) rd_st9_866  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[866]), .rdlo_in(a9_wr[867]),  .coef_in(coef[0]), .rdup_out(a10_wr[866]), .rdlo_out(a10_wr[867]));
			radix2 #(.width(width)) rd_st9_868  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[868]), .rdlo_in(a9_wr[869]),  .coef_in(coef[0]), .rdup_out(a10_wr[868]), .rdlo_out(a10_wr[869]));
			radix2 #(.width(width)) rd_st9_870  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[870]), .rdlo_in(a9_wr[871]),  .coef_in(coef[0]), .rdup_out(a10_wr[870]), .rdlo_out(a10_wr[871]));
			radix2 #(.width(width)) rd_st9_872  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[872]), .rdlo_in(a9_wr[873]),  .coef_in(coef[0]), .rdup_out(a10_wr[872]), .rdlo_out(a10_wr[873]));
			radix2 #(.width(width)) rd_st9_874  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[874]), .rdlo_in(a9_wr[875]),  .coef_in(coef[0]), .rdup_out(a10_wr[874]), .rdlo_out(a10_wr[875]));
			radix2 #(.width(width)) rd_st9_876  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[876]), .rdlo_in(a9_wr[877]),  .coef_in(coef[0]), .rdup_out(a10_wr[876]), .rdlo_out(a10_wr[877]));
			radix2 #(.width(width)) rd_st9_878  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[878]), .rdlo_in(a9_wr[879]),  .coef_in(coef[0]), .rdup_out(a10_wr[878]), .rdlo_out(a10_wr[879]));
			radix2 #(.width(width)) rd_st9_880  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[880]), .rdlo_in(a9_wr[881]),  .coef_in(coef[0]), .rdup_out(a10_wr[880]), .rdlo_out(a10_wr[881]));
			radix2 #(.width(width)) rd_st9_882  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[882]), .rdlo_in(a9_wr[883]),  .coef_in(coef[0]), .rdup_out(a10_wr[882]), .rdlo_out(a10_wr[883]));
			radix2 #(.width(width)) rd_st9_884  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[884]), .rdlo_in(a9_wr[885]),  .coef_in(coef[0]), .rdup_out(a10_wr[884]), .rdlo_out(a10_wr[885]));
			radix2 #(.width(width)) rd_st9_886  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[886]), .rdlo_in(a9_wr[887]),  .coef_in(coef[0]), .rdup_out(a10_wr[886]), .rdlo_out(a10_wr[887]));
			radix2 #(.width(width)) rd_st9_888  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[888]), .rdlo_in(a9_wr[889]),  .coef_in(coef[0]), .rdup_out(a10_wr[888]), .rdlo_out(a10_wr[889]));
			radix2 #(.width(width)) rd_st9_890  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[890]), .rdlo_in(a9_wr[891]),  .coef_in(coef[0]), .rdup_out(a10_wr[890]), .rdlo_out(a10_wr[891]));
			radix2 #(.width(width)) rd_st9_892  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[892]), .rdlo_in(a9_wr[893]),  .coef_in(coef[0]), .rdup_out(a10_wr[892]), .rdlo_out(a10_wr[893]));
			radix2 #(.width(width)) rd_st9_894  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[894]), .rdlo_in(a9_wr[895]),  .coef_in(coef[0]), .rdup_out(a10_wr[894]), .rdlo_out(a10_wr[895]));
			radix2 #(.width(width)) rd_st9_896  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[896]), .rdlo_in(a9_wr[897]),  .coef_in(coef[0]), .rdup_out(a10_wr[896]), .rdlo_out(a10_wr[897]));
			radix2 #(.width(width)) rd_st9_898  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[898]), .rdlo_in(a9_wr[899]),  .coef_in(coef[0]), .rdup_out(a10_wr[898]), .rdlo_out(a10_wr[899]));
			radix2 #(.width(width)) rd_st9_900  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[900]), .rdlo_in(a9_wr[901]),  .coef_in(coef[0]), .rdup_out(a10_wr[900]), .rdlo_out(a10_wr[901]));
			radix2 #(.width(width)) rd_st9_902  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[902]), .rdlo_in(a9_wr[903]),  .coef_in(coef[0]), .rdup_out(a10_wr[902]), .rdlo_out(a10_wr[903]));
			radix2 #(.width(width)) rd_st9_904  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[904]), .rdlo_in(a9_wr[905]),  .coef_in(coef[0]), .rdup_out(a10_wr[904]), .rdlo_out(a10_wr[905]));
			radix2 #(.width(width)) rd_st9_906  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[906]), .rdlo_in(a9_wr[907]),  .coef_in(coef[0]), .rdup_out(a10_wr[906]), .rdlo_out(a10_wr[907]));
			radix2 #(.width(width)) rd_st9_908  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[908]), .rdlo_in(a9_wr[909]),  .coef_in(coef[0]), .rdup_out(a10_wr[908]), .rdlo_out(a10_wr[909]));
			radix2 #(.width(width)) rd_st9_910  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[910]), .rdlo_in(a9_wr[911]),  .coef_in(coef[0]), .rdup_out(a10_wr[910]), .rdlo_out(a10_wr[911]));
			radix2 #(.width(width)) rd_st9_912  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[912]), .rdlo_in(a9_wr[913]),  .coef_in(coef[0]), .rdup_out(a10_wr[912]), .rdlo_out(a10_wr[913]));
			radix2 #(.width(width)) rd_st9_914  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[914]), .rdlo_in(a9_wr[915]),  .coef_in(coef[0]), .rdup_out(a10_wr[914]), .rdlo_out(a10_wr[915]));
			radix2 #(.width(width)) rd_st9_916  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[916]), .rdlo_in(a9_wr[917]),  .coef_in(coef[0]), .rdup_out(a10_wr[916]), .rdlo_out(a10_wr[917]));
			radix2 #(.width(width)) rd_st9_918  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[918]), .rdlo_in(a9_wr[919]),  .coef_in(coef[0]), .rdup_out(a10_wr[918]), .rdlo_out(a10_wr[919]));
			radix2 #(.width(width)) rd_st9_920  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[920]), .rdlo_in(a9_wr[921]),  .coef_in(coef[0]), .rdup_out(a10_wr[920]), .rdlo_out(a10_wr[921]));
			radix2 #(.width(width)) rd_st9_922  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[922]), .rdlo_in(a9_wr[923]),  .coef_in(coef[0]), .rdup_out(a10_wr[922]), .rdlo_out(a10_wr[923]));
			radix2 #(.width(width)) rd_st9_924  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[924]), .rdlo_in(a9_wr[925]),  .coef_in(coef[0]), .rdup_out(a10_wr[924]), .rdlo_out(a10_wr[925]));
			radix2 #(.width(width)) rd_st9_926  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[926]), .rdlo_in(a9_wr[927]),  .coef_in(coef[0]), .rdup_out(a10_wr[926]), .rdlo_out(a10_wr[927]));
			radix2 #(.width(width)) rd_st9_928  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[928]), .rdlo_in(a9_wr[929]),  .coef_in(coef[0]), .rdup_out(a10_wr[928]), .rdlo_out(a10_wr[929]));
			radix2 #(.width(width)) rd_st9_930  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[930]), .rdlo_in(a9_wr[931]),  .coef_in(coef[0]), .rdup_out(a10_wr[930]), .rdlo_out(a10_wr[931]));
			radix2 #(.width(width)) rd_st9_932  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[932]), .rdlo_in(a9_wr[933]),  .coef_in(coef[0]), .rdup_out(a10_wr[932]), .rdlo_out(a10_wr[933]));
			radix2 #(.width(width)) rd_st9_934  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[934]), .rdlo_in(a9_wr[935]),  .coef_in(coef[0]), .rdup_out(a10_wr[934]), .rdlo_out(a10_wr[935]));
			radix2 #(.width(width)) rd_st9_936  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[936]), .rdlo_in(a9_wr[937]),  .coef_in(coef[0]), .rdup_out(a10_wr[936]), .rdlo_out(a10_wr[937]));
			radix2 #(.width(width)) rd_st9_938  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[938]), .rdlo_in(a9_wr[939]),  .coef_in(coef[0]), .rdup_out(a10_wr[938]), .rdlo_out(a10_wr[939]));
			radix2 #(.width(width)) rd_st9_940  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[940]), .rdlo_in(a9_wr[941]),  .coef_in(coef[0]), .rdup_out(a10_wr[940]), .rdlo_out(a10_wr[941]));
			radix2 #(.width(width)) rd_st9_942  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[942]), .rdlo_in(a9_wr[943]),  .coef_in(coef[0]), .rdup_out(a10_wr[942]), .rdlo_out(a10_wr[943]));
			radix2 #(.width(width)) rd_st9_944  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[944]), .rdlo_in(a9_wr[945]),  .coef_in(coef[0]), .rdup_out(a10_wr[944]), .rdlo_out(a10_wr[945]));
			radix2 #(.width(width)) rd_st9_946  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[946]), .rdlo_in(a9_wr[947]),  .coef_in(coef[0]), .rdup_out(a10_wr[946]), .rdlo_out(a10_wr[947]));
			radix2 #(.width(width)) rd_st9_948  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[948]), .rdlo_in(a9_wr[949]),  .coef_in(coef[0]), .rdup_out(a10_wr[948]), .rdlo_out(a10_wr[949]));
			radix2 #(.width(width)) rd_st9_950  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[950]), .rdlo_in(a9_wr[951]),  .coef_in(coef[0]), .rdup_out(a10_wr[950]), .rdlo_out(a10_wr[951]));
			radix2 #(.width(width)) rd_st9_952  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[952]), .rdlo_in(a9_wr[953]),  .coef_in(coef[0]), .rdup_out(a10_wr[952]), .rdlo_out(a10_wr[953]));
			radix2 #(.width(width)) rd_st9_954  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[954]), .rdlo_in(a9_wr[955]),  .coef_in(coef[0]), .rdup_out(a10_wr[954]), .rdlo_out(a10_wr[955]));
			radix2 #(.width(width)) rd_st9_956  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[956]), .rdlo_in(a9_wr[957]),  .coef_in(coef[0]), .rdup_out(a10_wr[956]), .rdlo_out(a10_wr[957]));
			radix2 #(.width(width)) rd_st9_958  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[958]), .rdlo_in(a9_wr[959]),  .coef_in(coef[0]), .rdup_out(a10_wr[958]), .rdlo_out(a10_wr[959]));
			radix2 #(.width(width)) rd_st9_960  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[960]), .rdlo_in(a9_wr[961]),  .coef_in(coef[0]), .rdup_out(a10_wr[960]), .rdlo_out(a10_wr[961]));
			radix2 #(.width(width)) rd_st9_962  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[962]), .rdlo_in(a9_wr[963]),  .coef_in(coef[0]), .rdup_out(a10_wr[962]), .rdlo_out(a10_wr[963]));
			radix2 #(.width(width)) rd_st9_964  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[964]), .rdlo_in(a9_wr[965]),  .coef_in(coef[0]), .rdup_out(a10_wr[964]), .rdlo_out(a10_wr[965]));
			radix2 #(.width(width)) rd_st9_966  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[966]), .rdlo_in(a9_wr[967]),  .coef_in(coef[0]), .rdup_out(a10_wr[966]), .rdlo_out(a10_wr[967]));
			radix2 #(.width(width)) rd_st9_968  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[968]), .rdlo_in(a9_wr[969]),  .coef_in(coef[0]), .rdup_out(a10_wr[968]), .rdlo_out(a10_wr[969]));
			radix2 #(.width(width)) rd_st9_970  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[970]), .rdlo_in(a9_wr[971]),  .coef_in(coef[0]), .rdup_out(a10_wr[970]), .rdlo_out(a10_wr[971]));
			radix2 #(.width(width)) rd_st9_972  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[972]), .rdlo_in(a9_wr[973]),  .coef_in(coef[0]), .rdup_out(a10_wr[972]), .rdlo_out(a10_wr[973]));
			radix2 #(.width(width)) rd_st9_974  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[974]), .rdlo_in(a9_wr[975]),  .coef_in(coef[0]), .rdup_out(a10_wr[974]), .rdlo_out(a10_wr[975]));
			radix2 #(.width(width)) rd_st9_976  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[976]), .rdlo_in(a9_wr[977]),  .coef_in(coef[0]), .rdup_out(a10_wr[976]), .rdlo_out(a10_wr[977]));
			radix2 #(.width(width)) rd_st9_978  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[978]), .rdlo_in(a9_wr[979]),  .coef_in(coef[0]), .rdup_out(a10_wr[978]), .rdlo_out(a10_wr[979]));
			radix2 #(.width(width)) rd_st9_980  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[980]), .rdlo_in(a9_wr[981]),  .coef_in(coef[0]), .rdup_out(a10_wr[980]), .rdlo_out(a10_wr[981]));
			radix2 #(.width(width)) rd_st9_982  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[982]), .rdlo_in(a9_wr[983]),  .coef_in(coef[0]), .rdup_out(a10_wr[982]), .rdlo_out(a10_wr[983]));
			radix2 #(.width(width)) rd_st9_984  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[984]), .rdlo_in(a9_wr[985]),  .coef_in(coef[0]), .rdup_out(a10_wr[984]), .rdlo_out(a10_wr[985]));
			radix2 #(.width(width)) rd_st9_986  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[986]), .rdlo_in(a9_wr[987]),  .coef_in(coef[0]), .rdup_out(a10_wr[986]), .rdlo_out(a10_wr[987]));
			radix2 #(.width(width)) rd_st9_988  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[988]), .rdlo_in(a9_wr[989]),  .coef_in(coef[0]), .rdup_out(a10_wr[988]), .rdlo_out(a10_wr[989]));
			radix2 #(.width(width)) rd_st9_990  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[990]), .rdlo_in(a9_wr[991]),  .coef_in(coef[0]), .rdup_out(a10_wr[990]), .rdlo_out(a10_wr[991]));
			radix2 #(.width(width)) rd_st9_992  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[992]), .rdlo_in(a9_wr[993]),  .coef_in(coef[0]), .rdup_out(a10_wr[992]), .rdlo_out(a10_wr[993]));
			radix2 #(.width(width)) rd_st9_994  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[994]), .rdlo_in(a9_wr[995]),  .coef_in(coef[0]), .rdup_out(a10_wr[994]), .rdlo_out(a10_wr[995]));
			radix2 #(.width(width)) rd_st9_996  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[996]), .rdlo_in(a9_wr[997]),  .coef_in(coef[0]), .rdup_out(a10_wr[996]), .rdlo_out(a10_wr[997]));
			radix2 #(.width(width)) rd_st9_998  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[998]), .rdlo_in(a9_wr[999]),  .coef_in(coef[0]), .rdup_out(a10_wr[998]), .rdlo_out(a10_wr[999]));
			radix2 #(.width(width)) rd_st9_1000  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1000]), .rdlo_in(a9_wr[1001]),  .coef_in(coef[0]), .rdup_out(a10_wr[1000]), .rdlo_out(a10_wr[1001]));
			radix2 #(.width(width)) rd_st9_1002  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1002]), .rdlo_in(a9_wr[1003]),  .coef_in(coef[0]), .rdup_out(a10_wr[1002]), .rdlo_out(a10_wr[1003]));
			radix2 #(.width(width)) rd_st9_1004  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1004]), .rdlo_in(a9_wr[1005]),  .coef_in(coef[0]), .rdup_out(a10_wr[1004]), .rdlo_out(a10_wr[1005]));
			radix2 #(.width(width)) rd_st9_1006  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1006]), .rdlo_in(a9_wr[1007]),  .coef_in(coef[0]), .rdup_out(a10_wr[1006]), .rdlo_out(a10_wr[1007]));
			radix2 #(.width(width)) rd_st9_1008  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1008]), .rdlo_in(a9_wr[1009]),  .coef_in(coef[0]), .rdup_out(a10_wr[1008]), .rdlo_out(a10_wr[1009]));
			radix2 #(.width(width)) rd_st9_1010  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1010]), .rdlo_in(a9_wr[1011]),  .coef_in(coef[0]), .rdup_out(a10_wr[1010]), .rdlo_out(a10_wr[1011]));
			radix2 #(.width(width)) rd_st9_1012  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1012]), .rdlo_in(a9_wr[1013]),  .coef_in(coef[0]), .rdup_out(a10_wr[1012]), .rdlo_out(a10_wr[1013]));
			radix2 #(.width(width)) rd_st9_1014  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1014]), .rdlo_in(a9_wr[1015]),  .coef_in(coef[0]), .rdup_out(a10_wr[1014]), .rdlo_out(a10_wr[1015]));
			radix2 #(.width(width)) rd_st9_1016  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1016]), .rdlo_in(a9_wr[1017]),  .coef_in(coef[0]), .rdup_out(a10_wr[1016]), .rdlo_out(a10_wr[1017]));
			radix2 #(.width(width)) rd_st9_1018  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1018]), .rdlo_in(a9_wr[1019]),  .coef_in(coef[0]), .rdup_out(a10_wr[1018]), .rdlo_out(a10_wr[1019]));
			radix2 #(.width(width)) rd_st9_1020  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1020]), .rdlo_in(a9_wr[1021]),  .coef_in(coef[0]), .rdup_out(a10_wr[1020]), .rdlo_out(a10_wr[1021]));
			radix2 #(.width(width)) rd_st9_1022  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1022]), .rdlo_in(a9_wr[1023]),  .coef_in(coef[0]), .rdup_out(a10_wr[1022]), .rdlo_out(a10_wr[1023]));

		//--- output stage (bit reversal)
			assign x0_out       = a10_wr[0];                   
			assign x1_out       = a10_wr[512];                 
			assign x2_out       = a10_wr[256];                 
			assign x3_out       = a10_wr[768];                 
			assign x4_out       = a10_wr[128];                 
			assign x5_out       = a10_wr[640];                 
			assign x6_out       = a10_wr[384];                 
			assign x7_out       = a10_wr[896];                 
			assign x8_out       = a10_wr[64];                  
			assign x9_out       = a10_wr[576];                 
			assign x10_out      = a10_wr[320];                 
			assign x11_out      = a10_wr[832];                 
			assign x12_out      = a10_wr[192];                 
			assign x13_out      = a10_wr[704];                 
			assign x14_out      = a10_wr[448];                 
			assign x15_out      = a10_wr[960];                 
			assign x16_out      = a10_wr[32];                  
			assign x17_out      = a10_wr[544];                 
			assign x18_out      = a10_wr[288];                 
			assign x19_out      = a10_wr[800];                 
			assign x20_out      = a10_wr[160];                 
			assign x21_out      = a10_wr[672];                 
			assign x22_out      = a10_wr[416];                 
			assign x23_out      = a10_wr[928];                 
			assign x24_out      = a10_wr[96];                  
			assign x25_out      = a10_wr[608];                 
			assign x26_out      = a10_wr[352];                 
			assign x27_out      = a10_wr[864];                 
			assign x28_out      = a10_wr[224];                 
			assign x29_out      = a10_wr[736];                 
			assign x30_out      = a10_wr[480];                 
			assign x31_out      = a10_wr[992];                 
			assign x32_out      = a10_wr[16];                  
			assign x33_out      = a10_wr[528];                 
			assign x34_out      = a10_wr[272];                 
			assign x35_out      = a10_wr[784];                 
			assign x36_out      = a10_wr[144];                 
			assign x37_out      = a10_wr[656];                 
			assign x38_out      = a10_wr[400];                 
			assign x39_out      = a10_wr[912];                 
			assign x40_out      = a10_wr[80];                  
			assign x41_out      = a10_wr[592];                 
			assign x42_out      = a10_wr[336];                 
			assign x43_out      = a10_wr[848];                 
			assign x44_out      = a10_wr[208];                 
			assign x45_out      = a10_wr[720];                 
			assign x46_out      = a10_wr[464];                 
			assign x47_out      = a10_wr[976];                 
			assign x48_out      = a10_wr[48];                  
			assign x49_out      = a10_wr[560];                 
			assign x50_out      = a10_wr[304];                 
			assign x51_out      = a10_wr[816];                 
			assign x52_out      = a10_wr[176];                 
			assign x53_out      = a10_wr[688];                 
			assign x54_out      = a10_wr[432];                 
			assign x55_out      = a10_wr[944];                 
			assign x56_out      = a10_wr[112];                 
			assign x57_out      = a10_wr[624];                 
			assign x58_out      = a10_wr[368];                 
			assign x59_out      = a10_wr[880];                 
			assign x60_out      = a10_wr[240];                 
			assign x61_out      = a10_wr[752];                 
			assign x62_out      = a10_wr[496];                 
			assign x63_out      = a10_wr[1008];                
			assign x64_out      = a10_wr[8];                   
			assign x65_out      = a10_wr[520];                 
			assign x66_out      = a10_wr[264];                 
			assign x67_out      = a10_wr[776];                 
			assign x68_out      = a10_wr[136];                 
			assign x69_out      = a10_wr[648];                 
			assign x70_out      = a10_wr[392];                 
			assign x71_out      = a10_wr[904];                 
			assign x72_out      = a10_wr[72];                  
			assign x73_out      = a10_wr[584];                 
			assign x74_out      = a10_wr[328];                 
			assign x75_out      = a10_wr[840];                 
			assign x76_out      = a10_wr[200];                 
			assign x77_out      = a10_wr[712];                 
			assign x78_out      = a10_wr[456];                 
			assign x79_out      = a10_wr[968];                 
			assign x80_out      = a10_wr[40];                  
			assign x81_out      = a10_wr[552];                 
			assign x82_out      = a10_wr[296];                 
			assign x83_out      = a10_wr[808];                 
			assign x84_out      = a10_wr[168];                 
			assign x85_out      = a10_wr[680];                 
			assign x86_out      = a10_wr[424];                 
			assign x87_out      = a10_wr[936];                 
			assign x88_out      = a10_wr[104];                 
			assign x89_out      = a10_wr[616];                 
			assign x90_out      = a10_wr[360];                 
			assign x91_out      = a10_wr[872];                 
			assign x92_out      = a10_wr[232];                 
			assign x93_out      = a10_wr[744];                 
			assign x94_out      = a10_wr[488];                 
			assign x95_out      = a10_wr[1000];                
			assign x96_out      = a10_wr[24];                  
			assign x97_out      = a10_wr[536];                 
			assign x98_out      = a10_wr[280];                 
			assign x99_out      = a10_wr[792];                 
			assign x100_out     = a10_wr[152];                 
			assign x101_out     = a10_wr[664];                 
			assign x102_out     = a10_wr[408];                 
			assign x103_out     = a10_wr[920];                 
			assign x104_out     = a10_wr[88];                  
			assign x105_out     = a10_wr[600];                 
			assign x106_out     = a10_wr[344];                 
			assign x107_out     = a10_wr[856];                 
			assign x108_out     = a10_wr[216];                 
			assign x109_out     = a10_wr[728];                 
			assign x110_out     = a10_wr[472];                 
			assign x111_out     = a10_wr[984];                 
			assign x112_out     = a10_wr[56];                  
			assign x113_out     = a10_wr[568];                 
			assign x114_out     = a10_wr[312];                 
			assign x115_out     = a10_wr[824];                 
			assign x116_out     = a10_wr[184];                 
			assign x117_out     = a10_wr[696];                 
			assign x118_out     = a10_wr[440];                 
			assign x119_out     = a10_wr[952];                 
			assign x120_out     = a10_wr[120];                 
			assign x121_out     = a10_wr[632];                 
			assign x122_out     = a10_wr[376];                 
			assign x123_out     = a10_wr[888];                 
			assign x124_out     = a10_wr[248];                 
			assign x125_out     = a10_wr[760];                 
			assign x126_out     = a10_wr[504];                 
			assign x127_out     = a10_wr[1016];                
			assign x128_out     = a10_wr[4];                   
			assign x129_out     = a10_wr[516];                 
			assign x130_out     = a10_wr[260];                 
			assign x131_out     = a10_wr[772];                 
			assign x132_out     = a10_wr[132];                 
			assign x133_out     = a10_wr[644];                 
			assign x134_out     = a10_wr[388];                 
			assign x135_out     = a10_wr[900];                 
			assign x136_out     = a10_wr[68];                  
			assign x137_out     = a10_wr[580];                 
			assign x138_out     = a10_wr[324];                 
			assign x139_out     = a10_wr[836];                 
			assign x140_out     = a10_wr[196];                 
			assign x141_out     = a10_wr[708];                 
			assign x142_out     = a10_wr[452];                 
			assign x143_out     = a10_wr[964];                 
			assign x144_out     = a10_wr[36];                  
			assign x145_out     = a10_wr[548];                 
			assign x146_out     = a10_wr[292];                 
			assign x147_out     = a10_wr[804];                 
			assign x148_out     = a10_wr[164];                 
			assign x149_out     = a10_wr[676];                 
			assign x150_out     = a10_wr[420];                 
			assign x151_out     = a10_wr[932];                 
			assign x152_out     = a10_wr[100];                 
			assign x153_out     = a10_wr[612];                 
			assign x154_out     = a10_wr[356];                 
			assign x155_out     = a10_wr[868];                 
			assign x156_out     = a10_wr[228];                 
			assign x157_out     = a10_wr[740];                 
			assign x158_out     = a10_wr[484];                 
			assign x159_out     = a10_wr[996];                 
			assign x160_out     = a10_wr[20];                  
			assign x161_out     = a10_wr[532];                 
			assign x162_out     = a10_wr[276];                 
			assign x163_out     = a10_wr[788];                 
			assign x164_out     = a10_wr[148];                 
			assign x165_out     = a10_wr[660];                 
			assign x166_out     = a10_wr[404];                 
			assign x167_out     = a10_wr[916];                 
			assign x168_out     = a10_wr[84];                  
			assign x169_out     = a10_wr[596];                 
			assign x170_out     = a10_wr[340];                 
			assign x171_out     = a10_wr[852];                 
			assign x172_out     = a10_wr[212];                 
			assign x173_out     = a10_wr[724];                 
			assign x174_out     = a10_wr[468];                 
			assign x175_out     = a10_wr[980];                 
			assign x176_out     = a10_wr[52];                  
			assign x177_out     = a10_wr[564];                 
			assign x178_out     = a10_wr[308];                 
			assign x179_out     = a10_wr[820];                 
			assign x180_out     = a10_wr[180];                 
			assign x181_out     = a10_wr[692];                 
			assign x182_out     = a10_wr[436];                 
			assign x183_out     = a10_wr[948];                 
			assign x184_out     = a10_wr[116];                 
			assign x185_out     = a10_wr[628];                 
			assign x186_out     = a10_wr[372];                 
			assign x187_out     = a10_wr[884];                 
			assign x188_out     = a10_wr[244];                 
			assign x189_out     = a10_wr[756];                 
			assign x190_out     = a10_wr[500];                 
			assign x191_out     = a10_wr[1012];                
			assign x192_out     = a10_wr[12];                  
			assign x193_out     = a10_wr[524];                 
			assign x194_out     = a10_wr[268];                 
			assign x195_out     = a10_wr[780];                 
			assign x196_out     = a10_wr[140];                 
			assign x197_out     = a10_wr[652];                 
			assign x198_out     = a10_wr[396];                 
			assign x199_out     = a10_wr[908];                 
			assign x200_out     = a10_wr[76];                  
			assign x201_out     = a10_wr[588];                 
			assign x202_out     = a10_wr[332];                 
			assign x203_out     = a10_wr[844];                 
			assign x204_out     = a10_wr[204];                 
			assign x205_out     = a10_wr[716];                 
			assign x206_out     = a10_wr[460];                 
			assign x207_out     = a10_wr[972];                 
			assign x208_out     = a10_wr[44];                  
			assign x209_out     = a10_wr[556];                 
			assign x210_out     = a10_wr[300];                 
			assign x211_out     = a10_wr[812];                 
			assign x212_out     = a10_wr[172];                 
			assign x213_out     = a10_wr[684];                 
			assign x214_out     = a10_wr[428];                 
			assign x215_out     = a10_wr[940];                 
			assign x216_out     = a10_wr[108];                 
			assign x217_out     = a10_wr[620];                 
			assign x218_out     = a10_wr[364];                 
			assign x219_out     = a10_wr[876];                 
			assign x220_out     = a10_wr[236];                 
			assign x221_out     = a10_wr[748];                 
			assign x222_out     = a10_wr[492];                 
			assign x223_out     = a10_wr[1004];                
			assign x224_out     = a10_wr[28];                  
			assign x225_out     = a10_wr[540];                 
			assign x226_out     = a10_wr[284];                 
			assign x227_out     = a10_wr[796];                 
			assign x228_out     = a10_wr[156];                 
			assign x229_out     = a10_wr[668];                 
			assign x230_out     = a10_wr[412];                 
			assign x231_out     = a10_wr[924];                 
			assign x232_out     = a10_wr[92];                  
			assign x233_out     = a10_wr[604];                 
			assign x234_out     = a10_wr[348];                 
			assign x235_out     = a10_wr[860];                 
			assign x236_out     = a10_wr[220];                 
			assign x237_out     = a10_wr[732];                 
			assign x238_out     = a10_wr[476];                 
			assign x239_out     = a10_wr[988];                 
			assign x240_out     = a10_wr[60];                  
			assign x241_out     = a10_wr[572];                 
			assign x242_out     = a10_wr[316];                 
			assign x243_out     = a10_wr[828];                 
			assign x244_out     = a10_wr[188];                 
			assign x245_out     = a10_wr[700];                 
			assign x246_out     = a10_wr[444];                 
			assign x247_out     = a10_wr[956];                 
			assign x248_out     = a10_wr[124];                 
			assign x249_out     = a10_wr[636];                 
			assign x250_out     = a10_wr[380];                 
			assign x251_out     = a10_wr[892];                 
			assign x252_out     = a10_wr[252];                 
			assign x253_out     = a10_wr[764];                 
			assign x254_out     = a10_wr[508];                 
			assign x255_out     = a10_wr[1020];                
			assign x256_out     = a10_wr[2];                   
			assign x257_out     = a10_wr[514];                 
			assign x258_out     = a10_wr[258];                 
			assign x259_out     = a10_wr[770];                 
			assign x260_out     = a10_wr[130];                 
			assign x261_out     = a10_wr[642];                 
			assign x262_out     = a10_wr[386];                 
			assign x263_out     = a10_wr[898];                 
			assign x264_out     = a10_wr[66];                  
			assign x265_out     = a10_wr[578];                 
			assign x266_out     = a10_wr[322];                 
			assign x267_out     = a10_wr[834];                 
			assign x268_out     = a10_wr[194];                 
			assign x269_out     = a10_wr[706];                 
			assign x270_out     = a10_wr[450];                 
			assign x271_out     = a10_wr[962];                 
			assign x272_out     = a10_wr[34];                  
			assign x273_out     = a10_wr[546];                 
			assign x274_out     = a10_wr[290];                 
			assign x275_out     = a10_wr[802];                 
			assign x276_out     = a10_wr[162];                 
			assign x277_out     = a10_wr[674];                 
			assign x278_out     = a10_wr[418];                 
			assign x279_out     = a10_wr[930];                 
			assign x280_out     = a10_wr[98];                  
			assign x281_out     = a10_wr[610];                 
			assign x282_out     = a10_wr[354];                 
			assign x283_out     = a10_wr[866];                 
			assign x284_out     = a10_wr[226];                 
			assign x285_out     = a10_wr[738];                 
			assign x286_out     = a10_wr[482];                 
			assign x287_out     = a10_wr[994];                 
			assign x288_out     = a10_wr[18];                  
			assign x289_out     = a10_wr[530];                 
			assign x290_out     = a10_wr[274];                 
			assign x291_out     = a10_wr[786];                 
			assign x292_out     = a10_wr[146];                 
			assign x293_out     = a10_wr[658];                 
			assign x294_out     = a10_wr[402];                 
			assign x295_out     = a10_wr[914];                 
			assign x296_out     = a10_wr[82];                  
			assign x297_out     = a10_wr[594];                 
			assign x298_out     = a10_wr[338];                 
			assign x299_out     = a10_wr[850];                 
			assign x300_out     = a10_wr[210];                 
			assign x301_out     = a10_wr[722];                 
			assign x302_out     = a10_wr[466];                 
			assign x303_out     = a10_wr[978];                 
			assign x304_out     = a10_wr[50];                  
			assign x305_out     = a10_wr[562];                 
			assign x306_out     = a10_wr[306];                 
			assign x307_out     = a10_wr[818];                 
			assign x308_out     = a10_wr[178];                 
			assign x309_out     = a10_wr[690];                 
			assign x310_out     = a10_wr[434];                 
			assign x311_out     = a10_wr[946];                 
			assign x312_out     = a10_wr[114];                 
			assign x313_out     = a10_wr[626];                 
			assign x314_out     = a10_wr[370];                 
			assign x315_out     = a10_wr[882];                 
			assign x316_out     = a10_wr[242];                 
			assign x317_out     = a10_wr[754];                 
			assign x318_out     = a10_wr[498];                 
			assign x319_out     = a10_wr[1010];                
			assign x320_out     = a10_wr[10];                  
			assign x321_out     = a10_wr[522];                 
			assign x322_out     = a10_wr[266];                 
			assign x323_out     = a10_wr[778];                 
			assign x324_out     = a10_wr[138];                 
			assign x325_out     = a10_wr[650];                 
			assign x326_out     = a10_wr[394];                 
			assign x327_out     = a10_wr[906];                 
			assign x328_out     = a10_wr[74];                  
			assign x329_out     = a10_wr[586];                 
			assign x330_out     = a10_wr[330];                 
			assign x331_out     = a10_wr[842];                 
			assign x332_out     = a10_wr[202];                 
			assign x333_out     = a10_wr[714];                 
			assign x334_out     = a10_wr[458];                 
			assign x335_out     = a10_wr[970];                 
			assign x336_out     = a10_wr[42];                  
			assign x337_out     = a10_wr[554];                 
			assign x338_out     = a10_wr[298];                 
			assign x339_out     = a10_wr[810];                 
			assign x340_out     = a10_wr[170];                 
			assign x341_out     = a10_wr[682];                 
			assign x342_out     = a10_wr[426];                 
			assign x343_out     = a10_wr[938];                 
			assign x344_out     = a10_wr[106];                 
			assign x345_out     = a10_wr[618];                 
			assign x346_out     = a10_wr[362];                 
			assign x347_out     = a10_wr[874];                 
			assign x348_out     = a10_wr[234];                 
			assign x349_out     = a10_wr[746];                 
			assign x350_out     = a10_wr[490];                 
			assign x351_out     = a10_wr[1002];                
			assign x352_out     = a10_wr[26];                  
			assign x353_out     = a10_wr[538];                 
			assign x354_out     = a10_wr[282];                 
			assign x355_out     = a10_wr[794];                 
			assign x356_out     = a10_wr[154];                 
			assign x357_out     = a10_wr[666];                 
			assign x358_out     = a10_wr[410];                 
			assign x359_out     = a10_wr[922];                 
			assign x360_out     = a10_wr[90];                  
			assign x361_out     = a10_wr[602];                 
			assign x362_out     = a10_wr[346];                 
			assign x363_out     = a10_wr[858];                 
			assign x364_out     = a10_wr[218];                 
			assign x365_out     = a10_wr[730];                 
			assign x366_out     = a10_wr[474];                 
			assign x367_out     = a10_wr[986];                 
			assign x368_out     = a10_wr[58];                  
			assign x369_out     = a10_wr[570];                 
			assign x370_out     = a10_wr[314];                 
			assign x371_out     = a10_wr[826];                 
			assign x372_out     = a10_wr[186];                 
			assign x373_out     = a10_wr[698];                 
			assign x374_out     = a10_wr[442];                 
			assign x375_out     = a10_wr[954];                 
			assign x376_out     = a10_wr[122];                 
			assign x377_out     = a10_wr[634];                 
			assign x378_out     = a10_wr[378];                 
			assign x379_out     = a10_wr[890];                 
			assign x380_out     = a10_wr[250];                 
			assign x381_out     = a10_wr[762];                 
			assign x382_out     = a10_wr[506];                 
			assign x383_out     = a10_wr[1018];                
			assign x384_out     = a10_wr[6];                   
			assign x385_out     = a10_wr[518];                 
			assign x386_out     = a10_wr[262];                 
			assign x387_out     = a10_wr[774];                 
			assign x388_out     = a10_wr[134];                 
			assign x389_out     = a10_wr[646];                 
			assign x390_out     = a10_wr[390];                 
			assign x391_out     = a10_wr[902];                 
			assign x392_out     = a10_wr[70];                  
			assign x393_out     = a10_wr[582];                 
			assign x394_out     = a10_wr[326];                 
			assign x395_out     = a10_wr[838];                 
			assign x396_out     = a10_wr[198];                 
			assign x397_out     = a10_wr[710];                 
			assign x398_out     = a10_wr[454];                 
			assign x399_out     = a10_wr[966];                 
			assign x400_out     = a10_wr[38];                  
			assign x401_out     = a10_wr[550];                 
			assign x402_out     = a10_wr[294];                 
			assign x403_out     = a10_wr[806];                 
			assign x404_out     = a10_wr[166];                 
			assign x405_out     = a10_wr[678];                 
			assign x406_out     = a10_wr[422];                 
			assign x407_out     = a10_wr[934];                 
			assign x408_out     = a10_wr[102];                 
			assign x409_out     = a10_wr[614];                 
			assign x410_out     = a10_wr[358];                 
			assign x411_out     = a10_wr[870];                 
			assign x412_out     = a10_wr[230];                 
			assign x413_out     = a10_wr[742];                 
			assign x414_out     = a10_wr[486];                 
			assign x415_out     = a10_wr[998];                 
			assign x416_out     = a10_wr[22];                  
			assign x417_out     = a10_wr[534];                 
			assign x418_out     = a10_wr[278];                 
			assign x419_out     = a10_wr[790];                 
			assign x420_out     = a10_wr[150];                 
			assign x421_out     = a10_wr[662];                 
			assign x422_out     = a10_wr[406];                 
			assign x423_out     = a10_wr[918];                 
			assign x424_out     = a10_wr[86];                  
			assign x425_out     = a10_wr[598];                 
			assign x426_out     = a10_wr[342];                 
			assign x427_out     = a10_wr[854];                 
			assign x428_out     = a10_wr[214];                 
			assign x429_out     = a10_wr[726];                 
			assign x430_out     = a10_wr[470];                 
			assign x431_out     = a10_wr[982];                 
			assign x432_out     = a10_wr[54];                  
			assign x433_out     = a10_wr[566];                 
			assign x434_out     = a10_wr[310];                 
			assign x435_out     = a10_wr[822];                 
			assign x436_out     = a10_wr[182];                 
			assign x437_out     = a10_wr[694];                 
			assign x438_out     = a10_wr[438];                 
			assign x439_out     = a10_wr[950];                 
			assign x440_out     = a10_wr[118];                 
			assign x441_out     = a10_wr[630];                 
			assign x442_out     = a10_wr[374];                 
			assign x443_out     = a10_wr[886];                 
			assign x444_out     = a10_wr[246];                 
			assign x445_out     = a10_wr[758];                 
			assign x446_out     = a10_wr[502];                 
			assign x447_out     = a10_wr[1014];                
			assign x448_out     = a10_wr[14];                  
			assign x449_out     = a10_wr[526];                 
			assign x450_out     = a10_wr[270];                 
			assign x451_out     = a10_wr[782];                 
			assign x452_out     = a10_wr[142];                 
			assign x453_out     = a10_wr[654];                 
			assign x454_out     = a10_wr[398];                 
			assign x455_out     = a10_wr[910];                 
			assign x456_out     = a10_wr[78];                  
			assign x457_out     = a10_wr[590];                 
			assign x458_out     = a10_wr[334];                 
			assign x459_out     = a10_wr[846];                 
			assign x460_out     = a10_wr[206];                 
			assign x461_out     = a10_wr[718];                 
			assign x462_out     = a10_wr[462];                 
			assign x463_out     = a10_wr[974];                 
			assign x464_out     = a10_wr[46];                  
			assign x465_out     = a10_wr[558];                 
			assign x466_out     = a10_wr[302];                 
			assign x467_out     = a10_wr[814];                 
			assign x468_out     = a10_wr[174];                 
			assign x469_out     = a10_wr[686];                 
			assign x470_out     = a10_wr[430];                 
			assign x471_out     = a10_wr[942];                 
			assign x472_out     = a10_wr[110];                 
			assign x473_out     = a10_wr[622];                 
			assign x474_out     = a10_wr[366];                 
			assign x475_out     = a10_wr[878];                 
			assign x476_out     = a10_wr[238];                 
			assign x477_out     = a10_wr[750];                 
			assign x478_out     = a10_wr[494];                 
			assign x479_out     = a10_wr[1006];                
			assign x480_out     = a10_wr[30];                  
			assign x481_out     = a10_wr[542];                 
			assign x482_out     = a10_wr[286];                 
			assign x483_out     = a10_wr[798];                 
			assign x484_out     = a10_wr[158];                 
			assign x485_out     = a10_wr[670];                 
			assign x486_out     = a10_wr[414];                 
			assign x487_out     = a10_wr[926];                 
			assign x488_out     = a10_wr[94];                  
			assign x489_out     = a10_wr[606];                 
			assign x490_out     = a10_wr[350];                 
			assign x491_out     = a10_wr[862];                 
			assign x492_out     = a10_wr[222];                 
			assign x493_out     = a10_wr[734];                 
			assign x494_out     = a10_wr[478];                 
			assign x495_out     = a10_wr[990];                 
			assign x496_out     = a10_wr[62];                  
			assign x497_out     = a10_wr[574];                 
			assign x498_out     = a10_wr[318];                 
			assign x499_out     = a10_wr[830];                 
			assign x500_out     = a10_wr[190];                 
			assign x501_out     = a10_wr[702];                 
			assign x502_out     = a10_wr[446];                 
			assign x503_out     = a10_wr[958];                 
			assign x504_out     = a10_wr[126];                 
			assign x505_out     = a10_wr[638];                 
			assign x506_out     = a10_wr[382];                 
			assign x507_out     = a10_wr[894];                 
			assign x508_out     = a10_wr[254];                 
			assign x509_out     = a10_wr[766];                 
			assign x510_out     = a10_wr[510];                 
			assign x511_out     = a10_wr[1022];                
			assign x512_out     = a10_wr[1];                   
			assign x513_out     = a10_wr[513];                 
			assign x514_out     = a10_wr[257];                 
			assign x515_out     = a10_wr[769];                 
			assign x516_out     = a10_wr[129];                 
			assign x517_out     = a10_wr[641];                 
			assign x518_out     = a10_wr[385];                 
			assign x519_out     = a10_wr[897];                 
			assign x520_out     = a10_wr[65];                  
			assign x521_out     = a10_wr[577];                 
			assign x522_out     = a10_wr[321];                 
			assign x523_out     = a10_wr[833];                 
			assign x524_out     = a10_wr[193];                 
			assign x525_out     = a10_wr[705];                 
			assign x526_out     = a10_wr[449];                 
			assign x527_out     = a10_wr[961];                 
			assign x528_out     = a10_wr[33];                  
			assign x529_out     = a10_wr[545];                 
			assign x530_out     = a10_wr[289];                 
			assign x531_out     = a10_wr[801];                 
			assign x532_out     = a10_wr[161];                 
			assign x533_out     = a10_wr[673];                 
			assign x534_out     = a10_wr[417];                 
			assign x535_out     = a10_wr[929];                 
			assign x536_out     = a10_wr[97];                  
			assign x537_out     = a10_wr[609];                 
			assign x538_out     = a10_wr[353];                 
			assign x539_out     = a10_wr[865];                 
			assign x540_out     = a10_wr[225];                 
			assign x541_out     = a10_wr[737];                 
			assign x542_out     = a10_wr[481];                 
			assign x543_out     = a10_wr[993];                 
			assign x544_out     = a10_wr[17];                  
			assign x545_out     = a10_wr[529];                 
			assign x546_out     = a10_wr[273];                 
			assign x547_out     = a10_wr[785];                 
			assign x548_out     = a10_wr[145];                 
			assign x549_out     = a10_wr[657];                 
			assign x550_out     = a10_wr[401];                 
			assign x551_out     = a10_wr[913];                 
			assign x552_out     = a10_wr[81];                  
			assign x553_out     = a10_wr[593];                 
			assign x554_out     = a10_wr[337];                 
			assign x555_out     = a10_wr[849];                 
			assign x556_out     = a10_wr[209];                 
			assign x557_out     = a10_wr[721];                 
			assign x558_out     = a10_wr[465];                 
			assign x559_out     = a10_wr[977];                 
			assign x560_out     = a10_wr[49];                  
			assign x561_out     = a10_wr[561];                 
			assign x562_out     = a10_wr[305];                 
			assign x563_out     = a10_wr[817];                 
			assign x564_out     = a10_wr[177];                 
			assign x565_out     = a10_wr[689];                 
			assign x566_out     = a10_wr[433];                 
			assign x567_out     = a10_wr[945];                 
			assign x568_out     = a10_wr[113];                 
			assign x569_out     = a10_wr[625];                 
			assign x570_out     = a10_wr[369];                 
			assign x571_out     = a10_wr[881];                 
			assign x572_out     = a10_wr[241];                 
			assign x573_out     = a10_wr[753];                 
			assign x574_out     = a10_wr[497];                 
			assign x575_out     = a10_wr[1009];                
			assign x576_out     = a10_wr[9];                   
			assign x577_out     = a10_wr[521];                 
			assign x578_out     = a10_wr[265];                 
			assign x579_out     = a10_wr[777];                 
			assign x580_out     = a10_wr[137];                 
			assign x581_out     = a10_wr[649];                 
			assign x582_out     = a10_wr[393];                 
			assign x583_out     = a10_wr[905];                 
			assign x584_out     = a10_wr[73];                  
			assign x585_out     = a10_wr[585];                 
			assign x586_out     = a10_wr[329];                 
			assign x587_out     = a10_wr[841];                 
			assign x588_out     = a10_wr[201];                 
			assign x589_out     = a10_wr[713];                 
			assign x590_out     = a10_wr[457];                 
			assign x591_out     = a10_wr[969];                 
			assign x592_out     = a10_wr[41];                  
			assign x593_out     = a10_wr[553];                 
			assign x594_out     = a10_wr[297];                 
			assign x595_out     = a10_wr[809];                 
			assign x596_out     = a10_wr[169];                 
			assign x597_out     = a10_wr[681];                 
			assign x598_out     = a10_wr[425];                 
			assign x599_out     = a10_wr[937];                 
			assign x600_out     = a10_wr[105];                 
			assign x601_out     = a10_wr[617];                 
			assign x602_out     = a10_wr[361];                 
			assign x603_out     = a10_wr[873];                 
			assign x604_out     = a10_wr[233];                 
			assign x605_out     = a10_wr[745];                 
			assign x606_out     = a10_wr[489];                 
			assign x607_out     = a10_wr[1001];                
			assign x608_out     = a10_wr[25];                  
			assign x609_out     = a10_wr[537];                 
			assign x610_out     = a10_wr[281];                 
			assign x611_out     = a10_wr[793];                 
			assign x612_out     = a10_wr[153];                 
			assign x613_out     = a10_wr[665];                 
			assign x614_out     = a10_wr[409];                 
			assign x615_out     = a10_wr[921];                 
			assign x616_out     = a10_wr[89];                  
			assign x617_out     = a10_wr[601];                 
			assign x618_out     = a10_wr[345];                 
			assign x619_out     = a10_wr[857];                 
			assign x620_out     = a10_wr[217];                 
			assign x621_out     = a10_wr[729];                 
			assign x622_out     = a10_wr[473];                 
			assign x623_out     = a10_wr[985];                 
			assign x624_out     = a10_wr[57];                  
			assign x625_out     = a10_wr[569];                 
			assign x626_out     = a10_wr[313];                 
			assign x627_out     = a10_wr[825];                 
			assign x628_out     = a10_wr[185];                 
			assign x629_out     = a10_wr[697];                 
			assign x630_out     = a10_wr[441];                 
			assign x631_out     = a10_wr[953];                 
			assign x632_out     = a10_wr[121];                 
			assign x633_out     = a10_wr[633];                 
			assign x634_out     = a10_wr[377];                 
			assign x635_out     = a10_wr[889];                 
			assign x636_out     = a10_wr[249];                 
			assign x637_out     = a10_wr[761];                 
			assign x638_out     = a10_wr[505];                 
			assign x639_out     = a10_wr[1017];                
			assign x640_out     = a10_wr[5];                   
			assign x641_out     = a10_wr[517];                 
			assign x642_out     = a10_wr[261];                 
			assign x643_out     = a10_wr[773];                 
			assign x644_out     = a10_wr[133];                 
			assign x645_out     = a10_wr[645];                 
			assign x646_out     = a10_wr[389];                 
			assign x647_out     = a10_wr[901];                 
			assign x648_out     = a10_wr[69];                  
			assign x649_out     = a10_wr[581];                 
			assign x650_out     = a10_wr[325];                 
			assign x651_out     = a10_wr[837];                 
			assign x652_out     = a10_wr[197];                 
			assign x653_out     = a10_wr[709];                 
			assign x654_out     = a10_wr[453];                 
			assign x655_out     = a10_wr[965];                 
			assign x656_out     = a10_wr[37];                  
			assign x657_out     = a10_wr[549];                 
			assign x658_out     = a10_wr[293];                 
			assign x659_out     = a10_wr[805];                 
			assign x660_out     = a10_wr[165];                 
			assign x661_out     = a10_wr[677];                 
			assign x662_out     = a10_wr[421];                 
			assign x663_out     = a10_wr[933];                 
			assign x664_out     = a10_wr[101];                 
			assign x665_out     = a10_wr[613];                 
			assign x666_out     = a10_wr[357];                 
			assign x667_out     = a10_wr[869];                 
			assign x668_out     = a10_wr[229];                 
			assign x669_out     = a10_wr[741];                 
			assign x670_out     = a10_wr[485];                 
			assign x671_out     = a10_wr[997];                 
			assign x672_out     = a10_wr[21];                  
			assign x673_out     = a10_wr[533];                 
			assign x674_out     = a10_wr[277];                 
			assign x675_out     = a10_wr[789];                 
			assign x676_out     = a10_wr[149];                 
			assign x677_out     = a10_wr[661];                 
			assign x678_out     = a10_wr[405];                 
			assign x679_out     = a10_wr[917];                 
			assign x680_out     = a10_wr[85];                  
			assign x681_out     = a10_wr[597];                 
			assign x682_out     = a10_wr[341];                 
			assign x683_out     = a10_wr[853];                 
			assign x684_out     = a10_wr[213];                 
			assign x685_out     = a10_wr[725];                 
			assign x686_out     = a10_wr[469];                 
			assign x687_out     = a10_wr[981];                 
			assign x688_out     = a10_wr[53];                  
			assign x689_out     = a10_wr[565];                 
			assign x690_out     = a10_wr[309];                 
			assign x691_out     = a10_wr[821];                 
			assign x692_out     = a10_wr[181];                 
			assign x693_out     = a10_wr[693];                 
			assign x694_out     = a10_wr[437];                 
			assign x695_out     = a10_wr[949];                 
			assign x696_out     = a10_wr[117];                 
			assign x697_out     = a10_wr[629];                 
			assign x698_out     = a10_wr[373];                 
			assign x699_out     = a10_wr[885];                 
			assign x700_out     = a10_wr[245];                 
			assign x701_out     = a10_wr[757];                 
			assign x702_out     = a10_wr[501];                 
			assign x703_out     = a10_wr[1013];                
			assign x704_out     = a10_wr[13];                  
			assign x705_out     = a10_wr[525];                 
			assign x706_out     = a10_wr[269];                 
			assign x707_out     = a10_wr[781];                 
			assign x708_out     = a10_wr[141];                 
			assign x709_out     = a10_wr[653];                 
			assign x710_out     = a10_wr[397];                 
			assign x711_out     = a10_wr[909];                 
			assign x712_out     = a10_wr[77];                  
			assign x713_out     = a10_wr[589];                 
			assign x714_out     = a10_wr[333];                 
			assign x715_out     = a10_wr[845];                 
			assign x716_out     = a10_wr[205];                 
			assign x717_out     = a10_wr[717];                 
			assign x718_out     = a10_wr[461];                 
			assign x719_out     = a10_wr[973];                 
			assign x720_out     = a10_wr[45];                  
			assign x721_out     = a10_wr[557];                 
			assign x722_out     = a10_wr[301];                 
			assign x723_out     = a10_wr[813];                 
			assign x724_out     = a10_wr[173];                 
			assign x725_out     = a10_wr[685];                 
			assign x726_out     = a10_wr[429];                 
			assign x727_out     = a10_wr[941];                 
			assign x728_out     = a10_wr[109];                 
			assign x729_out     = a10_wr[621];                 
			assign x730_out     = a10_wr[365];                 
			assign x731_out     = a10_wr[877];                 
			assign x732_out     = a10_wr[237];                 
			assign x733_out     = a10_wr[749];                 
			assign x734_out     = a10_wr[493];                 
			assign x735_out     = a10_wr[1005];                
			assign x736_out     = a10_wr[29];                  
			assign x737_out     = a10_wr[541];                 
			assign x738_out     = a10_wr[285];                 
			assign x739_out     = a10_wr[797];                 
			assign x740_out     = a10_wr[157];                 
			assign x741_out     = a10_wr[669];                 
			assign x742_out     = a10_wr[413];                 
			assign x743_out     = a10_wr[925];                 
			assign x744_out     = a10_wr[93];                  
			assign x745_out     = a10_wr[605];                 
			assign x746_out     = a10_wr[349];                 
			assign x747_out     = a10_wr[861];                 
			assign x748_out     = a10_wr[221];                 
			assign x749_out     = a10_wr[733];                 
			assign x750_out     = a10_wr[477];                 
			assign x751_out     = a10_wr[989];                 
			assign x752_out     = a10_wr[61];                  
			assign x753_out     = a10_wr[573];                 
			assign x754_out     = a10_wr[317];                 
			assign x755_out     = a10_wr[829];                 
			assign x756_out     = a10_wr[189];                 
			assign x757_out     = a10_wr[701];                 
			assign x758_out     = a10_wr[445];                 
			assign x759_out     = a10_wr[957];                 
			assign x760_out     = a10_wr[125];                 
			assign x761_out     = a10_wr[637];                 
			assign x762_out     = a10_wr[381];                 
			assign x763_out     = a10_wr[893];                 
			assign x764_out     = a10_wr[253];                 
			assign x765_out     = a10_wr[765];                 
			assign x766_out     = a10_wr[509];                 
			assign x767_out     = a10_wr[1021];                
			assign x768_out     = a10_wr[3];                   
			assign x769_out     = a10_wr[515];                 
			assign x770_out     = a10_wr[259];                 
			assign x771_out     = a10_wr[771];                 
			assign x772_out     = a10_wr[131];                 
			assign x773_out     = a10_wr[643];                 
			assign x774_out     = a10_wr[387];                 
			assign x775_out     = a10_wr[899];                 
			assign x776_out     = a10_wr[67];                  
			assign x777_out     = a10_wr[579];                 
			assign x778_out     = a10_wr[323];                 
			assign x779_out     = a10_wr[835];                 
			assign x780_out     = a10_wr[195];                 
			assign x781_out     = a10_wr[707];                 
			assign x782_out     = a10_wr[451];                 
			assign x783_out     = a10_wr[963];                 
			assign x784_out     = a10_wr[35];                  
			assign x785_out     = a10_wr[547];                 
			assign x786_out     = a10_wr[291];                 
			assign x787_out     = a10_wr[803];                 
			assign x788_out     = a10_wr[163];                 
			assign x789_out     = a10_wr[675];                 
			assign x790_out     = a10_wr[419];                 
			assign x791_out     = a10_wr[931];                 
			assign x792_out     = a10_wr[99];                  
			assign x793_out     = a10_wr[611];                 
			assign x794_out     = a10_wr[355];                 
			assign x795_out     = a10_wr[867];                 
			assign x796_out     = a10_wr[227];                 
			assign x797_out     = a10_wr[739];                 
			assign x798_out     = a10_wr[483];                 
			assign x799_out     = a10_wr[995];                 
			assign x800_out     = a10_wr[19];                  
			assign x801_out     = a10_wr[531];                 
			assign x802_out     = a10_wr[275];                 
			assign x803_out     = a10_wr[787];                 
			assign x804_out     = a10_wr[147];                 
			assign x805_out     = a10_wr[659];                 
			assign x806_out     = a10_wr[403];                 
			assign x807_out     = a10_wr[915];                 
			assign x808_out     = a10_wr[83];                  
			assign x809_out     = a10_wr[595];                 
			assign x810_out     = a10_wr[339];                 
			assign x811_out     = a10_wr[851];                 
			assign x812_out     = a10_wr[211];                 
			assign x813_out     = a10_wr[723];                 
			assign x814_out     = a10_wr[467];                 
			assign x815_out     = a10_wr[979];                 
			assign x816_out     = a10_wr[51];                  
			assign x817_out     = a10_wr[563];                 
			assign x818_out     = a10_wr[307];                 
			assign x819_out     = a10_wr[819];                 
			assign x820_out     = a10_wr[179];                 
			assign x821_out     = a10_wr[691];                 
			assign x822_out     = a10_wr[435];                 
			assign x823_out     = a10_wr[947];                 
			assign x824_out     = a10_wr[115];                 
			assign x825_out     = a10_wr[627];                 
			assign x826_out     = a10_wr[371];                 
			assign x827_out     = a10_wr[883];                 
			assign x828_out     = a10_wr[243];                 
			assign x829_out     = a10_wr[755];                 
			assign x830_out     = a10_wr[499];                 
			assign x831_out     = a10_wr[1011];                
			assign x832_out     = a10_wr[11];                  
			assign x833_out     = a10_wr[523];                 
			assign x834_out     = a10_wr[267];                 
			assign x835_out     = a10_wr[779];                 
			assign x836_out     = a10_wr[139];                 
			assign x837_out     = a10_wr[651];                 
			assign x838_out     = a10_wr[395];                 
			assign x839_out     = a10_wr[907];                 
			assign x840_out     = a10_wr[75];                  
			assign x841_out     = a10_wr[587];                 
			assign x842_out     = a10_wr[331];                 
			assign x843_out     = a10_wr[843];                 
			assign x844_out     = a10_wr[203];                 
			assign x845_out     = a10_wr[715];                 
			assign x846_out     = a10_wr[459];                 
			assign x847_out     = a10_wr[971];                 
			assign x848_out     = a10_wr[43];                  
			assign x849_out     = a10_wr[555];                 
			assign x850_out     = a10_wr[299];                 
			assign x851_out     = a10_wr[811];                 
			assign x852_out     = a10_wr[171];                 
			assign x853_out     = a10_wr[683];                 
			assign x854_out     = a10_wr[427];                 
			assign x855_out     = a10_wr[939];                 
			assign x856_out     = a10_wr[107];                 
			assign x857_out     = a10_wr[619];                 
			assign x858_out     = a10_wr[363];                 
			assign x859_out     = a10_wr[875];                 
			assign x860_out     = a10_wr[235];                 
			assign x861_out     = a10_wr[747];                 
			assign x862_out     = a10_wr[491];                 
			assign x863_out     = a10_wr[1003];                
			assign x864_out     = a10_wr[27];                  
			assign x865_out     = a10_wr[539];                 
			assign x866_out     = a10_wr[283];                 
			assign x867_out     = a10_wr[795];                 
			assign x868_out     = a10_wr[155];                 
			assign x869_out     = a10_wr[667];                 
			assign x870_out     = a10_wr[411];                 
			assign x871_out     = a10_wr[923];                 
			assign x872_out     = a10_wr[91];                  
			assign x873_out     = a10_wr[603];                 
			assign x874_out     = a10_wr[347];                 
			assign x875_out     = a10_wr[859];                 
			assign x876_out     = a10_wr[219];                 
			assign x877_out     = a10_wr[731];                 
			assign x878_out     = a10_wr[475];                 
			assign x879_out     = a10_wr[987];                 
			assign x880_out     = a10_wr[59];                  
			assign x881_out     = a10_wr[571];                 
			assign x882_out     = a10_wr[315];                 
			assign x883_out     = a10_wr[827];                 
			assign x884_out     = a10_wr[187];                 
			assign x885_out     = a10_wr[699];                 
			assign x886_out     = a10_wr[443];                 
			assign x887_out     = a10_wr[955];                 
			assign x888_out     = a10_wr[123];                 
			assign x889_out     = a10_wr[635];                 
			assign x890_out     = a10_wr[379];                 
			assign x891_out     = a10_wr[891];                 
			assign x892_out     = a10_wr[251];                 
			assign x893_out     = a10_wr[763];                 
			assign x894_out     = a10_wr[507];                 
			assign x895_out     = a10_wr[1019];                
			assign x896_out     = a10_wr[7];                   
			assign x897_out     = a10_wr[519];                 
			assign x898_out     = a10_wr[263];                 
			assign x899_out     = a10_wr[775];                 
			assign x900_out     = a10_wr[135];                 
			assign x901_out     = a10_wr[647];                 
			assign x902_out     = a10_wr[391];                 
			assign x903_out     = a10_wr[903];                 
			assign x904_out     = a10_wr[71];                  
			assign x905_out     = a10_wr[583];                 
			assign x906_out     = a10_wr[327];                 
			assign x907_out     = a10_wr[839];                 
			assign x908_out     = a10_wr[199];                 
			assign x909_out     = a10_wr[711];                 
			assign x910_out     = a10_wr[455];                 
			assign x911_out     = a10_wr[967];                 
			assign x912_out     = a10_wr[39];                  
			assign x913_out     = a10_wr[551];                 
			assign x914_out     = a10_wr[295];                 
			assign x915_out     = a10_wr[807];                 
			assign x916_out     = a10_wr[167];                 
			assign x917_out     = a10_wr[679];                 
			assign x918_out     = a10_wr[423];                 
			assign x919_out     = a10_wr[935];                 
			assign x920_out     = a10_wr[103];                 
			assign x921_out     = a10_wr[615];                 
			assign x922_out     = a10_wr[359];                 
			assign x923_out     = a10_wr[871];                 
			assign x924_out     = a10_wr[231];                 
			assign x925_out     = a10_wr[743];                 
			assign x926_out     = a10_wr[487];                 
			assign x927_out     = a10_wr[999];                 
			assign x928_out     = a10_wr[23];                  
			assign x929_out     = a10_wr[535];                 
			assign x930_out     = a10_wr[279];                 
			assign x931_out     = a10_wr[791];                 
			assign x932_out     = a10_wr[151];                 
			assign x933_out     = a10_wr[663];                 
			assign x934_out     = a10_wr[407];                 
			assign x935_out     = a10_wr[919];                 
			assign x936_out     = a10_wr[87];                  
			assign x937_out     = a10_wr[599];                 
			assign x938_out     = a10_wr[343];                 
			assign x939_out     = a10_wr[855];                 
			assign x940_out     = a10_wr[215];                 
			assign x941_out     = a10_wr[727];                 
			assign x942_out     = a10_wr[471];                 
			assign x943_out     = a10_wr[983];                 
			assign x944_out     = a10_wr[55];                  
			assign x945_out     = a10_wr[567];                 
			assign x946_out     = a10_wr[311];                 
			assign x947_out     = a10_wr[823];                 
			assign x948_out     = a10_wr[183];                 
			assign x949_out     = a10_wr[695];                 
			assign x950_out     = a10_wr[439];                 
			assign x951_out     = a10_wr[951];                 
			assign x952_out     = a10_wr[119];                 
			assign x953_out     = a10_wr[631];                 
			assign x954_out     = a10_wr[375];                 
			assign x955_out     = a10_wr[887];                 
			assign x956_out     = a10_wr[247];                 
			assign x957_out     = a10_wr[759];                 
			assign x958_out     = a10_wr[503];                 
			assign x959_out     = a10_wr[1015];                
			assign x960_out     = a10_wr[15];                  
			assign x961_out     = a10_wr[527];                 
			assign x962_out     = a10_wr[271];                 
			assign x963_out     = a10_wr[783];                 
			assign x964_out     = a10_wr[143];                 
			assign x965_out     = a10_wr[655];                 
			assign x966_out     = a10_wr[399];                 
			assign x967_out     = a10_wr[911];                 
			assign x968_out     = a10_wr[79];                  
			assign x969_out     = a10_wr[591];                 
			assign x970_out     = a10_wr[335];                 
			assign x971_out     = a10_wr[847];                 
			assign x972_out     = a10_wr[207];                 
			assign x973_out     = a10_wr[719];                 
			assign x974_out     = a10_wr[463];                 
			assign x975_out     = a10_wr[975];                 
			assign x976_out     = a10_wr[47];                  
			assign x977_out     = a10_wr[559];                 
			assign x978_out     = a10_wr[303];                 
			assign x979_out     = a10_wr[815];                 
			assign x980_out     = a10_wr[175];                 
			assign x981_out     = a10_wr[687];                 
			assign x982_out     = a10_wr[431];                 
			assign x983_out     = a10_wr[943];                 
			assign x984_out     = a10_wr[111];                 
			assign x985_out     = a10_wr[623];                 
			assign x986_out     = a10_wr[367];                 
			assign x987_out     = a10_wr[879];                 
			assign x988_out     = a10_wr[239];                 
			assign x989_out     = a10_wr[751];                 
			assign x990_out     = a10_wr[495];                 
			assign x991_out     = a10_wr[1007];                
			assign x992_out     = a10_wr[31];                  
			assign x993_out     = a10_wr[543];                 
			assign x994_out     = a10_wr[287];                 
			assign x995_out     = a10_wr[799];                 
			assign x996_out     = a10_wr[159];                 
			assign x997_out     = a10_wr[671];                 
			assign x998_out     = a10_wr[415];                 
			assign x999_out     = a10_wr[927];                 
			assign x1000_out    = a10_wr[95];                  
			assign x1001_out    = a10_wr[607];                 
			assign x1002_out    = a10_wr[351];                 
			assign x1003_out    = a10_wr[863];                 
			assign x1004_out    = a10_wr[223];                 
			assign x1005_out    = a10_wr[735];                 
			assign x1006_out    = a10_wr[479];                 
			assign x1007_out    = a10_wr[991];                 
			assign x1008_out    = a10_wr[63];                  
			assign x1009_out    = a10_wr[575];                 
			assign x1010_out    = a10_wr[319];                 
			assign x1011_out    = a10_wr[831];                 
			assign x1012_out    = a10_wr[191];                 
			assign x1013_out    = a10_wr[703];                 
			assign x1014_out    = a10_wr[447];                 
			assign x1015_out    = a10_wr[959];                 
			assign x1016_out    = a10_wr[127];                 
			assign x1017_out    = a10_wr[639];                 
			assign x1018_out    = a10_wr[383];                 
			assign x1019_out    = a10_wr[895];                 
			assign x1020_out    = a10_wr[255];                 
			assign x1021_out    = a10_wr[767];                 
			assign x1022_out    = a10_wr[511];                 
			assign x1023_out    = a10_wr[1023];                


endmodule
