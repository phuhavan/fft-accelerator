//=====================================================
//
//
//=====================================================
`include "defines.h"
`include "macros.h"

module adderTestBench
#(
	//--- complex data width
		parameter	width 		= 24,
	//--- number of simulation cycle (# inputs)
		parameter simcycle 	= 100000
);
	localparam						hwidth 			= width/2;

	wire							clk, n_rst, n_stall, n_stall_out;
	wire 	signed [31:0]			cur_cycle;

	wire signed [hwidth-1:0] 		dt_in0, dt_in1, dt_in2, dt_in3, dt_in4, dt_in5, dt_in6, dt_in7, dt_in8, dt_in9, dt_in10, dt_in11, dt_in12, dt_in13, dt_in14, dt_in15, 
									dt_in16, dt_in17, dt_in18, dt_in19, dt_in20, dt_in21, dt_in22, dt_in23, dt_in24, dt_in25, dt_in26, dt_in27, dt_in28, dt_in29, dt_in30, dt_in31, 
									dt_in32, dt_in33, dt_in34, dt_in35, dt_in36, dt_in37, dt_in38, dt_in39, dt_in40, dt_in41, dt_in42, dt_in43, dt_in44, dt_in45, dt_in46, dt_in47, 
									dt_in48, dt_in49, dt_in50, dt_in51, dt_in52, dt_in53, dt_in54, dt_in55, dt_in56, dt_in57, dt_in58, dt_in59, dt_in60, dt_in61, dt_in62, dt_in63, 
									dt_in64, dt_in65, dt_in66, dt_in67, dt_in68, dt_in69, dt_in70, dt_in71, dt_in72, dt_in73, dt_in74, dt_in75, dt_in76, dt_in77, dt_in78, dt_in79, 
									dt_in80, dt_in81, dt_in82, dt_in83, dt_in84, dt_in85, dt_in86, dt_in87, dt_in88, dt_in89, dt_in90, dt_in91, dt_in92, dt_in93, dt_in94, dt_in95, 
									dt_in96, dt_in97, dt_in98, dt_in99, dt_in100, dt_in101, dt_in102, dt_in103, dt_in104, dt_in105, dt_in106, dt_in107, dt_in108, dt_in109, dt_in110, dt_in111, 
									dt_in112, dt_in113, dt_in114, dt_in115, dt_in116, dt_in117, dt_in118, dt_in119, dt_in120, dt_in121, dt_in122, dt_in123, dt_in124, dt_in125, dt_in126, dt_in127, 
									dt_in128, dt_in129, dt_in130, dt_in131, dt_in132, dt_in133, dt_in134, dt_in135, dt_in136, dt_in137, dt_in138, dt_in139, dt_in140, dt_in141, dt_in142, dt_in143, 
									dt_in144, dt_in145, dt_in146, dt_in147, dt_in148, dt_in149, dt_in150, dt_in151, dt_in152, dt_in153, dt_in154, dt_in155, dt_in156, dt_in157, dt_in158, dt_in159, 
									dt_in160, dt_in161, dt_in162, dt_in163, dt_in164, dt_in165, dt_in166, dt_in167, dt_in168, dt_in169, dt_in170, dt_in171, dt_in172, dt_in173, dt_in174, dt_in175, 
									dt_in176, dt_in177, dt_in178, dt_in179, dt_in180, dt_in181, dt_in182, dt_in183, dt_in184, dt_in185, dt_in186, dt_in187, dt_in188, dt_in189, dt_in190, dt_in191, 
									dt_in192, dt_in193, dt_in194, dt_in195, dt_in196, dt_in197, dt_in198, dt_in199, dt_in200, dt_in201, dt_in202, dt_in203, dt_in204, dt_in205, dt_in206, dt_in207, 
									dt_in208, dt_in209, dt_in210, dt_in211, dt_in212, dt_in213, dt_in214, dt_in215, dt_in216, dt_in217, dt_in218, dt_in219, dt_in220, dt_in221, dt_in222, dt_in223, 
									dt_in224, dt_in225, dt_in226, dt_in227, dt_in228, dt_in229, dt_in230, dt_in231, dt_in232, dt_in233, dt_in234, dt_in235, dt_in236, dt_in237, dt_in238, dt_in239, 
									dt_in240, dt_in241, dt_in242, dt_in243, dt_in244, dt_in245, dt_in246, dt_in247, dt_in248, dt_in249, dt_in250, dt_in251, dt_in252, dt_in253, dt_in254, dt_in255, 
									dt_in256, dt_in257, dt_in258, dt_in259, dt_in260, dt_in261, dt_in262, dt_in263, dt_in264, dt_in265, dt_in266, dt_in267, dt_in268, dt_in269, dt_in270, dt_in271, 
									dt_in272, dt_in273, dt_in274, dt_in275, dt_in276, dt_in277, dt_in278, dt_in279, dt_in280, dt_in281, dt_in282, dt_in283, dt_in284, dt_in285, dt_in286, dt_in287, 
									dt_in288, dt_in289, dt_in290, dt_in291, dt_in292, dt_in293, dt_in294, dt_in295, dt_in296, dt_in297, dt_in298, dt_in299, dt_in300, dt_in301, dt_in302, dt_in303, 
									dt_in304, dt_in305, dt_in306, dt_in307, dt_in308, dt_in309, dt_in310, dt_in311, dt_in312, dt_in313, dt_in314, dt_in315, dt_in316, dt_in317, dt_in318, dt_in319, 
									dt_in320, dt_in321, dt_in322, dt_in323, dt_in324, dt_in325, dt_in326, dt_in327, dt_in328, dt_in329, dt_in330, dt_in331, dt_in332, dt_in333, dt_in334, dt_in335, 
									dt_in336, dt_in337, dt_in338, dt_in339, dt_in340, dt_in341, dt_in342, dt_in343, dt_in344, dt_in345, dt_in346, dt_in347, dt_in348, dt_in349, dt_in350, dt_in351, 
									dt_in352, dt_in353, dt_in354, dt_in355, dt_in356, dt_in357, dt_in358, dt_in359, dt_in360, dt_in361, dt_in362, dt_in363, dt_in364, dt_in365, dt_in366, dt_in367, 
									dt_in368, dt_in369, dt_in370, dt_in371, dt_in372, dt_in373, dt_in374, dt_in375, dt_in376, dt_in377, dt_in378, dt_in379, dt_in380, dt_in381, dt_in382, dt_in383, 
									dt_in384, dt_in385, dt_in386, dt_in387, dt_in388, dt_in389, dt_in390, dt_in391, dt_in392, dt_in393, dt_in394, dt_in395, dt_in396, dt_in397, dt_in398, dt_in399, 
									dt_in400, dt_in401, dt_in402, dt_in403, dt_in404, dt_in405, dt_in406, dt_in407, dt_in408, dt_in409, dt_in410, dt_in411, dt_in412, dt_in413, dt_in414, dt_in415, 
									dt_in416, dt_in417, dt_in418, dt_in419, dt_in420, dt_in421, dt_in422, dt_in423, dt_in424, dt_in425, dt_in426, dt_in427, dt_in428, dt_in429, dt_in430, dt_in431, 
									dt_in432, dt_in433, dt_in434, dt_in435, dt_in436, dt_in437, dt_in438, dt_in439, dt_in440, dt_in441, dt_in442, dt_in443, dt_in444, dt_in445, dt_in446, dt_in447, 
									dt_in448, dt_in449, dt_in450, dt_in451, dt_in452, dt_in453, dt_in454, dt_in455, dt_in456, dt_in457, dt_in458, dt_in459, dt_in460, dt_in461, dt_in462, dt_in463, 
									dt_in464, dt_in465, dt_in466, dt_in467, dt_in468, dt_in469, dt_in470, dt_in471, dt_in472, dt_in473, dt_in474, dt_in475, dt_in476, dt_in477, dt_in478, dt_in479, 
									dt_in480, dt_in481, dt_in482, dt_in483, dt_in484, dt_in485, dt_in486, dt_in487, dt_in488, dt_in489, dt_in490, dt_in491, dt_in492, dt_in493, dt_in494, dt_in495, 
									dt_in496, dt_in497, dt_in498, dt_in499, dt_in500, dt_in501, dt_in502, dt_in503, dt_in504, dt_in505, dt_in506, dt_in507, dt_in508, dt_in509, dt_in510, dt_in511, 
									dt_in512, dt_in513, dt_in514, dt_in515, dt_in516, dt_in517, dt_in518, dt_in519, dt_in520, dt_in521, dt_in522, dt_in523, dt_in524, dt_in525, dt_in526, dt_in527, 
									dt_in528, dt_in529, dt_in530, dt_in531, dt_in532, dt_in533, dt_in534, dt_in535, dt_in536, dt_in537, dt_in538, dt_in539, dt_in540, dt_in541, dt_in542, dt_in543, 
									dt_in544, dt_in545, dt_in546, dt_in547, dt_in548, dt_in549, dt_in550, dt_in551, dt_in552, dt_in553, dt_in554, dt_in555, dt_in556, dt_in557, dt_in558, dt_in559, 
									dt_in560, dt_in561, dt_in562, dt_in563, dt_in564, dt_in565, dt_in566, dt_in567, dt_in568, dt_in569, dt_in570, dt_in571, dt_in572, dt_in573, dt_in574, dt_in575, 
									dt_in576, dt_in577, dt_in578, dt_in579, dt_in580, dt_in581, dt_in582, dt_in583, dt_in584, dt_in585, dt_in586, dt_in587, dt_in588, dt_in589, dt_in590, dt_in591, 
									dt_in592, dt_in593, dt_in594, dt_in595, dt_in596, dt_in597, dt_in598, dt_in599, dt_in600, dt_in601, dt_in602, dt_in603, dt_in604, dt_in605, dt_in606, dt_in607, 
									dt_in608, dt_in609, dt_in610, dt_in611, dt_in612, dt_in613, dt_in614, dt_in615, dt_in616, dt_in617, dt_in618, dt_in619, dt_in620, dt_in621, dt_in622, dt_in623, 
									dt_in624, dt_in625, dt_in626, dt_in627, dt_in628, dt_in629, dt_in630, dt_in631, dt_in632, dt_in633, dt_in634, dt_in635, dt_in636, dt_in637, dt_in638, dt_in639, 
									dt_in640, dt_in641, dt_in642, dt_in643, dt_in644, dt_in645, dt_in646, dt_in647, dt_in648, dt_in649, dt_in650, dt_in651, dt_in652, dt_in653, dt_in654, dt_in655, 
									dt_in656, dt_in657, dt_in658, dt_in659, dt_in660, dt_in661, dt_in662, dt_in663, dt_in664, dt_in665, dt_in666, dt_in667, dt_in668, dt_in669, dt_in670, dt_in671, 
									dt_in672, dt_in673, dt_in674, dt_in675, dt_in676, dt_in677, dt_in678, dt_in679, dt_in680, dt_in681, dt_in682, dt_in683, dt_in684, dt_in685, dt_in686, dt_in687, 
									dt_in688, dt_in689, dt_in690, dt_in691, dt_in692, dt_in693, dt_in694, dt_in695, dt_in696, dt_in697, dt_in698, dt_in699, dt_in700, dt_in701, dt_in702, dt_in703, 
									dt_in704, dt_in705, dt_in706, dt_in707, dt_in708, dt_in709, dt_in710, dt_in711, dt_in712, dt_in713, dt_in714, dt_in715, dt_in716, dt_in717, dt_in718, dt_in719, 
									dt_in720, dt_in721, dt_in722, dt_in723, dt_in724, dt_in725, dt_in726, dt_in727, dt_in728, dt_in729, dt_in730, dt_in731, dt_in732, dt_in733, dt_in734, dt_in735, 
									dt_in736, dt_in737, dt_in738, dt_in739, dt_in740, dt_in741, dt_in742, dt_in743, dt_in744, dt_in745, dt_in746, dt_in747, dt_in748, dt_in749, dt_in750, dt_in751, 
									dt_in752, dt_in753, dt_in754, dt_in755, dt_in756, dt_in757, dt_in758, dt_in759, dt_in760, dt_in761, dt_in762, dt_in763, dt_in764, dt_in765, dt_in766, dt_in767, 
									dt_in768, dt_in769, dt_in770, dt_in771, dt_in772, dt_in773, dt_in774, dt_in775, dt_in776, dt_in777, dt_in778, dt_in779, dt_in780, dt_in781, dt_in782, dt_in783, 
									dt_in784, dt_in785, dt_in786, dt_in787, dt_in788, dt_in789, dt_in790, dt_in791, dt_in792, dt_in793, dt_in794, dt_in795, dt_in796, dt_in797, dt_in798, dt_in799, 
									dt_in800, dt_in801, dt_in802, dt_in803, dt_in804, dt_in805, dt_in806, dt_in807, dt_in808, dt_in809, dt_in810, dt_in811, dt_in812, dt_in813, dt_in814, dt_in815, 
									dt_in816, dt_in817, dt_in818, dt_in819, dt_in820, dt_in821, dt_in822, dt_in823, dt_in824, dt_in825, dt_in826, dt_in827, dt_in828, dt_in829, dt_in830, dt_in831, 
									dt_in832, dt_in833, dt_in834, dt_in835, dt_in836, dt_in837, dt_in838, dt_in839, dt_in840, dt_in841, dt_in842, dt_in843, dt_in844, dt_in845, dt_in846, dt_in847, 
									dt_in848, dt_in849, dt_in850, dt_in851, dt_in852, dt_in853, dt_in854, dt_in855, dt_in856, dt_in857, dt_in858, dt_in859, dt_in860, dt_in861, dt_in862, dt_in863, 
									dt_in864, dt_in865, dt_in866, dt_in867, dt_in868, dt_in869, dt_in870, dt_in871, dt_in872, dt_in873, dt_in874, dt_in875, dt_in876, dt_in877, dt_in878, dt_in879, 
									dt_in880, dt_in881, dt_in882, dt_in883, dt_in884, dt_in885, dt_in886, dt_in887, dt_in888, dt_in889, dt_in890, dt_in891, dt_in892, dt_in893, dt_in894, dt_in895, 
									dt_in896, dt_in897, dt_in898, dt_in899, dt_in900, dt_in901, dt_in902, dt_in903, dt_in904, dt_in905, dt_in906, dt_in907, dt_in908, dt_in909, dt_in910, dt_in911, 
									dt_in912, dt_in913, dt_in914, dt_in915, dt_in916, dt_in917, dt_in918, dt_in919, dt_in920, dt_in921, dt_in922, dt_in923, dt_in924, dt_in925, dt_in926, dt_in927, 
									dt_in928, dt_in929, dt_in930, dt_in931, dt_in932, dt_in933, dt_in934, dt_in935, dt_in936, dt_in937, dt_in938, dt_in939, dt_in940, dt_in941, dt_in942, dt_in943, 
									dt_in944, dt_in945, dt_in946, dt_in947, dt_in948, dt_in949, dt_in950, dt_in951, dt_in952, dt_in953, dt_in954, dt_in955, dt_in956, dt_in957, dt_in958, dt_in959, 
									dt_in960, dt_in961, dt_in962, dt_in963, dt_in964, dt_in965, dt_in966, dt_in967, dt_in968, dt_in969, dt_in970, dt_in971, dt_in972, dt_in973, dt_in974, dt_in975, 
									dt_in976, dt_in977, dt_in978, dt_in979, dt_in980, dt_in981, dt_in982, dt_in983, dt_in984, dt_in985, dt_in986, dt_in987, dt_in988, dt_in989, dt_in990, dt_in991, 
									dt_in992, dt_in993, dt_in994, dt_in995, dt_in996, dt_in997, dt_in998, dt_in999, dt_in1000, dt_in1001, dt_in1002, dt_in1003, dt_in1004, dt_in1005, dt_in1006, dt_in1007, 
									dt_in1008, dt_in1009, dt_in1010, dt_in1011, dt_in1012, dt_in1013, dt_in1014, dt_in1015, dt_in1016, dt_in1017, dt_in1018, dt_in1019, dt_in1020, dt_in1021, dt_in1022, dt_in1023;


	wire signed [hwidth-1:0] 		dt_out0, dt_out1, dt_out2, dt_out3, dt_out4, dt_out5, dt_out6, dt_out7, dt_out8, dt_out9, dt_out10, dt_out11, dt_out12, dt_out13, dt_out14, dt_out15, 
									dt_out16, dt_out17, dt_out18, dt_out19, dt_out20, dt_out21, dt_out22, dt_out23, dt_out24, dt_out25, dt_out26, dt_out27, dt_out28, dt_out29, dt_out30, dt_out31, 
									dt_out32, dt_out33, dt_out34, dt_out35, dt_out36, dt_out37, dt_out38, dt_out39, dt_out40, dt_out41, dt_out42, dt_out43, dt_out44, dt_out45, dt_out46, dt_out47, 
									dt_out48, dt_out49, dt_out50, dt_out51, dt_out52, dt_out53, dt_out54, dt_out55, dt_out56, dt_out57, dt_out58, dt_out59, dt_out60, dt_out61, dt_out62, dt_out63, 
									dt_out64, dt_out65, dt_out66, dt_out67, dt_out68, dt_out69, dt_out70, dt_out71, dt_out72, dt_out73, dt_out74, dt_out75, dt_out76, dt_out77, dt_out78, dt_out79, 
									dt_out80, dt_out81, dt_out82, dt_out83, dt_out84, dt_out85, dt_out86, dt_out87, dt_out88, dt_out89, dt_out90, dt_out91, dt_out92, dt_out93, dt_out94, dt_out95, 
									dt_out96, dt_out97, dt_out98, dt_out99, dt_out100, dt_out101, dt_out102, dt_out103, dt_out104, dt_out105, dt_out106, dt_out107, dt_out108, dt_out109, dt_out110, dt_out111, 
									dt_out112, dt_out113, dt_out114, dt_out115, dt_out116, dt_out117, dt_out118, dt_out119, dt_out120, dt_out121, dt_out122, dt_out123, dt_out124, dt_out125, dt_out126, dt_out127, 
									dt_out128, dt_out129, dt_out130, dt_out131, dt_out132, dt_out133, dt_out134, dt_out135, dt_out136, dt_out137, dt_out138, dt_out139, dt_out140, dt_out141, dt_out142, dt_out143, 
									dt_out144, dt_out145, dt_out146, dt_out147, dt_out148, dt_out149, dt_out150, dt_out151, dt_out152, dt_out153, dt_out154, dt_out155, dt_out156, dt_out157, dt_out158, dt_out159, 
									dt_out160, dt_out161, dt_out162, dt_out163, dt_out164, dt_out165, dt_out166, dt_out167, dt_out168, dt_out169, dt_out170, dt_out171, dt_out172, dt_out173, dt_out174, dt_out175, 
									dt_out176, dt_out177, dt_out178, dt_out179, dt_out180, dt_out181, dt_out182, dt_out183, dt_out184, dt_out185, dt_out186, dt_out187, dt_out188, dt_out189, dt_out190, dt_out191, 
									dt_out192, dt_out193, dt_out194, dt_out195, dt_out196, dt_out197, dt_out198, dt_out199, dt_out200, dt_out201, dt_out202, dt_out203, dt_out204, dt_out205, dt_out206, dt_out207, 
									dt_out208, dt_out209, dt_out210, dt_out211, dt_out212, dt_out213, dt_out214, dt_out215, dt_out216, dt_out217, dt_out218, dt_out219, dt_out220, dt_out221, dt_out222, dt_out223, 
									dt_out224, dt_out225, dt_out226, dt_out227, dt_out228, dt_out229, dt_out230, dt_out231, dt_out232, dt_out233, dt_out234, dt_out235, dt_out236, dt_out237, dt_out238, dt_out239, 
									dt_out240, dt_out241, dt_out242, dt_out243, dt_out244, dt_out245, dt_out246, dt_out247, dt_out248, dt_out249, dt_out250, dt_out251, dt_out252, dt_out253, dt_out254, dt_out255, 
									dt_out256, dt_out257, dt_out258, dt_out259, dt_out260, dt_out261, dt_out262, dt_out263, dt_out264, dt_out265, dt_out266, dt_out267, dt_out268, dt_out269, dt_out270, dt_out271, 
									dt_out272, dt_out273, dt_out274, dt_out275, dt_out276, dt_out277, dt_out278, dt_out279, dt_out280, dt_out281, dt_out282, dt_out283, dt_out284, dt_out285, dt_out286, dt_out287, 
									dt_out288, dt_out289, dt_out290, dt_out291, dt_out292, dt_out293, dt_out294, dt_out295, dt_out296, dt_out297, dt_out298, dt_out299, dt_out300, dt_out301, dt_out302, dt_out303, 
									dt_out304, dt_out305, dt_out306, dt_out307, dt_out308, dt_out309, dt_out310, dt_out311, dt_out312, dt_out313, dt_out314, dt_out315, dt_out316, dt_out317, dt_out318, dt_out319, 
									dt_out320, dt_out321, dt_out322, dt_out323, dt_out324, dt_out325, dt_out326, dt_out327, dt_out328, dt_out329, dt_out330, dt_out331, dt_out332, dt_out333, dt_out334, dt_out335, 
									dt_out336, dt_out337, dt_out338, dt_out339, dt_out340, dt_out341, dt_out342, dt_out343, dt_out344, dt_out345, dt_out346, dt_out347, dt_out348, dt_out349, dt_out350, dt_out351, 
									dt_out352, dt_out353, dt_out354, dt_out355, dt_out356, dt_out357, dt_out358, dt_out359, dt_out360, dt_out361, dt_out362, dt_out363, dt_out364, dt_out365, dt_out366, dt_out367, 
									dt_out368, dt_out369, dt_out370, dt_out371, dt_out372, dt_out373, dt_out374, dt_out375, dt_out376, dt_out377, dt_out378, dt_out379, dt_out380, dt_out381, dt_out382, dt_out383, 
									dt_out384, dt_out385, dt_out386, dt_out387, dt_out388, dt_out389, dt_out390, dt_out391, dt_out392, dt_out393, dt_out394, dt_out395, dt_out396, dt_out397, dt_out398, dt_out399, 
									dt_out400, dt_out401, dt_out402, dt_out403, dt_out404, dt_out405, dt_out406, dt_out407, dt_out408, dt_out409, dt_out410, dt_out411, dt_out412, dt_out413, dt_out414, dt_out415, 
									dt_out416, dt_out417, dt_out418, dt_out419, dt_out420, dt_out421, dt_out422, dt_out423, dt_out424, dt_out425, dt_out426, dt_out427, dt_out428, dt_out429, dt_out430, dt_out431, 
									dt_out432, dt_out433, dt_out434, dt_out435, dt_out436, dt_out437, dt_out438, dt_out439, dt_out440, dt_out441, dt_out442, dt_out443, dt_out444, dt_out445, dt_out446, dt_out447, 
									dt_out448, dt_out449, dt_out450, dt_out451, dt_out452, dt_out453, dt_out454, dt_out455, dt_out456, dt_out457, dt_out458, dt_out459, dt_out460, dt_out461, dt_out462, dt_out463, 
									dt_out464, dt_out465, dt_out466, dt_out467, dt_out468, dt_out469, dt_out470, dt_out471, dt_out472, dt_out473, dt_out474, dt_out475, dt_out476, dt_out477, dt_out478, dt_out479, 
									dt_out480, dt_out481, dt_out482, dt_out483, dt_out484, dt_out485, dt_out486, dt_out487, dt_out488, dt_out489, dt_out490, dt_out491, dt_out492, dt_out493, dt_out494, dt_out495, 
									dt_out496, dt_out497, dt_out498, dt_out499, dt_out500, dt_out501, dt_out502, dt_out503, dt_out504, dt_out505, dt_out506, dt_out507, dt_out508, dt_out509, dt_out510, dt_out511, 
									dt_out512, dt_out513, dt_out514, dt_out515, dt_out516, dt_out517, dt_out518, dt_out519, dt_out520, dt_out521, dt_out522, dt_out523, dt_out524, dt_out525, dt_out526, dt_out527, 
									dt_out528, dt_out529, dt_out530, dt_out531, dt_out532, dt_out533, dt_out534, dt_out535, dt_out536, dt_out537, dt_out538, dt_out539, dt_out540, dt_out541, dt_out542, dt_out543, 
									dt_out544, dt_out545, dt_out546, dt_out547, dt_out548, dt_out549, dt_out550, dt_out551, dt_out552, dt_out553, dt_out554, dt_out555, dt_out556, dt_out557, dt_out558, dt_out559, 
									dt_out560, dt_out561, dt_out562, dt_out563, dt_out564, dt_out565, dt_out566, dt_out567, dt_out568, dt_out569, dt_out570, dt_out571, dt_out572, dt_out573, dt_out574, dt_out575, 
									dt_out576, dt_out577, dt_out578, dt_out579, dt_out580, dt_out581, dt_out582, dt_out583, dt_out584, dt_out585, dt_out586, dt_out587, dt_out588, dt_out589, dt_out590, dt_out591, 
									dt_out592, dt_out593, dt_out594, dt_out595, dt_out596, dt_out597, dt_out598, dt_out599, dt_out600, dt_out601, dt_out602, dt_out603, dt_out604, dt_out605, dt_out606, dt_out607, 
									dt_out608, dt_out609, dt_out610, dt_out611, dt_out612, dt_out613, dt_out614, dt_out615, dt_out616, dt_out617, dt_out618, dt_out619, dt_out620, dt_out621, dt_out622, dt_out623, 
									dt_out624, dt_out625, dt_out626, dt_out627, dt_out628, dt_out629, dt_out630, dt_out631, dt_out632, dt_out633, dt_out634, dt_out635, dt_out636, dt_out637, dt_out638, dt_out639, 
									dt_out640, dt_out641, dt_out642, dt_out643, dt_out644, dt_out645, dt_out646, dt_out647, dt_out648, dt_out649, dt_out650, dt_out651, dt_out652, dt_out653, dt_out654, dt_out655, 
									dt_out656, dt_out657, dt_out658, dt_out659, dt_out660, dt_out661, dt_out662, dt_out663, dt_out664, dt_out665, dt_out666, dt_out667, dt_out668, dt_out669, dt_out670, dt_out671, 
									dt_out672, dt_out673, dt_out674, dt_out675, dt_out676, dt_out677, dt_out678, dt_out679, dt_out680, dt_out681, dt_out682, dt_out683, dt_out684, dt_out685, dt_out686, dt_out687, 
									dt_out688, dt_out689, dt_out690, dt_out691, dt_out692, dt_out693, dt_out694, dt_out695, dt_out696, dt_out697, dt_out698, dt_out699, dt_out700, dt_out701, dt_out702, dt_out703, 
									dt_out704, dt_out705, dt_out706, dt_out707, dt_out708, dt_out709, dt_out710, dt_out711, dt_out712, dt_out713, dt_out714, dt_out715, dt_out716, dt_out717, dt_out718, dt_out719, 
									dt_out720, dt_out721, dt_out722, dt_out723, dt_out724, dt_out725, dt_out726, dt_out727, dt_out728, dt_out729, dt_out730, dt_out731, dt_out732, dt_out733, dt_out734, dt_out735, 
									dt_out736, dt_out737, dt_out738, dt_out739, dt_out740, dt_out741, dt_out742, dt_out743, dt_out744, dt_out745, dt_out746, dt_out747, dt_out748, dt_out749, dt_out750, dt_out751, 
									dt_out752, dt_out753, dt_out754, dt_out755, dt_out756, dt_out757, dt_out758, dt_out759, dt_out760, dt_out761, dt_out762, dt_out763, dt_out764, dt_out765, dt_out766, dt_out767, 
									dt_out768, dt_out769, dt_out770, dt_out771, dt_out772, dt_out773, dt_out774, dt_out775, dt_out776, dt_out777, dt_out778, dt_out779, dt_out780, dt_out781, dt_out782, dt_out783, 
									dt_out784, dt_out785, dt_out786, dt_out787, dt_out788, dt_out789, dt_out790, dt_out791, dt_out792, dt_out793, dt_out794, dt_out795, dt_out796, dt_out797, dt_out798, dt_out799, 
									dt_out800, dt_out801, dt_out802, dt_out803, dt_out804, dt_out805, dt_out806, dt_out807, dt_out808, dt_out809, dt_out810, dt_out811, dt_out812, dt_out813, dt_out814, dt_out815, 
									dt_out816, dt_out817, dt_out818, dt_out819, dt_out820, dt_out821, dt_out822, dt_out823, dt_out824, dt_out825, dt_out826, dt_out827, dt_out828, dt_out829, dt_out830, dt_out831, 
									dt_out832, dt_out833, dt_out834, dt_out835, dt_out836, dt_out837, dt_out838, dt_out839, dt_out840, dt_out841, dt_out842, dt_out843, dt_out844, dt_out845, dt_out846, dt_out847, 
									dt_out848, dt_out849, dt_out850, dt_out851, dt_out852, dt_out853, dt_out854, dt_out855, dt_out856, dt_out857, dt_out858, dt_out859, dt_out860, dt_out861, dt_out862, dt_out863, 
									dt_out864, dt_out865, dt_out866, dt_out867, dt_out868, dt_out869, dt_out870, dt_out871, dt_out872, dt_out873, dt_out874, dt_out875, dt_out876, dt_out877, dt_out878, dt_out879, 
									dt_out880, dt_out881, dt_out882, dt_out883, dt_out884, dt_out885, dt_out886, dt_out887, dt_out888, dt_out889, dt_out890, dt_out891, dt_out892, dt_out893, dt_out894, dt_out895, 
									dt_out896, dt_out897, dt_out898, dt_out899, dt_out900, dt_out901, dt_out902, dt_out903, dt_out904, dt_out905, dt_out906, dt_out907, dt_out908, dt_out909, dt_out910, dt_out911, 
									dt_out912, dt_out913, dt_out914, dt_out915, dt_out916, dt_out917, dt_out918, dt_out919, dt_out920, dt_out921, dt_out922, dt_out923, dt_out924, dt_out925, dt_out926, dt_out927, 
									dt_out928, dt_out929, dt_out930, dt_out931, dt_out932, dt_out933, dt_out934, dt_out935, dt_out936, dt_out937, dt_out938, dt_out939, dt_out940, dt_out941, dt_out942, dt_out943, 
									dt_out944, dt_out945, dt_out946, dt_out947, dt_out948, dt_out949, dt_out950, dt_out951, dt_out952, dt_out953, dt_out954, dt_out955, dt_out956, dt_out957, dt_out958, dt_out959, 
									dt_out960, dt_out961, dt_out962, dt_out963, dt_out964, dt_out965, dt_out966, dt_out967, dt_out968, dt_out969, dt_out970, dt_out971, dt_out972, dt_out973, dt_out974, dt_out975, 
									dt_out976, dt_out977, dt_out978, dt_out979, dt_out980, dt_out981, dt_out982, dt_out983, dt_out984, dt_out985, dt_out986, dt_out987, dt_out988, dt_out989, dt_out990, dt_out991, 
									dt_out992, dt_out993, dt_out994, dt_out995, dt_out996, dt_out997, dt_out998, dt_out999, dt_out1000, dt_out1001, dt_out1002, dt_out1003, dt_out1004, dt_out1005, dt_out1006, dt_out1007, 
									dt_out1008, dt_out1009, dt_out1010, dt_out1011, dt_out1012, dt_out1013, dt_out1014, dt_out1015, dt_out1016, dt_out1017, dt_out1018, dt_out1019, dt_out1020, dt_out1021, dt_out1022, dt_out1023;

// read input from file
		vcReadFile #(.size(1), .filename(`TV_INFILE), .hwidth(hwidth))
			inst_vcReadFile (clk, n_rst, 
							n_stall, 
			 				dt_in0, dt_in1, dt_in2, dt_in3, dt_in4, dt_in5, dt_in6, dt_in7, dt_in8, dt_in9, dt_in10, dt_in11, dt_in12, dt_in13, dt_in14, dt_in15, 
							dt_in16, dt_in17, dt_in18, dt_in19, dt_in20, dt_in21, dt_in22, dt_in23, dt_in24, dt_in25, dt_in26, dt_in27, dt_in28, dt_in29, dt_in30, dt_in31, 
							dt_in32, dt_in33, dt_in34, dt_in35, dt_in36, dt_in37, dt_in38, dt_in39, dt_in40, dt_in41, dt_in42, dt_in43, dt_in44, dt_in45, dt_in46, dt_in47, 
							dt_in48, dt_in49, dt_in50, dt_in51, dt_in52, dt_in53, dt_in54, dt_in55, dt_in56, dt_in57, dt_in58, dt_in59, dt_in60, dt_in61, dt_in62, dt_in63, 
							dt_in64, dt_in65, dt_in66, dt_in67, dt_in68, dt_in69, dt_in70, dt_in71, dt_in72, dt_in73, dt_in74, dt_in75, dt_in76, dt_in77, dt_in78, dt_in79, 
							dt_in80, dt_in81, dt_in82, dt_in83, dt_in84, dt_in85, dt_in86, dt_in87, dt_in88, dt_in89, dt_in90, dt_in91, dt_in92, dt_in93, dt_in94, dt_in95, 
							dt_in96, dt_in97, dt_in98, dt_in99, dt_in100, dt_in101, dt_in102, dt_in103, dt_in104, dt_in105, dt_in106, dt_in107, dt_in108, dt_in109, dt_in110, dt_in111, 
							dt_in112, dt_in113, dt_in114, dt_in115, dt_in116, dt_in117, dt_in118, dt_in119, dt_in120, dt_in121, dt_in122, dt_in123, dt_in124, dt_in125, dt_in126, dt_in127, 
							dt_in128, dt_in129, dt_in130, dt_in131, dt_in132, dt_in133, dt_in134, dt_in135, dt_in136, dt_in137, dt_in138, dt_in139, dt_in140, dt_in141, dt_in142, dt_in143, 
							dt_in144, dt_in145, dt_in146, dt_in147, dt_in148, dt_in149, dt_in150, dt_in151, dt_in152, dt_in153, dt_in154, dt_in155, dt_in156, dt_in157, dt_in158, dt_in159, 
							dt_in160, dt_in161, dt_in162, dt_in163, dt_in164, dt_in165, dt_in166, dt_in167, dt_in168, dt_in169, dt_in170, dt_in171, dt_in172, dt_in173, dt_in174, dt_in175, 
							dt_in176, dt_in177, dt_in178, dt_in179, dt_in180, dt_in181, dt_in182, dt_in183, dt_in184, dt_in185, dt_in186, dt_in187, dt_in188, dt_in189, dt_in190, dt_in191, 
							dt_in192, dt_in193, dt_in194, dt_in195, dt_in196, dt_in197, dt_in198, dt_in199, dt_in200, dt_in201, dt_in202, dt_in203, dt_in204, dt_in205, dt_in206, dt_in207, 
							dt_in208, dt_in209, dt_in210, dt_in211, dt_in212, dt_in213, dt_in214, dt_in215, dt_in216, dt_in217, dt_in218, dt_in219, dt_in220, dt_in221, dt_in222, dt_in223, 
							dt_in224, dt_in225, dt_in226, dt_in227, dt_in228, dt_in229, dt_in230, dt_in231, dt_in232, dt_in233, dt_in234, dt_in235, dt_in236, dt_in237, dt_in238, dt_in239, 
							dt_in240, dt_in241, dt_in242, dt_in243, dt_in244, dt_in245, dt_in246, dt_in247, dt_in248, dt_in249, dt_in250, dt_in251, dt_in252, dt_in253, dt_in254, dt_in255, 
							dt_in256, dt_in257, dt_in258, dt_in259, dt_in260, dt_in261, dt_in262, dt_in263, dt_in264, dt_in265, dt_in266, dt_in267, dt_in268, dt_in269, dt_in270, dt_in271, 
							dt_in272, dt_in273, dt_in274, dt_in275, dt_in276, dt_in277, dt_in278, dt_in279, dt_in280, dt_in281, dt_in282, dt_in283, dt_in284, dt_in285, dt_in286, dt_in287, 
							dt_in288, dt_in289, dt_in290, dt_in291, dt_in292, dt_in293, dt_in294, dt_in295, dt_in296, dt_in297, dt_in298, dt_in299, dt_in300, dt_in301, dt_in302, dt_in303, 
							dt_in304, dt_in305, dt_in306, dt_in307, dt_in308, dt_in309, dt_in310, dt_in311, dt_in312, dt_in313, dt_in314, dt_in315, dt_in316, dt_in317, dt_in318, dt_in319, 
							dt_in320, dt_in321, dt_in322, dt_in323, dt_in324, dt_in325, dt_in326, dt_in327, dt_in328, dt_in329, dt_in330, dt_in331, dt_in332, dt_in333, dt_in334, dt_in335, 
							dt_in336, dt_in337, dt_in338, dt_in339, dt_in340, dt_in341, dt_in342, dt_in343, dt_in344, dt_in345, dt_in346, dt_in347, dt_in348, dt_in349, dt_in350, dt_in351, 
							dt_in352, dt_in353, dt_in354, dt_in355, dt_in356, dt_in357, dt_in358, dt_in359, dt_in360, dt_in361, dt_in362, dt_in363, dt_in364, dt_in365, dt_in366, dt_in367, 
							dt_in368, dt_in369, dt_in370, dt_in371, dt_in372, dt_in373, dt_in374, dt_in375, dt_in376, dt_in377, dt_in378, dt_in379, dt_in380, dt_in381, dt_in382, dt_in383, 
							dt_in384, dt_in385, dt_in386, dt_in387, dt_in388, dt_in389, dt_in390, dt_in391, dt_in392, dt_in393, dt_in394, dt_in395, dt_in396, dt_in397, dt_in398, dt_in399, 
							dt_in400, dt_in401, dt_in402, dt_in403, dt_in404, dt_in405, dt_in406, dt_in407, dt_in408, dt_in409, dt_in410, dt_in411, dt_in412, dt_in413, dt_in414, dt_in415, 
							dt_in416, dt_in417, dt_in418, dt_in419, dt_in420, dt_in421, dt_in422, dt_in423, dt_in424, dt_in425, dt_in426, dt_in427, dt_in428, dt_in429, dt_in430, dt_in431, 
							dt_in432, dt_in433, dt_in434, dt_in435, dt_in436, dt_in437, dt_in438, dt_in439, dt_in440, dt_in441, dt_in442, dt_in443, dt_in444, dt_in445, dt_in446, dt_in447, 
							dt_in448, dt_in449, dt_in450, dt_in451, dt_in452, dt_in453, dt_in454, dt_in455, dt_in456, dt_in457, dt_in458, dt_in459, dt_in460, dt_in461, dt_in462, dt_in463, 
							dt_in464, dt_in465, dt_in466, dt_in467, dt_in468, dt_in469, dt_in470, dt_in471, dt_in472, dt_in473, dt_in474, dt_in475, dt_in476, dt_in477, dt_in478, dt_in479, 
							dt_in480, dt_in481, dt_in482, dt_in483, dt_in484, dt_in485, dt_in486, dt_in487, dt_in488, dt_in489, dt_in490, dt_in491, dt_in492, dt_in493, dt_in494, dt_in495, 
							dt_in496, dt_in497, dt_in498, dt_in499, dt_in500, dt_in501, dt_in502, dt_in503, dt_in504, dt_in505, dt_in506, dt_in507, dt_in508, dt_in509, dt_in510, dt_in511, 
							dt_in512, dt_in513, dt_in514, dt_in515, dt_in516, dt_in517, dt_in518, dt_in519, dt_in520, dt_in521, dt_in522, dt_in523, dt_in524, dt_in525, dt_in526, dt_in527, 
							dt_in528, dt_in529, dt_in530, dt_in531, dt_in532, dt_in533, dt_in534, dt_in535, dt_in536, dt_in537, dt_in538, dt_in539, dt_in540, dt_in541, dt_in542, dt_in543, 
							dt_in544, dt_in545, dt_in546, dt_in547, dt_in548, dt_in549, dt_in550, dt_in551, dt_in552, dt_in553, dt_in554, dt_in555, dt_in556, dt_in557, dt_in558, dt_in559, 
							dt_in560, dt_in561, dt_in562, dt_in563, dt_in564, dt_in565, dt_in566, dt_in567, dt_in568, dt_in569, dt_in570, dt_in571, dt_in572, dt_in573, dt_in574, dt_in575, 
							dt_in576, dt_in577, dt_in578, dt_in579, dt_in580, dt_in581, dt_in582, dt_in583, dt_in584, dt_in585, dt_in586, dt_in587, dt_in588, dt_in589, dt_in590, dt_in591, 
							dt_in592, dt_in593, dt_in594, dt_in595, dt_in596, dt_in597, dt_in598, dt_in599, dt_in600, dt_in601, dt_in602, dt_in603, dt_in604, dt_in605, dt_in606, dt_in607, 
							dt_in608, dt_in609, dt_in610, dt_in611, dt_in612, dt_in613, dt_in614, dt_in615, dt_in616, dt_in617, dt_in618, dt_in619, dt_in620, dt_in621, dt_in622, dt_in623, 
							dt_in624, dt_in625, dt_in626, dt_in627, dt_in628, dt_in629, dt_in630, dt_in631, dt_in632, dt_in633, dt_in634, dt_in635, dt_in636, dt_in637, dt_in638, dt_in639, 
							dt_in640, dt_in641, dt_in642, dt_in643, dt_in644, dt_in645, dt_in646, dt_in647, dt_in648, dt_in649, dt_in650, dt_in651, dt_in652, dt_in653, dt_in654, dt_in655, 
							dt_in656, dt_in657, dt_in658, dt_in659, dt_in660, dt_in661, dt_in662, dt_in663, dt_in664, dt_in665, dt_in666, dt_in667, dt_in668, dt_in669, dt_in670, dt_in671, 
							dt_in672, dt_in673, dt_in674, dt_in675, dt_in676, dt_in677, dt_in678, dt_in679, dt_in680, dt_in681, dt_in682, dt_in683, dt_in684, dt_in685, dt_in686, dt_in687, 
							dt_in688, dt_in689, dt_in690, dt_in691, dt_in692, dt_in693, dt_in694, dt_in695, dt_in696, dt_in697, dt_in698, dt_in699, dt_in700, dt_in701, dt_in702, dt_in703, 
							dt_in704, dt_in705, dt_in706, dt_in707, dt_in708, dt_in709, dt_in710, dt_in711, dt_in712, dt_in713, dt_in714, dt_in715, dt_in716, dt_in717, dt_in718, dt_in719, 
							dt_in720, dt_in721, dt_in722, dt_in723, dt_in724, dt_in725, dt_in726, dt_in727, dt_in728, dt_in729, dt_in730, dt_in731, dt_in732, dt_in733, dt_in734, dt_in735, 
							dt_in736, dt_in737, dt_in738, dt_in739, dt_in740, dt_in741, dt_in742, dt_in743, dt_in744, dt_in745, dt_in746, dt_in747, dt_in748, dt_in749, dt_in750, dt_in751, 
							dt_in752, dt_in753, dt_in754, dt_in755, dt_in756, dt_in757, dt_in758, dt_in759, dt_in760, dt_in761, dt_in762, dt_in763, dt_in764, dt_in765, dt_in766, dt_in767, 
							dt_in768, dt_in769, dt_in770, dt_in771, dt_in772, dt_in773, dt_in774, dt_in775, dt_in776, dt_in777, dt_in778, dt_in779, dt_in780, dt_in781, dt_in782, dt_in783, 
							dt_in784, dt_in785, dt_in786, dt_in787, dt_in788, dt_in789, dt_in790, dt_in791, dt_in792, dt_in793, dt_in794, dt_in795, dt_in796, dt_in797, dt_in798, dt_in799, 
							dt_in800, dt_in801, dt_in802, dt_in803, dt_in804, dt_in805, dt_in806, dt_in807, dt_in808, dt_in809, dt_in810, dt_in811, dt_in812, dt_in813, dt_in814, dt_in815, 
							dt_in816, dt_in817, dt_in818, dt_in819, dt_in820, dt_in821, dt_in822, dt_in823, dt_in824, dt_in825, dt_in826, dt_in827, dt_in828, dt_in829, dt_in830, dt_in831, 
							dt_in832, dt_in833, dt_in834, dt_in835, dt_in836, dt_in837, dt_in838, dt_in839, dt_in840, dt_in841, dt_in842, dt_in843, dt_in844, dt_in845, dt_in846, dt_in847, 
							dt_in848, dt_in849, dt_in850, dt_in851, dt_in852, dt_in853, dt_in854, dt_in855, dt_in856, dt_in857, dt_in858, dt_in859, dt_in860, dt_in861, dt_in862, dt_in863, 
							dt_in864, dt_in865, dt_in866, dt_in867, dt_in868, dt_in869, dt_in870, dt_in871, dt_in872, dt_in873, dt_in874, dt_in875, dt_in876, dt_in877, dt_in878, dt_in879, 
							dt_in880, dt_in881, dt_in882, dt_in883, dt_in884, dt_in885, dt_in886, dt_in887, dt_in888, dt_in889, dt_in890, dt_in891, dt_in892, dt_in893, dt_in894, dt_in895, 
							dt_in896, dt_in897, dt_in898, dt_in899, dt_in900, dt_in901, dt_in902, dt_in903, dt_in904, dt_in905, dt_in906, dt_in907, dt_in908, dt_in909, dt_in910, dt_in911, 
							dt_in912, dt_in913, dt_in914, dt_in915, dt_in916, dt_in917, dt_in918, dt_in919, dt_in920, dt_in921, dt_in922, dt_in923, dt_in924, dt_in925, dt_in926, dt_in927, 
							dt_in928, dt_in929, dt_in930, dt_in931, dt_in932, dt_in933, dt_in934, dt_in935, dt_in936, dt_in937, dt_in938, dt_in939, dt_in940, dt_in941, dt_in942, dt_in943, 
							dt_in944, dt_in945, dt_in946, dt_in947, dt_in948, dt_in949, dt_in950, dt_in951, dt_in952, dt_in953, dt_in954, dt_in955, dt_in956, dt_in957, dt_in958, dt_in959, 
							dt_in960, dt_in961, dt_in962, dt_in963, dt_in964, dt_in965, dt_in966, dt_in967, dt_in968, dt_in969, dt_in970, dt_in971, dt_in972, dt_in973, dt_in974, dt_in975, 
							dt_in976, dt_in977, dt_in978, dt_in979, dt_in980, dt_in981, dt_in982, dt_in983, dt_in984, dt_in985, dt_in986, dt_in987, dt_in988, dt_in989, dt_in990, dt_in991, 
							dt_in992, dt_in993, dt_in994, dt_in995, dt_in996, dt_in997, dt_in998, dt_in999, dt_in1000, dt_in1001, dt_in1002, dt_in1003, dt_in1004, dt_in1005, dt_in1006, dt_in1007, 
							dt_in1008, dt_in1009, dt_in1010, dt_in1011, dt_in1012, dt_in1013, dt_in1014, dt_in1015, dt_in1016, dt_in1017, dt_in1018, dt_in1019, dt_in1020, dt_in1021, dt_in1022, dt_in1023);

	// write output data to file
		vcWriteFile #(.size(1), .filename(`TV_OUTFILE), .hwidth(hwidth))
			inst_vcWriteFile (clk, n_rst, 
							n_stall_out, 
			 				dt_out0, dt_out1, dt_out2, dt_out3, dt_out4, dt_out5, dt_out6, dt_out7, dt_out8, dt_out9, dt_out10, dt_out11, dt_out12, dt_out13, dt_out14, dt_out15, 
							dt_out16, dt_out17, dt_out18, dt_out19, dt_out20, dt_out21, dt_out22, dt_out23, dt_out24, dt_out25, dt_out26, dt_out27, dt_out28, dt_out29, dt_out30, dt_out31, 
							dt_out32, dt_out33, dt_out34, dt_out35, dt_out36, dt_out37, dt_out38, dt_out39, dt_out40, dt_out41, dt_out42, dt_out43, dt_out44, dt_out45, dt_out46, dt_out47, 
							dt_out48, dt_out49, dt_out50, dt_out51, dt_out52, dt_out53, dt_out54, dt_out55, dt_out56, dt_out57, dt_out58, dt_out59, dt_out60, dt_out61, dt_out62, dt_out63, 
							dt_out64, dt_out65, dt_out66, dt_out67, dt_out68, dt_out69, dt_out70, dt_out71, dt_out72, dt_out73, dt_out74, dt_out75, dt_out76, dt_out77, dt_out78, dt_out79, 
							dt_out80, dt_out81, dt_out82, dt_out83, dt_out84, dt_out85, dt_out86, dt_out87, dt_out88, dt_out89, dt_out90, dt_out91, dt_out92, dt_out93, dt_out94, dt_out95, 
							dt_out96, dt_out97, dt_out98, dt_out99, dt_out100, dt_out101, dt_out102, dt_out103, dt_out104, dt_out105, dt_out106, dt_out107, dt_out108, dt_out109, dt_out110, dt_out111, 
							dt_out112, dt_out113, dt_out114, dt_out115, dt_out116, dt_out117, dt_out118, dt_out119, dt_out120, dt_out121, dt_out122, dt_out123, dt_out124, dt_out125, dt_out126, dt_out127, 
							dt_out128, dt_out129, dt_out130, dt_out131, dt_out132, dt_out133, dt_out134, dt_out135, dt_out136, dt_out137, dt_out138, dt_out139, dt_out140, dt_out141, dt_out142, dt_out143, 
							dt_out144, dt_out145, dt_out146, dt_out147, dt_out148, dt_out149, dt_out150, dt_out151, dt_out152, dt_out153, dt_out154, dt_out155, dt_out156, dt_out157, dt_out158, dt_out159, 
							dt_out160, dt_out161, dt_out162, dt_out163, dt_out164, dt_out165, dt_out166, dt_out167, dt_out168, dt_out169, dt_out170, dt_out171, dt_out172, dt_out173, dt_out174, dt_out175, 
							dt_out176, dt_out177, dt_out178, dt_out179, dt_out180, dt_out181, dt_out182, dt_out183, dt_out184, dt_out185, dt_out186, dt_out187, dt_out188, dt_out189, dt_out190, dt_out191, 
							dt_out192, dt_out193, dt_out194, dt_out195, dt_out196, dt_out197, dt_out198, dt_out199, dt_out200, dt_out201, dt_out202, dt_out203, dt_out204, dt_out205, dt_out206, dt_out207, 
							dt_out208, dt_out209, dt_out210, dt_out211, dt_out212, dt_out213, dt_out214, dt_out215, dt_out216, dt_out217, dt_out218, dt_out219, dt_out220, dt_out221, dt_out222, dt_out223, 
							dt_out224, dt_out225, dt_out226, dt_out227, dt_out228, dt_out229, dt_out230, dt_out231, dt_out232, dt_out233, dt_out234, dt_out235, dt_out236, dt_out237, dt_out238, dt_out239, 
							dt_out240, dt_out241, dt_out242, dt_out243, dt_out244, dt_out245, dt_out246, dt_out247, dt_out248, dt_out249, dt_out250, dt_out251, dt_out252, dt_out253, dt_out254, dt_out255, 
							dt_out256, dt_out257, dt_out258, dt_out259, dt_out260, dt_out261, dt_out262, dt_out263, dt_out264, dt_out265, dt_out266, dt_out267, dt_out268, dt_out269, dt_out270, dt_out271, 
							dt_out272, dt_out273, dt_out274, dt_out275, dt_out276, dt_out277, dt_out278, dt_out279, dt_out280, dt_out281, dt_out282, dt_out283, dt_out284, dt_out285, dt_out286, dt_out287, 
							dt_out288, dt_out289, dt_out290, dt_out291, dt_out292, dt_out293, dt_out294, dt_out295, dt_out296, dt_out297, dt_out298, dt_out299, dt_out300, dt_out301, dt_out302, dt_out303, 
							dt_out304, dt_out305, dt_out306, dt_out307, dt_out308, dt_out309, dt_out310, dt_out311, dt_out312, dt_out313, dt_out314, dt_out315, dt_out316, dt_out317, dt_out318, dt_out319, 
							dt_out320, dt_out321, dt_out322, dt_out323, dt_out324, dt_out325, dt_out326, dt_out327, dt_out328, dt_out329, dt_out330, dt_out331, dt_out332, dt_out333, dt_out334, dt_out335, 
							dt_out336, dt_out337, dt_out338, dt_out339, dt_out340, dt_out341, dt_out342, dt_out343, dt_out344, dt_out345, dt_out346, dt_out347, dt_out348, dt_out349, dt_out350, dt_out351, 
							dt_out352, dt_out353, dt_out354, dt_out355, dt_out356, dt_out357, dt_out358, dt_out359, dt_out360, dt_out361, dt_out362, dt_out363, dt_out364, dt_out365, dt_out366, dt_out367, 
							dt_out368, dt_out369, dt_out370, dt_out371, dt_out372, dt_out373, dt_out374, dt_out375, dt_out376, dt_out377, dt_out378, dt_out379, dt_out380, dt_out381, dt_out382, dt_out383, 
							dt_out384, dt_out385, dt_out386, dt_out387, dt_out388, dt_out389, dt_out390, dt_out391, dt_out392, dt_out393, dt_out394, dt_out395, dt_out396, dt_out397, dt_out398, dt_out399, 
							dt_out400, dt_out401, dt_out402, dt_out403, dt_out404, dt_out405, dt_out406, dt_out407, dt_out408, dt_out409, dt_out410, dt_out411, dt_out412, dt_out413, dt_out414, dt_out415, 
							dt_out416, dt_out417, dt_out418, dt_out419, dt_out420, dt_out421, dt_out422, dt_out423, dt_out424, dt_out425, dt_out426, dt_out427, dt_out428, dt_out429, dt_out430, dt_out431, 
							dt_out432, dt_out433, dt_out434, dt_out435, dt_out436, dt_out437, dt_out438, dt_out439, dt_out440, dt_out441, dt_out442, dt_out443, dt_out444, dt_out445, dt_out446, dt_out447, 
							dt_out448, dt_out449, dt_out450, dt_out451, dt_out452, dt_out453, dt_out454, dt_out455, dt_out456, dt_out457, dt_out458, dt_out459, dt_out460, dt_out461, dt_out462, dt_out463, 
							dt_out464, dt_out465, dt_out466, dt_out467, dt_out468, dt_out469, dt_out470, dt_out471, dt_out472, dt_out473, dt_out474, dt_out475, dt_out476, dt_out477, dt_out478, dt_out479, 
							dt_out480, dt_out481, dt_out482, dt_out483, dt_out484, dt_out485, dt_out486, dt_out487, dt_out488, dt_out489, dt_out490, dt_out491, dt_out492, dt_out493, dt_out494, dt_out495, 
							dt_out496, dt_out497, dt_out498, dt_out499, dt_out500, dt_out501, dt_out502, dt_out503, dt_out504, dt_out505, dt_out506, dt_out507, dt_out508, dt_out509, dt_out510, dt_out511, 
							dt_out512, dt_out513, dt_out514, dt_out515, dt_out516, dt_out517, dt_out518, dt_out519, dt_out520, dt_out521, dt_out522, dt_out523, dt_out524, dt_out525, dt_out526, dt_out527, 
							dt_out528, dt_out529, dt_out530, dt_out531, dt_out532, dt_out533, dt_out534, dt_out535, dt_out536, dt_out537, dt_out538, dt_out539, dt_out540, dt_out541, dt_out542, dt_out543, 
							dt_out544, dt_out545, dt_out546, dt_out547, dt_out548, dt_out549, dt_out550, dt_out551, dt_out552, dt_out553, dt_out554, dt_out555, dt_out556, dt_out557, dt_out558, dt_out559, 
							dt_out560, dt_out561, dt_out562, dt_out563, dt_out564, dt_out565, dt_out566, dt_out567, dt_out568, dt_out569, dt_out570, dt_out571, dt_out572, dt_out573, dt_out574, dt_out575, 
							dt_out576, dt_out577, dt_out578, dt_out579, dt_out580, dt_out581, dt_out582, dt_out583, dt_out584, dt_out585, dt_out586, dt_out587, dt_out588, dt_out589, dt_out590, dt_out591, 
							dt_out592, dt_out593, dt_out594, dt_out595, dt_out596, dt_out597, dt_out598, dt_out599, dt_out600, dt_out601, dt_out602, dt_out603, dt_out604, dt_out605, dt_out606, dt_out607, 
							dt_out608, dt_out609, dt_out610, dt_out611, dt_out612, dt_out613, dt_out614, dt_out615, dt_out616, dt_out617, dt_out618, dt_out619, dt_out620, dt_out621, dt_out622, dt_out623, 
							dt_out624, dt_out625, dt_out626, dt_out627, dt_out628, dt_out629, dt_out630, dt_out631, dt_out632, dt_out633, dt_out634, dt_out635, dt_out636, dt_out637, dt_out638, dt_out639, 
							dt_out640, dt_out641, dt_out642, dt_out643, dt_out644, dt_out645, dt_out646, dt_out647, dt_out648, dt_out649, dt_out650, dt_out651, dt_out652, dt_out653, dt_out654, dt_out655, 
							dt_out656, dt_out657, dt_out658, dt_out659, dt_out660, dt_out661, dt_out662, dt_out663, dt_out664, dt_out665, dt_out666, dt_out667, dt_out668, dt_out669, dt_out670, dt_out671, 
							dt_out672, dt_out673, dt_out674, dt_out675, dt_out676, dt_out677, dt_out678, dt_out679, dt_out680, dt_out681, dt_out682, dt_out683, dt_out684, dt_out685, dt_out686, dt_out687, 
							dt_out688, dt_out689, dt_out690, dt_out691, dt_out692, dt_out693, dt_out694, dt_out695, dt_out696, dt_out697, dt_out698, dt_out699, dt_out700, dt_out701, dt_out702, dt_out703, 
							dt_out704, dt_out705, dt_out706, dt_out707, dt_out708, dt_out709, dt_out710, dt_out711, dt_out712, dt_out713, dt_out714, dt_out715, dt_out716, dt_out717, dt_out718, dt_out719, 
							dt_out720, dt_out721, dt_out722, dt_out723, dt_out724, dt_out725, dt_out726, dt_out727, dt_out728, dt_out729, dt_out730, dt_out731, dt_out732, dt_out733, dt_out734, dt_out735, 
							dt_out736, dt_out737, dt_out738, dt_out739, dt_out740, dt_out741, dt_out742, dt_out743, dt_out744, dt_out745, dt_out746, dt_out747, dt_out748, dt_out749, dt_out750, dt_out751, 
							dt_out752, dt_out753, dt_out754, dt_out755, dt_out756, dt_out757, dt_out758, dt_out759, dt_out760, dt_out761, dt_out762, dt_out763, dt_out764, dt_out765, dt_out766, dt_out767, 
							dt_out768, dt_out769, dt_out770, dt_out771, dt_out772, dt_out773, dt_out774, dt_out775, dt_out776, dt_out777, dt_out778, dt_out779, dt_out780, dt_out781, dt_out782, dt_out783, 
							dt_out784, dt_out785, dt_out786, dt_out787, dt_out788, dt_out789, dt_out790, dt_out791, dt_out792, dt_out793, dt_out794, dt_out795, dt_out796, dt_out797, dt_out798, dt_out799, 
							dt_out800, dt_out801, dt_out802, dt_out803, dt_out804, dt_out805, dt_out806, dt_out807, dt_out808, dt_out809, dt_out810, dt_out811, dt_out812, dt_out813, dt_out814, dt_out815, 
							dt_out816, dt_out817, dt_out818, dt_out819, dt_out820, dt_out821, dt_out822, dt_out823, dt_out824, dt_out825, dt_out826, dt_out827, dt_out828, dt_out829, dt_out830, dt_out831, 
							dt_out832, dt_out833, dt_out834, dt_out835, dt_out836, dt_out837, dt_out838, dt_out839, dt_out840, dt_out841, dt_out842, dt_out843, dt_out844, dt_out845, dt_out846, dt_out847, 
							dt_out848, dt_out849, dt_out850, dt_out851, dt_out852, dt_out853, dt_out854, dt_out855, dt_out856, dt_out857, dt_out858, dt_out859, dt_out860, dt_out861, dt_out862, dt_out863, 
							dt_out864, dt_out865, dt_out866, dt_out867, dt_out868, dt_out869, dt_out870, dt_out871, dt_out872, dt_out873, dt_out874, dt_out875, dt_out876, dt_out877, dt_out878, dt_out879, 
							dt_out880, dt_out881, dt_out882, dt_out883, dt_out884, dt_out885, dt_out886, dt_out887, dt_out888, dt_out889, dt_out890, dt_out891, dt_out892, dt_out893, dt_out894, dt_out895, 
							dt_out896, dt_out897, dt_out898, dt_out899, dt_out900, dt_out901, dt_out902, dt_out903, dt_out904, dt_out905, dt_out906, dt_out907, dt_out908, dt_out909, dt_out910, dt_out911, 
							dt_out912, dt_out913, dt_out914, dt_out915, dt_out916, dt_out917, dt_out918, dt_out919, dt_out920, dt_out921, dt_out922, dt_out923, dt_out924, dt_out925, dt_out926, dt_out927, 
							dt_out928, dt_out929, dt_out930, dt_out931, dt_out932, dt_out933, dt_out934, dt_out935, dt_out936, dt_out937, dt_out938, dt_out939, dt_out940, dt_out941, dt_out942, dt_out943, 
							dt_out944, dt_out945, dt_out946, dt_out947, dt_out948, dt_out949, dt_out950, dt_out951, dt_out952, dt_out953, dt_out954, dt_out955, dt_out956, dt_out957, dt_out958, dt_out959, 
							dt_out960, dt_out961, dt_out962, dt_out963, dt_out964, dt_out965, dt_out966, dt_out967, dt_out968, dt_out969, dt_out970, dt_out971, dt_out972, dt_out973, dt_out974, dt_out975, 
							dt_out976, dt_out977, dt_out978, dt_out979, dt_out980, dt_out981, dt_out982, dt_out983, dt_out984, dt_out985, dt_out986, dt_out987, dt_out988, dt_out989, dt_out990, dt_out991, 
							dt_out992, dt_out993, dt_out994, dt_out995, dt_out996, dt_out997, dt_out998, dt_out999, dt_out1000, dt_out1001, dt_out1002, dt_out1003, dt_out1004, dt_out1005, dt_out1006, dt_out1007, 
							dt_out1008, dt_out1009, dt_out1010, dt_out1011, dt_out1012, dt_out1013, dt_out1014, dt_out1015, dt_out1016, dt_out1017, dt_out1018, dt_out1019, dt_out1020, dt_out1021, dt_out1022, dt_out1023);

	always @(posedge clk or negedge n_stall_out) begin
		if (!n_stall_out && cur_cycle > `LOG2(4)+4) begin	
			`ifdef GEN_VCD
				$display ("WARNS --- Generate VCD file !");
				`ifdef MODELSIM						// defined in <designs.h> file
					$dumpflush;
					$dumpoff;
				`elsif VCS
					$vcdplusflush;
					$vcdplusoff;
				`else
					$display ("ERROR --- Simulation tool is not supported (ModelSim or Synopsys VCS");
				`endif
			`else
				$display ("WARNS --- No VCD file is generated !");
			`endif
			$display ("INFOR --- Simulation is finished at cycle   %d", cur_cycle);
			$display ("INFOR --- CLOCK_PERIOD:                          %.3f", `CLOCK_PERIOD); 

			//$stop;
			$finish;
		end
	end

	// clock generator
		vcClockGen	 #(.clockperiod(`CLOCK_PERIOD)) 
			inst_vcClockGen(.clk(clk), .n_clk(n_clk), .n_rst(n_rst), .cur_cycle(cur_cycle));

	// start generating VCD file for power estimation
		initial
  		begin  			
			`ifdef GEN_VCD
				$dumpfile(`VCD_FILE);
				$dumpvars(0, dut_adder);			// dump all variables inside dut_fft4 into VCD file

				`ifdef MODELSIM
					$display ("INFOR --- Using ModelSim simulator");
				`elsif VCS
					$display ("INFOR --- Using Synopsys VCS simulator");
					$vcdpluson;
				`else
					$display ("ERROR --- Simulation tool is not supported (ModelSim or Synopsys VCS)");
				`endif				
			`endif
		end

	// FIFO
		fifo #(.depth(2)) inst_fifo(.clk(n_clk), .n_rst(n_rst), .n_stall_in(n_stall), .n_stall_out(n_stall_out));

	// Design Under Test
		adder dut_adder(.clk(n_clk), .n_rst(n_rst), .n_stall(n_stall),
						  .a0(dt_in0), .b0(dt_in1), .a1(dt_in2), .b1(dt_in3), .out0(dt_out0), .out1(dt_out1));

endmodule