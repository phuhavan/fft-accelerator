`include "macros.h"

module fft2048
#(
		//--- data bit-width
			parameter width = 24,
		//--- fft size
			parameter size=2048
)
(
		//--- control
			input                   clk, rst, stall,              
		//--- inputs
			input    [width-1:0]    x0_in,                        
			input    [width-1:0]    x1_in,                        
			input    [width-1:0]    x2_in,                        
			input    [width-1:0]    x3_in,                        
			input    [width-1:0]    x4_in,                        
			input    [width-1:0]    x5_in,                        
			input    [width-1:0]    x6_in,                        
			input    [width-1:0]    x7_in,                        
			input    [width-1:0]    x8_in,                        
			input    [width-1:0]    x9_in,                        
			input    [width-1:0]    x10_in,                       
			input    [width-1:0]    x11_in,                       
			input    [width-1:0]    x12_in,                       
			input    [width-1:0]    x13_in,                       
			input    [width-1:0]    x14_in,                       
			input    [width-1:0]    x15_in,                       
			input    [width-1:0]    x16_in,                       
			input    [width-1:0]    x17_in,                       
			input    [width-1:0]    x18_in,                       
			input    [width-1:0]    x19_in,                       
			input    [width-1:0]    x20_in,                       
			input    [width-1:0]    x21_in,                       
			input    [width-1:0]    x22_in,                       
			input    [width-1:0]    x23_in,                       
			input    [width-1:0]    x24_in,                       
			input    [width-1:0]    x25_in,                       
			input    [width-1:0]    x26_in,                       
			input    [width-1:0]    x27_in,                       
			input    [width-1:0]    x28_in,                       
			input    [width-1:0]    x29_in,                       
			input    [width-1:0]    x30_in,                       
			input    [width-1:0]    x31_in,                       
			input    [width-1:0]    x32_in,                       
			input    [width-1:0]    x33_in,                       
			input    [width-1:0]    x34_in,                       
			input    [width-1:0]    x35_in,                       
			input    [width-1:0]    x36_in,                       
			input    [width-1:0]    x37_in,                       
			input    [width-1:0]    x38_in,                       
			input    [width-1:0]    x39_in,                       
			input    [width-1:0]    x40_in,                       
			input    [width-1:0]    x41_in,                       
			input    [width-1:0]    x42_in,                       
			input    [width-1:0]    x43_in,                       
			input    [width-1:0]    x44_in,                       
			input    [width-1:0]    x45_in,                       
			input    [width-1:0]    x46_in,                       
			input    [width-1:0]    x47_in,                       
			input    [width-1:0]    x48_in,                       
			input    [width-1:0]    x49_in,                       
			input    [width-1:0]    x50_in,                       
			input    [width-1:0]    x51_in,                       
			input    [width-1:0]    x52_in,                       
			input    [width-1:0]    x53_in,                       
			input    [width-1:0]    x54_in,                       
			input    [width-1:0]    x55_in,                       
			input    [width-1:0]    x56_in,                       
			input    [width-1:0]    x57_in,                       
			input    [width-1:0]    x58_in,                       
			input    [width-1:0]    x59_in,                       
			input    [width-1:0]    x60_in,                       
			input    [width-1:0]    x61_in,                       
			input    [width-1:0]    x62_in,                       
			input    [width-1:0]    x63_in,                       
			input    [width-1:0]    x64_in,                       
			input    [width-1:0]    x65_in,                       
			input    [width-1:0]    x66_in,                       
			input    [width-1:0]    x67_in,                       
			input    [width-1:0]    x68_in,                       
			input    [width-1:0]    x69_in,                       
			input    [width-1:0]    x70_in,                       
			input    [width-1:0]    x71_in,                       
			input    [width-1:0]    x72_in,                       
			input    [width-1:0]    x73_in,                       
			input    [width-1:0]    x74_in,                       
			input    [width-1:0]    x75_in,                       
			input    [width-1:0]    x76_in,                       
			input    [width-1:0]    x77_in,                       
			input    [width-1:0]    x78_in,                       
			input    [width-1:0]    x79_in,                       
			input    [width-1:0]    x80_in,                       
			input    [width-1:0]    x81_in,                       
			input    [width-1:0]    x82_in,                       
			input    [width-1:0]    x83_in,                       
			input    [width-1:0]    x84_in,                       
			input    [width-1:0]    x85_in,                       
			input    [width-1:0]    x86_in,                       
			input    [width-1:0]    x87_in,                       
			input    [width-1:0]    x88_in,                       
			input    [width-1:0]    x89_in,                       
			input    [width-1:0]    x90_in,                       
			input    [width-1:0]    x91_in,                       
			input    [width-1:0]    x92_in,                       
			input    [width-1:0]    x93_in,                       
			input    [width-1:0]    x94_in,                       
			input    [width-1:0]    x95_in,                       
			input    [width-1:0]    x96_in,                       
			input    [width-1:0]    x97_in,                       
			input    [width-1:0]    x98_in,                       
			input    [width-1:0]    x99_in,                       
			input    [width-1:0]    x100_in,                      
			input    [width-1:0]    x101_in,                      
			input    [width-1:0]    x102_in,                      
			input    [width-1:0]    x103_in,                      
			input    [width-1:0]    x104_in,                      
			input    [width-1:0]    x105_in,                      
			input    [width-1:0]    x106_in,                      
			input    [width-1:0]    x107_in,                      
			input    [width-1:0]    x108_in,                      
			input    [width-1:0]    x109_in,                      
			input    [width-1:0]    x110_in,                      
			input    [width-1:0]    x111_in,                      
			input    [width-1:0]    x112_in,                      
			input    [width-1:0]    x113_in,                      
			input    [width-1:0]    x114_in,                      
			input    [width-1:0]    x115_in,                      
			input    [width-1:0]    x116_in,                      
			input    [width-1:0]    x117_in,                      
			input    [width-1:0]    x118_in,                      
			input    [width-1:0]    x119_in,                      
			input    [width-1:0]    x120_in,                      
			input    [width-1:0]    x121_in,                      
			input    [width-1:0]    x122_in,                      
			input    [width-1:0]    x123_in,                      
			input    [width-1:0]    x124_in,                      
			input    [width-1:0]    x125_in,                      
			input    [width-1:0]    x126_in,                      
			input    [width-1:0]    x127_in,                      
			input    [width-1:0]    x128_in,                      
			input    [width-1:0]    x129_in,                      
			input    [width-1:0]    x130_in,                      
			input    [width-1:0]    x131_in,                      
			input    [width-1:0]    x132_in,                      
			input    [width-1:0]    x133_in,                      
			input    [width-1:0]    x134_in,                      
			input    [width-1:0]    x135_in,                      
			input    [width-1:0]    x136_in,                      
			input    [width-1:0]    x137_in,                      
			input    [width-1:0]    x138_in,                      
			input    [width-1:0]    x139_in,                      
			input    [width-1:0]    x140_in,                      
			input    [width-1:0]    x141_in,                      
			input    [width-1:0]    x142_in,                      
			input    [width-1:0]    x143_in,                      
			input    [width-1:0]    x144_in,                      
			input    [width-1:0]    x145_in,                      
			input    [width-1:0]    x146_in,                      
			input    [width-1:0]    x147_in,                      
			input    [width-1:0]    x148_in,                      
			input    [width-1:0]    x149_in,                      
			input    [width-1:0]    x150_in,                      
			input    [width-1:0]    x151_in,                      
			input    [width-1:0]    x152_in,                      
			input    [width-1:0]    x153_in,                      
			input    [width-1:0]    x154_in,                      
			input    [width-1:0]    x155_in,                      
			input    [width-1:0]    x156_in,                      
			input    [width-1:0]    x157_in,                      
			input    [width-1:0]    x158_in,                      
			input    [width-1:0]    x159_in,                      
			input    [width-1:0]    x160_in,                      
			input    [width-1:0]    x161_in,                      
			input    [width-1:0]    x162_in,                      
			input    [width-1:0]    x163_in,                      
			input    [width-1:0]    x164_in,                      
			input    [width-1:0]    x165_in,                      
			input    [width-1:0]    x166_in,                      
			input    [width-1:0]    x167_in,                      
			input    [width-1:0]    x168_in,                      
			input    [width-1:0]    x169_in,                      
			input    [width-1:0]    x170_in,                      
			input    [width-1:0]    x171_in,                      
			input    [width-1:0]    x172_in,                      
			input    [width-1:0]    x173_in,                      
			input    [width-1:0]    x174_in,                      
			input    [width-1:0]    x175_in,                      
			input    [width-1:0]    x176_in,                      
			input    [width-1:0]    x177_in,                      
			input    [width-1:0]    x178_in,                      
			input    [width-1:0]    x179_in,                      
			input    [width-1:0]    x180_in,                      
			input    [width-1:0]    x181_in,                      
			input    [width-1:0]    x182_in,                      
			input    [width-1:0]    x183_in,                      
			input    [width-1:0]    x184_in,                      
			input    [width-1:0]    x185_in,                      
			input    [width-1:0]    x186_in,                      
			input    [width-1:0]    x187_in,                      
			input    [width-1:0]    x188_in,                      
			input    [width-1:0]    x189_in,                      
			input    [width-1:0]    x190_in,                      
			input    [width-1:0]    x191_in,                      
			input    [width-1:0]    x192_in,                      
			input    [width-1:0]    x193_in,                      
			input    [width-1:0]    x194_in,                      
			input    [width-1:0]    x195_in,                      
			input    [width-1:0]    x196_in,                      
			input    [width-1:0]    x197_in,                      
			input    [width-1:0]    x198_in,                      
			input    [width-1:0]    x199_in,                      
			input    [width-1:0]    x200_in,                      
			input    [width-1:0]    x201_in,                      
			input    [width-1:0]    x202_in,                      
			input    [width-1:0]    x203_in,                      
			input    [width-1:0]    x204_in,                      
			input    [width-1:0]    x205_in,                      
			input    [width-1:0]    x206_in,                      
			input    [width-1:0]    x207_in,                      
			input    [width-1:0]    x208_in,                      
			input    [width-1:0]    x209_in,                      
			input    [width-1:0]    x210_in,                      
			input    [width-1:0]    x211_in,                      
			input    [width-1:0]    x212_in,                      
			input    [width-1:0]    x213_in,                      
			input    [width-1:0]    x214_in,                      
			input    [width-1:0]    x215_in,                      
			input    [width-1:0]    x216_in,                      
			input    [width-1:0]    x217_in,                      
			input    [width-1:0]    x218_in,                      
			input    [width-1:0]    x219_in,                      
			input    [width-1:0]    x220_in,                      
			input    [width-1:0]    x221_in,                      
			input    [width-1:0]    x222_in,                      
			input    [width-1:0]    x223_in,                      
			input    [width-1:0]    x224_in,                      
			input    [width-1:0]    x225_in,                      
			input    [width-1:0]    x226_in,                      
			input    [width-1:0]    x227_in,                      
			input    [width-1:0]    x228_in,                      
			input    [width-1:0]    x229_in,                      
			input    [width-1:0]    x230_in,                      
			input    [width-1:0]    x231_in,                      
			input    [width-1:0]    x232_in,                      
			input    [width-1:0]    x233_in,                      
			input    [width-1:0]    x234_in,                      
			input    [width-1:0]    x235_in,                      
			input    [width-1:0]    x236_in,                      
			input    [width-1:0]    x237_in,                      
			input    [width-1:0]    x238_in,                      
			input    [width-1:0]    x239_in,                      
			input    [width-1:0]    x240_in,                      
			input    [width-1:0]    x241_in,                      
			input    [width-1:0]    x242_in,                      
			input    [width-1:0]    x243_in,                      
			input    [width-1:0]    x244_in,                      
			input    [width-1:0]    x245_in,                      
			input    [width-1:0]    x246_in,                      
			input    [width-1:0]    x247_in,                      
			input    [width-1:0]    x248_in,                      
			input    [width-1:0]    x249_in,                      
			input    [width-1:0]    x250_in,                      
			input    [width-1:0]    x251_in,                      
			input    [width-1:0]    x252_in,                      
			input    [width-1:0]    x253_in,                      
			input    [width-1:0]    x254_in,                      
			input    [width-1:0]    x255_in,                      
			input    [width-1:0]    x256_in,                      
			input    [width-1:0]    x257_in,                      
			input    [width-1:0]    x258_in,                      
			input    [width-1:0]    x259_in,                      
			input    [width-1:0]    x260_in,                      
			input    [width-1:0]    x261_in,                      
			input    [width-1:0]    x262_in,                      
			input    [width-1:0]    x263_in,                      
			input    [width-1:0]    x264_in,                      
			input    [width-1:0]    x265_in,                      
			input    [width-1:0]    x266_in,                      
			input    [width-1:0]    x267_in,                      
			input    [width-1:0]    x268_in,                      
			input    [width-1:0]    x269_in,                      
			input    [width-1:0]    x270_in,                      
			input    [width-1:0]    x271_in,                      
			input    [width-1:0]    x272_in,                      
			input    [width-1:0]    x273_in,                      
			input    [width-1:0]    x274_in,                      
			input    [width-1:0]    x275_in,                      
			input    [width-1:0]    x276_in,                      
			input    [width-1:0]    x277_in,                      
			input    [width-1:0]    x278_in,                      
			input    [width-1:0]    x279_in,                      
			input    [width-1:0]    x280_in,                      
			input    [width-1:0]    x281_in,                      
			input    [width-1:0]    x282_in,                      
			input    [width-1:0]    x283_in,                      
			input    [width-1:0]    x284_in,                      
			input    [width-1:0]    x285_in,                      
			input    [width-1:0]    x286_in,                      
			input    [width-1:0]    x287_in,                      
			input    [width-1:0]    x288_in,                      
			input    [width-1:0]    x289_in,                      
			input    [width-1:0]    x290_in,                      
			input    [width-1:0]    x291_in,                      
			input    [width-1:0]    x292_in,                      
			input    [width-1:0]    x293_in,                      
			input    [width-1:0]    x294_in,                      
			input    [width-1:0]    x295_in,                      
			input    [width-1:0]    x296_in,                      
			input    [width-1:0]    x297_in,                      
			input    [width-1:0]    x298_in,                      
			input    [width-1:0]    x299_in,                      
			input    [width-1:0]    x300_in,                      
			input    [width-1:0]    x301_in,                      
			input    [width-1:0]    x302_in,                      
			input    [width-1:0]    x303_in,                      
			input    [width-1:0]    x304_in,                      
			input    [width-1:0]    x305_in,                      
			input    [width-1:0]    x306_in,                      
			input    [width-1:0]    x307_in,                      
			input    [width-1:0]    x308_in,                      
			input    [width-1:0]    x309_in,                      
			input    [width-1:0]    x310_in,                      
			input    [width-1:0]    x311_in,                      
			input    [width-1:0]    x312_in,                      
			input    [width-1:0]    x313_in,                      
			input    [width-1:0]    x314_in,                      
			input    [width-1:0]    x315_in,                      
			input    [width-1:0]    x316_in,                      
			input    [width-1:0]    x317_in,                      
			input    [width-1:0]    x318_in,                      
			input    [width-1:0]    x319_in,                      
			input    [width-1:0]    x320_in,                      
			input    [width-1:0]    x321_in,                      
			input    [width-1:0]    x322_in,                      
			input    [width-1:0]    x323_in,                      
			input    [width-1:0]    x324_in,                      
			input    [width-1:0]    x325_in,                      
			input    [width-1:0]    x326_in,                      
			input    [width-1:0]    x327_in,                      
			input    [width-1:0]    x328_in,                      
			input    [width-1:0]    x329_in,                      
			input    [width-1:0]    x330_in,                      
			input    [width-1:0]    x331_in,                      
			input    [width-1:0]    x332_in,                      
			input    [width-1:0]    x333_in,                      
			input    [width-1:0]    x334_in,                      
			input    [width-1:0]    x335_in,                      
			input    [width-1:0]    x336_in,                      
			input    [width-1:0]    x337_in,                      
			input    [width-1:0]    x338_in,                      
			input    [width-1:0]    x339_in,                      
			input    [width-1:0]    x340_in,                      
			input    [width-1:0]    x341_in,                      
			input    [width-1:0]    x342_in,                      
			input    [width-1:0]    x343_in,                      
			input    [width-1:0]    x344_in,                      
			input    [width-1:0]    x345_in,                      
			input    [width-1:0]    x346_in,                      
			input    [width-1:0]    x347_in,                      
			input    [width-1:0]    x348_in,                      
			input    [width-1:0]    x349_in,                      
			input    [width-1:0]    x350_in,                      
			input    [width-1:0]    x351_in,                      
			input    [width-1:0]    x352_in,                      
			input    [width-1:0]    x353_in,                      
			input    [width-1:0]    x354_in,                      
			input    [width-1:0]    x355_in,                      
			input    [width-1:0]    x356_in,                      
			input    [width-1:0]    x357_in,                      
			input    [width-1:0]    x358_in,                      
			input    [width-1:0]    x359_in,                      
			input    [width-1:0]    x360_in,                      
			input    [width-1:0]    x361_in,                      
			input    [width-1:0]    x362_in,                      
			input    [width-1:0]    x363_in,                      
			input    [width-1:0]    x364_in,                      
			input    [width-1:0]    x365_in,                      
			input    [width-1:0]    x366_in,                      
			input    [width-1:0]    x367_in,                      
			input    [width-1:0]    x368_in,                      
			input    [width-1:0]    x369_in,                      
			input    [width-1:0]    x370_in,                      
			input    [width-1:0]    x371_in,                      
			input    [width-1:0]    x372_in,                      
			input    [width-1:0]    x373_in,                      
			input    [width-1:0]    x374_in,                      
			input    [width-1:0]    x375_in,                      
			input    [width-1:0]    x376_in,                      
			input    [width-1:0]    x377_in,                      
			input    [width-1:0]    x378_in,                      
			input    [width-1:0]    x379_in,                      
			input    [width-1:0]    x380_in,                      
			input    [width-1:0]    x381_in,                      
			input    [width-1:0]    x382_in,                      
			input    [width-1:0]    x383_in,                      
			input    [width-1:0]    x384_in,                      
			input    [width-1:0]    x385_in,                      
			input    [width-1:0]    x386_in,                      
			input    [width-1:0]    x387_in,                      
			input    [width-1:0]    x388_in,                      
			input    [width-1:0]    x389_in,                      
			input    [width-1:0]    x390_in,                      
			input    [width-1:0]    x391_in,                      
			input    [width-1:0]    x392_in,                      
			input    [width-1:0]    x393_in,                      
			input    [width-1:0]    x394_in,                      
			input    [width-1:0]    x395_in,                      
			input    [width-1:0]    x396_in,                      
			input    [width-1:0]    x397_in,                      
			input    [width-1:0]    x398_in,                      
			input    [width-1:0]    x399_in,                      
			input    [width-1:0]    x400_in,                      
			input    [width-1:0]    x401_in,                      
			input    [width-1:0]    x402_in,                      
			input    [width-1:0]    x403_in,                      
			input    [width-1:0]    x404_in,                      
			input    [width-1:0]    x405_in,                      
			input    [width-1:0]    x406_in,                      
			input    [width-1:0]    x407_in,                      
			input    [width-1:0]    x408_in,                      
			input    [width-1:0]    x409_in,                      
			input    [width-1:0]    x410_in,                      
			input    [width-1:0]    x411_in,                      
			input    [width-1:0]    x412_in,                      
			input    [width-1:0]    x413_in,                      
			input    [width-1:0]    x414_in,                      
			input    [width-1:0]    x415_in,                      
			input    [width-1:0]    x416_in,                      
			input    [width-1:0]    x417_in,                      
			input    [width-1:0]    x418_in,                      
			input    [width-1:0]    x419_in,                      
			input    [width-1:0]    x420_in,                      
			input    [width-1:0]    x421_in,                      
			input    [width-1:0]    x422_in,                      
			input    [width-1:0]    x423_in,                      
			input    [width-1:0]    x424_in,                      
			input    [width-1:0]    x425_in,                      
			input    [width-1:0]    x426_in,                      
			input    [width-1:0]    x427_in,                      
			input    [width-1:0]    x428_in,                      
			input    [width-1:0]    x429_in,                      
			input    [width-1:0]    x430_in,                      
			input    [width-1:0]    x431_in,                      
			input    [width-1:0]    x432_in,                      
			input    [width-1:0]    x433_in,                      
			input    [width-1:0]    x434_in,                      
			input    [width-1:0]    x435_in,                      
			input    [width-1:0]    x436_in,                      
			input    [width-1:0]    x437_in,                      
			input    [width-1:0]    x438_in,                      
			input    [width-1:0]    x439_in,                      
			input    [width-1:0]    x440_in,                      
			input    [width-1:0]    x441_in,                      
			input    [width-1:0]    x442_in,                      
			input    [width-1:0]    x443_in,                      
			input    [width-1:0]    x444_in,                      
			input    [width-1:0]    x445_in,                      
			input    [width-1:0]    x446_in,                      
			input    [width-1:0]    x447_in,                      
			input    [width-1:0]    x448_in,                      
			input    [width-1:0]    x449_in,                      
			input    [width-1:0]    x450_in,                      
			input    [width-1:0]    x451_in,                      
			input    [width-1:0]    x452_in,                      
			input    [width-1:0]    x453_in,                      
			input    [width-1:0]    x454_in,                      
			input    [width-1:0]    x455_in,                      
			input    [width-1:0]    x456_in,                      
			input    [width-1:0]    x457_in,                      
			input    [width-1:0]    x458_in,                      
			input    [width-1:0]    x459_in,                      
			input    [width-1:0]    x460_in,                      
			input    [width-1:0]    x461_in,                      
			input    [width-1:0]    x462_in,                      
			input    [width-1:0]    x463_in,                      
			input    [width-1:0]    x464_in,                      
			input    [width-1:0]    x465_in,                      
			input    [width-1:0]    x466_in,                      
			input    [width-1:0]    x467_in,                      
			input    [width-1:0]    x468_in,                      
			input    [width-1:0]    x469_in,                      
			input    [width-1:0]    x470_in,                      
			input    [width-1:0]    x471_in,                      
			input    [width-1:0]    x472_in,                      
			input    [width-1:0]    x473_in,                      
			input    [width-1:0]    x474_in,                      
			input    [width-1:0]    x475_in,                      
			input    [width-1:0]    x476_in,                      
			input    [width-1:0]    x477_in,                      
			input    [width-1:0]    x478_in,                      
			input    [width-1:0]    x479_in,                      
			input    [width-1:0]    x480_in,                      
			input    [width-1:0]    x481_in,                      
			input    [width-1:0]    x482_in,                      
			input    [width-1:0]    x483_in,                      
			input    [width-1:0]    x484_in,                      
			input    [width-1:0]    x485_in,                      
			input    [width-1:0]    x486_in,                      
			input    [width-1:0]    x487_in,                      
			input    [width-1:0]    x488_in,                      
			input    [width-1:0]    x489_in,                      
			input    [width-1:0]    x490_in,                      
			input    [width-1:0]    x491_in,                      
			input    [width-1:0]    x492_in,                      
			input    [width-1:0]    x493_in,                      
			input    [width-1:0]    x494_in,                      
			input    [width-1:0]    x495_in,                      
			input    [width-1:0]    x496_in,                      
			input    [width-1:0]    x497_in,                      
			input    [width-1:0]    x498_in,                      
			input    [width-1:0]    x499_in,                      
			input    [width-1:0]    x500_in,                      
			input    [width-1:0]    x501_in,                      
			input    [width-1:0]    x502_in,                      
			input    [width-1:0]    x503_in,                      
			input    [width-1:0]    x504_in,                      
			input    [width-1:0]    x505_in,                      
			input    [width-1:0]    x506_in,                      
			input    [width-1:0]    x507_in,                      
			input    [width-1:0]    x508_in,                      
			input    [width-1:0]    x509_in,                      
			input    [width-1:0]    x510_in,                      
			input    [width-1:0]    x511_in,                      
			input    [width-1:0]    x512_in,                      
			input    [width-1:0]    x513_in,                      
			input    [width-1:0]    x514_in,                      
			input    [width-1:0]    x515_in,                      
			input    [width-1:0]    x516_in,                      
			input    [width-1:0]    x517_in,                      
			input    [width-1:0]    x518_in,                      
			input    [width-1:0]    x519_in,                      
			input    [width-1:0]    x520_in,                      
			input    [width-1:0]    x521_in,                      
			input    [width-1:0]    x522_in,                      
			input    [width-1:0]    x523_in,                      
			input    [width-1:0]    x524_in,                      
			input    [width-1:0]    x525_in,                      
			input    [width-1:0]    x526_in,                      
			input    [width-1:0]    x527_in,                      
			input    [width-1:0]    x528_in,                      
			input    [width-1:0]    x529_in,                      
			input    [width-1:0]    x530_in,                      
			input    [width-1:0]    x531_in,                      
			input    [width-1:0]    x532_in,                      
			input    [width-1:0]    x533_in,                      
			input    [width-1:0]    x534_in,                      
			input    [width-1:0]    x535_in,                      
			input    [width-1:0]    x536_in,                      
			input    [width-1:0]    x537_in,                      
			input    [width-1:0]    x538_in,                      
			input    [width-1:0]    x539_in,                      
			input    [width-1:0]    x540_in,                      
			input    [width-1:0]    x541_in,                      
			input    [width-1:0]    x542_in,                      
			input    [width-1:0]    x543_in,                      
			input    [width-1:0]    x544_in,                      
			input    [width-1:0]    x545_in,                      
			input    [width-1:0]    x546_in,                      
			input    [width-1:0]    x547_in,                      
			input    [width-1:0]    x548_in,                      
			input    [width-1:0]    x549_in,                      
			input    [width-1:0]    x550_in,                      
			input    [width-1:0]    x551_in,                      
			input    [width-1:0]    x552_in,                      
			input    [width-1:0]    x553_in,                      
			input    [width-1:0]    x554_in,                      
			input    [width-1:0]    x555_in,                      
			input    [width-1:0]    x556_in,                      
			input    [width-1:0]    x557_in,                      
			input    [width-1:0]    x558_in,                      
			input    [width-1:0]    x559_in,                      
			input    [width-1:0]    x560_in,                      
			input    [width-1:0]    x561_in,                      
			input    [width-1:0]    x562_in,                      
			input    [width-1:0]    x563_in,                      
			input    [width-1:0]    x564_in,                      
			input    [width-1:0]    x565_in,                      
			input    [width-1:0]    x566_in,                      
			input    [width-1:0]    x567_in,                      
			input    [width-1:0]    x568_in,                      
			input    [width-1:0]    x569_in,                      
			input    [width-1:0]    x570_in,                      
			input    [width-1:0]    x571_in,                      
			input    [width-1:0]    x572_in,                      
			input    [width-1:0]    x573_in,                      
			input    [width-1:0]    x574_in,                      
			input    [width-1:0]    x575_in,                      
			input    [width-1:0]    x576_in,                      
			input    [width-1:0]    x577_in,                      
			input    [width-1:0]    x578_in,                      
			input    [width-1:0]    x579_in,                      
			input    [width-1:0]    x580_in,                      
			input    [width-1:0]    x581_in,                      
			input    [width-1:0]    x582_in,                      
			input    [width-1:0]    x583_in,                      
			input    [width-1:0]    x584_in,                      
			input    [width-1:0]    x585_in,                      
			input    [width-1:0]    x586_in,                      
			input    [width-1:0]    x587_in,                      
			input    [width-1:0]    x588_in,                      
			input    [width-1:0]    x589_in,                      
			input    [width-1:0]    x590_in,                      
			input    [width-1:0]    x591_in,                      
			input    [width-1:0]    x592_in,                      
			input    [width-1:0]    x593_in,                      
			input    [width-1:0]    x594_in,                      
			input    [width-1:0]    x595_in,                      
			input    [width-1:0]    x596_in,                      
			input    [width-1:0]    x597_in,                      
			input    [width-1:0]    x598_in,                      
			input    [width-1:0]    x599_in,                      
			input    [width-1:0]    x600_in,                      
			input    [width-1:0]    x601_in,                      
			input    [width-1:0]    x602_in,                      
			input    [width-1:0]    x603_in,                      
			input    [width-1:0]    x604_in,                      
			input    [width-1:0]    x605_in,                      
			input    [width-1:0]    x606_in,                      
			input    [width-1:0]    x607_in,                      
			input    [width-1:0]    x608_in,                      
			input    [width-1:0]    x609_in,                      
			input    [width-1:0]    x610_in,                      
			input    [width-1:0]    x611_in,                      
			input    [width-1:0]    x612_in,                      
			input    [width-1:0]    x613_in,                      
			input    [width-1:0]    x614_in,                      
			input    [width-1:0]    x615_in,                      
			input    [width-1:0]    x616_in,                      
			input    [width-1:0]    x617_in,                      
			input    [width-1:0]    x618_in,                      
			input    [width-1:0]    x619_in,                      
			input    [width-1:0]    x620_in,                      
			input    [width-1:0]    x621_in,                      
			input    [width-1:0]    x622_in,                      
			input    [width-1:0]    x623_in,                      
			input    [width-1:0]    x624_in,                      
			input    [width-1:0]    x625_in,                      
			input    [width-1:0]    x626_in,                      
			input    [width-1:0]    x627_in,                      
			input    [width-1:0]    x628_in,                      
			input    [width-1:0]    x629_in,                      
			input    [width-1:0]    x630_in,                      
			input    [width-1:0]    x631_in,                      
			input    [width-1:0]    x632_in,                      
			input    [width-1:0]    x633_in,                      
			input    [width-1:0]    x634_in,                      
			input    [width-1:0]    x635_in,                      
			input    [width-1:0]    x636_in,                      
			input    [width-1:0]    x637_in,                      
			input    [width-1:0]    x638_in,                      
			input    [width-1:0]    x639_in,                      
			input    [width-1:0]    x640_in,                      
			input    [width-1:0]    x641_in,                      
			input    [width-1:0]    x642_in,                      
			input    [width-1:0]    x643_in,                      
			input    [width-1:0]    x644_in,                      
			input    [width-1:0]    x645_in,                      
			input    [width-1:0]    x646_in,                      
			input    [width-1:0]    x647_in,                      
			input    [width-1:0]    x648_in,                      
			input    [width-1:0]    x649_in,                      
			input    [width-1:0]    x650_in,                      
			input    [width-1:0]    x651_in,                      
			input    [width-1:0]    x652_in,                      
			input    [width-1:0]    x653_in,                      
			input    [width-1:0]    x654_in,                      
			input    [width-1:0]    x655_in,                      
			input    [width-1:0]    x656_in,                      
			input    [width-1:0]    x657_in,                      
			input    [width-1:0]    x658_in,                      
			input    [width-1:0]    x659_in,                      
			input    [width-1:0]    x660_in,                      
			input    [width-1:0]    x661_in,                      
			input    [width-1:0]    x662_in,                      
			input    [width-1:0]    x663_in,                      
			input    [width-1:0]    x664_in,                      
			input    [width-1:0]    x665_in,                      
			input    [width-1:0]    x666_in,                      
			input    [width-1:0]    x667_in,                      
			input    [width-1:0]    x668_in,                      
			input    [width-1:0]    x669_in,                      
			input    [width-1:0]    x670_in,                      
			input    [width-1:0]    x671_in,                      
			input    [width-1:0]    x672_in,                      
			input    [width-1:0]    x673_in,                      
			input    [width-1:0]    x674_in,                      
			input    [width-1:0]    x675_in,                      
			input    [width-1:0]    x676_in,                      
			input    [width-1:0]    x677_in,                      
			input    [width-1:0]    x678_in,                      
			input    [width-1:0]    x679_in,                      
			input    [width-1:0]    x680_in,                      
			input    [width-1:0]    x681_in,                      
			input    [width-1:0]    x682_in,                      
			input    [width-1:0]    x683_in,                      
			input    [width-1:0]    x684_in,                      
			input    [width-1:0]    x685_in,                      
			input    [width-1:0]    x686_in,                      
			input    [width-1:0]    x687_in,                      
			input    [width-1:0]    x688_in,                      
			input    [width-1:0]    x689_in,                      
			input    [width-1:0]    x690_in,                      
			input    [width-1:0]    x691_in,                      
			input    [width-1:0]    x692_in,                      
			input    [width-1:0]    x693_in,                      
			input    [width-1:0]    x694_in,                      
			input    [width-1:0]    x695_in,                      
			input    [width-1:0]    x696_in,                      
			input    [width-1:0]    x697_in,                      
			input    [width-1:0]    x698_in,                      
			input    [width-1:0]    x699_in,                      
			input    [width-1:0]    x700_in,                      
			input    [width-1:0]    x701_in,                      
			input    [width-1:0]    x702_in,                      
			input    [width-1:0]    x703_in,                      
			input    [width-1:0]    x704_in,                      
			input    [width-1:0]    x705_in,                      
			input    [width-1:0]    x706_in,                      
			input    [width-1:0]    x707_in,                      
			input    [width-1:0]    x708_in,                      
			input    [width-1:0]    x709_in,                      
			input    [width-1:0]    x710_in,                      
			input    [width-1:0]    x711_in,                      
			input    [width-1:0]    x712_in,                      
			input    [width-1:0]    x713_in,                      
			input    [width-1:0]    x714_in,                      
			input    [width-1:0]    x715_in,                      
			input    [width-1:0]    x716_in,                      
			input    [width-1:0]    x717_in,                      
			input    [width-1:0]    x718_in,                      
			input    [width-1:0]    x719_in,                      
			input    [width-1:0]    x720_in,                      
			input    [width-1:0]    x721_in,                      
			input    [width-1:0]    x722_in,                      
			input    [width-1:0]    x723_in,                      
			input    [width-1:0]    x724_in,                      
			input    [width-1:0]    x725_in,                      
			input    [width-1:0]    x726_in,                      
			input    [width-1:0]    x727_in,                      
			input    [width-1:0]    x728_in,                      
			input    [width-1:0]    x729_in,                      
			input    [width-1:0]    x730_in,                      
			input    [width-1:0]    x731_in,                      
			input    [width-1:0]    x732_in,                      
			input    [width-1:0]    x733_in,                      
			input    [width-1:0]    x734_in,                      
			input    [width-1:0]    x735_in,                      
			input    [width-1:0]    x736_in,                      
			input    [width-1:0]    x737_in,                      
			input    [width-1:0]    x738_in,                      
			input    [width-1:0]    x739_in,                      
			input    [width-1:0]    x740_in,                      
			input    [width-1:0]    x741_in,                      
			input    [width-1:0]    x742_in,                      
			input    [width-1:0]    x743_in,                      
			input    [width-1:0]    x744_in,                      
			input    [width-1:0]    x745_in,                      
			input    [width-1:0]    x746_in,                      
			input    [width-1:0]    x747_in,                      
			input    [width-1:0]    x748_in,                      
			input    [width-1:0]    x749_in,                      
			input    [width-1:0]    x750_in,                      
			input    [width-1:0]    x751_in,                      
			input    [width-1:0]    x752_in,                      
			input    [width-1:0]    x753_in,                      
			input    [width-1:0]    x754_in,                      
			input    [width-1:0]    x755_in,                      
			input    [width-1:0]    x756_in,                      
			input    [width-1:0]    x757_in,                      
			input    [width-1:0]    x758_in,                      
			input    [width-1:0]    x759_in,                      
			input    [width-1:0]    x760_in,                      
			input    [width-1:0]    x761_in,                      
			input    [width-1:0]    x762_in,                      
			input    [width-1:0]    x763_in,                      
			input    [width-1:0]    x764_in,                      
			input    [width-1:0]    x765_in,                      
			input    [width-1:0]    x766_in,                      
			input    [width-1:0]    x767_in,                      
			input    [width-1:0]    x768_in,                      
			input    [width-1:0]    x769_in,                      
			input    [width-1:0]    x770_in,                      
			input    [width-1:0]    x771_in,                      
			input    [width-1:0]    x772_in,                      
			input    [width-1:0]    x773_in,                      
			input    [width-1:0]    x774_in,                      
			input    [width-1:0]    x775_in,                      
			input    [width-1:0]    x776_in,                      
			input    [width-1:0]    x777_in,                      
			input    [width-1:0]    x778_in,                      
			input    [width-1:0]    x779_in,                      
			input    [width-1:0]    x780_in,                      
			input    [width-1:0]    x781_in,                      
			input    [width-1:0]    x782_in,                      
			input    [width-1:0]    x783_in,                      
			input    [width-1:0]    x784_in,                      
			input    [width-1:0]    x785_in,                      
			input    [width-1:0]    x786_in,                      
			input    [width-1:0]    x787_in,                      
			input    [width-1:0]    x788_in,                      
			input    [width-1:0]    x789_in,                      
			input    [width-1:0]    x790_in,                      
			input    [width-1:0]    x791_in,                      
			input    [width-1:0]    x792_in,                      
			input    [width-1:0]    x793_in,                      
			input    [width-1:0]    x794_in,                      
			input    [width-1:0]    x795_in,                      
			input    [width-1:0]    x796_in,                      
			input    [width-1:0]    x797_in,                      
			input    [width-1:0]    x798_in,                      
			input    [width-1:0]    x799_in,                      
			input    [width-1:0]    x800_in,                      
			input    [width-1:0]    x801_in,                      
			input    [width-1:0]    x802_in,                      
			input    [width-1:0]    x803_in,                      
			input    [width-1:0]    x804_in,                      
			input    [width-1:0]    x805_in,                      
			input    [width-1:0]    x806_in,                      
			input    [width-1:0]    x807_in,                      
			input    [width-1:0]    x808_in,                      
			input    [width-1:0]    x809_in,                      
			input    [width-1:0]    x810_in,                      
			input    [width-1:0]    x811_in,                      
			input    [width-1:0]    x812_in,                      
			input    [width-1:0]    x813_in,                      
			input    [width-1:0]    x814_in,                      
			input    [width-1:0]    x815_in,                      
			input    [width-1:0]    x816_in,                      
			input    [width-1:0]    x817_in,                      
			input    [width-1:0]    x818_in,                      
			input    [width-1:0]    x819_in,                      
			input    [width-1:0]    x820_in,                      
			input    [width-1:0]    x821_in,                      
			input    [width-1:0]    x822_in,                      
			input    [width-1:0]    x823_in,                      
			input    [width-1:0]    x824_in,                      
			input    [width-1:0]    x825_in,                      
			input    [width-1:0]    x826_in,                      
			input    [width-1:0]    x827_in,                      
			input    [width-1:0]    x828_in,                      
			input    [width-1:0]    x829_in,                      
			input    [width-1:0]    x830_in,                      
			input    [width-1:0]    x831_in,                      
			input    [width-1:0]    x832_in,                      
			input    [width-1:0]    x833_in,                      
			input    [width-1:0]    x834_in,                      
			input    [width-1:0]    x835_in,                      
			input    [width-1:0]    x836_in,                      
			input    [width-1:0]    x837_in,                      
			input    [width-1:0]    x838_in,                      
			input    [width-1:0]    x839_in,                      
			input    [width-1:0]    x840_in,                      
			input    [width-1:0]    x841_in,                      
			input    [width-1:0]    x842_in,                      
			input    [width-1:0]    x843_in,                      
			input    [width-1:0]    x844_in,                      
			input    [width-1:0]    x845_in,                      
			input    [width-1:0]    x846_in,                      
			input    [width-1:0]    x847_in,                      
			input    [width-1:0]    x848_in,                      
			input    [width-1:0]    x849_in,                      
			input    [width-1:0]    x850_in,                      
			input    [width-1:0]    x851_in,                      
			input    [width-1:0]    x852_in,                      
			input    [width-1:0]    x853_in,                      
			input    [width-1:0]    x854_in,                      
			input    [width-1:0]    x855_in,                      
			input    [width-1:0]    x856_in,                      
			input    [width-1:0]    x857_in,                      
			input    [width-1:0]    x858_in,                      
			input    [width-1:0]    x859_in,                      
			input    [width-1:0]    x860_in,                      
			input    [width-1:0]    x861_in,                      
			input    [width-1:0]    x862_in,                      
			input    [width-1:0]    x863_in,                      
			input    [width-1:0]    x864_in,                      
			input    [width-1:0]    x865_in,                      
			input    [width-1:0]    x866_in,                      
			input    [width-1:0]    x867_in,                      
			input    [width-1:0]    x868_in,                      
			input    [width-1:0]    x869_in,                      
			input    [width-1:0]    x870_in,                      
			input    [width-1:0]    x871_in,                      
			input    [width-1:0]    x872_in,                      
			input    [width-1:0]    x873_in,                      
			input    [width-1:0]    x874_in,                      
			input    [width-1:0]    x875_in,                      
			input    [width-1:0]    x876_in,                      
			input    [width-1:0]    x877_in,                      
			input    [width-1:0]    x878_in,                      
			input    [width-1:0]    x879_in,                      
			input    [width-1:0]    x880_in,                      
			input    [width-1:0]    x881_in,                      
			input    [width-1:0]    x882_in,                      
			input    [width-1:0]    x883_in,                      
			input    [width-1:0]    x884_in,                      
			input    [width-1:0]    x885_in,                      
			input    [width-1:0]    x886_in,                      
			input    [width-1:0]    x887_in,                      
			input    [width-1:0]    x888_in,                      
			input    [width-1:0]    x889_in,                      
			input    [width-1:0]    x890_in,                      
			input    [width-1:0]    x891_in,                      
			input    [width-1:0]    x892_in,                      
			input    [width-1:0]    x893_in,                      
			input    [width-1:0]    x894_in,                      
			input    [width-1:0]    x895_in,                      
			input    [width-1:0]    x896_in,                      
			input    [width-1:0]    x897_in,                      
			input    [width-1:0]    x898_in,                      
			input    [width-1:0]    x899_in,                      
			input    [width-1:0]    x900_in,                      
			input    [width-1:0]    x901_in,                      
			input    [width-1:0]    x902_in,                      
			input    [width-1:0]    x903_in,                      
			input    [width-1:0]    x904_in,                      
			input    [width-1:0]    x905_in,                      
			input    [width-1:0]    x906_in,                      
			input    [width-1:0]    x907_in,                      
			input    [width-1:0]    x908_in,                      
			input    [width-1:0]    x909_in,                      
			input    [width-1:0]    x910_in,                      
			input    [width-1:0]    x911_in,                      
			input    [width-1:0]    x912_in,                      
			input    [width-1:0]    x913_in,                      
			input    [width-1:0]    x914_in,                      
			input    [width-1:0]    x915_in,                      
			input    [width-1:0]    x916_in,                      
			input    [width-1:0]    x917_in,                      
			input    [width-1:0]    x918_in,                      
			input    [width-1:0]    x919_in,                      
			input    [width-1:0]    x920_in,                      
			input    [width-1:0]    x921_in,                      
			input    [width-1:0]    x922_in,                      
			input    [width-1:0]    x923_in,                      
			input    [width-1:0]    x924_in,                      
			input    [width-1:0]    x925_in,                      
			input    [width-1:0]    x926_in,                      
			input    [width-1:0]    x927_in,                      
			input    [width-1:0]    x928_in,                      
			input    [width-1:0]    x929_in,                      
			input    [width-1:0]    x930_in,                      
			input    [width-1:0]    x931_in,                      
			input    [width-1:0]    x932_in,                      
			input    [width-1:0]    x933_in,                      
			input    [width-1:0]    x934_in,                      
			input    [width-1:0]    x935_in,                      
			input    [width-1:0]    x936_in,                      
			input    [width-1:0]    x937_in,                      
			input    [width-1:0]    x938_in,                      
			input    [width-1:0]    x939_in,                      
			input    [width-1:0]    x940_in,                      
			input    [width-1:0]    x941_in,                      
			input    [width-1:0]    x942_in,                      
			input    [width-1:0]    x943_in,                      
			input    [width-1:0]    x944_in,                      
			input    [width-1:0]    x945_in,                      
			input    [width-1:0]    x946_in,                      
			input    [width-1:0]    x947_in,                      
			input    [width-1:0]    x948_in,                      
			input    [width-1:0]    x949_in,                      
			input    [width-1:0]    x950_in,                      
			input    [width-1:0]    x951_in,                      
			input    [width-1:0]    x952_in,                      
			input    [width-1:0]    x953_in,                      
			input    [width-1:0]    x954_in,                      
			input    [width-1:0]    x955_in,                      
			input    [width-1:0]    x956_in,                      
			input    [width-1:0]    x957_in,                      
			input    [width-1:0]    x958_in,                      
			input    [width-1:0]    x959_in,                      
			input    [width-1:0]    x960_in,                      
			input    [width-1:0]    x961_in,                      
			input    [width-1:0]    x962_in,                      
			input    [width-1:0]    x963_in,                      
			input    [width-1:0]    x964_in,                      
			input    [width-1:0]    x965_in,                      
			input    [width-1:0]    x966_in,                      
			input    [width-1:0]    x967_in,                      
			input    [width-1:0]    x968_in,                      
			input    [width-1:0]    x969_in,                      
			input    [width-1:0]    x970_in,                      
			input    [width-1:0]    x971_in,                      
			input    [width-1:0]    x972_in,                      
			input    [width-1:0]    x973_in,                      
			input    [width-1:0]    x974_in,                      
			input    [width-1:0]    x975_in,                      
			input    [width-1:0]    x976_in,                      
			input    [width-1:0]    x977_in,                      
			input    [width-1:0]    x978_in,                      
			input    [width-1:0]    x979_in,                      
			input    [width-1:0]    x980_in,                      
			input    [width-1:0]    x981_in,                      
			input    [width-1:0]    x982_in,                      
			input    [width-1:0]    x983_in,                      
			input    [width-1:0]    x984_in,                      
			input    [width-1:0]    x985_in,                      
			input    [width-1:0]    x986_in,                      
			input    [width-1:0]    x987_in,                      
			input    [width-1:0]    x988_in,                      
			input    [width-1:0]    x989_in,                      
			input    [width-1:0]    x990_in,                      
			input    [width-1:0]    x991_in,                      
			input    [width-1:0]    x992_in,                      
			input    [width-1:0]    x993_in,                      
			input    [width-1:0]    x994_in,                      
			input    [width-1:0]    x995_in,                      
			input    [width-1:0]    x996_in,                      
			input    [width-1:0]    x997_in,                      
			input    [width-1:0]    x998_in,                      
			input    [width-1:0]    x999_in,                      
			input    [width-1:0]    x1000_in,                     
			input    [width-1:0]    x1001_in,                     
			input    [width-1:0]    x1002_in,                     
			input    [width-1:0]    x1003_in,                     
			input    [width-1:0]    x1004_in,                     
			input    [width-1:0]    x1005_in,                     
			input    [width-1:0]    x1006_in,                     
			input    [width-1:0]    x1007_in,                     
			input    [width-1:0]    x1008_in,                     
			input    [width-1:0]    x1009_in,                     
			input    [width-1:0]    x1010_in,                     
			input    [width-1:0]    x1011_in,                     
			input    [width-1:0]    x1012_in,                     
			input    [width-1:0]    x1013_in,                     
			input    [width-1:0]    x1014_in,                     
			input    [width-1:0]    x1015_in,                     
			input    [width-1:0]    x1016_in,                     
			input    [width-1:0]    x1017_in,                     
			input    [width-1:0]    x1018_in,                     
			input    [width-1:0]    x1019_in,                     
			input    [width-1:0]    x1020_in,                     
			input    [width-1:0]    x1021_in,                     
			input    [width-1:0]    x1022_in,                     
			input    [width-1:0]    x1023_in,                     
			input    [width-1:0]    x1024_in,                     
			input    [width-1:0]    x1025_in,                     
			input    [width-1:0]    x1026_in,                     
			input    [width-1:0]    x1027_in,                     
			input    [width-1:0]    x1028_in,                     
			input    [width-1:0]    x1029_in,                     
			input    [width-1:0]    x1030_in,                     
			input    [width-1:0]    x1031_in,                     
			input    [width-1:0]    x1032_in,                     
			input    [width-1:0]    x1033_in,                     
			input    [width-1:0]    x1034_in,                     
			input    [width-1:0]    x1035_in,                     
			input    [width-1:0]    x1036_in,                     
			input    [width-1:0]    x1037_in,                     
			input    [width-1:0]    x1038_in,                     
			input    [width-1:0]    x1039_in,                     
			input    [width-1:0]    x1040_in,                     
			input    [width-1:0]    x1041_in,                     
			input    [width-1:0]    x1042_in,                     
			input    [width-1:0]    x1043_in,                     
			input    [width-1:0]    x1044_in,                     
			input    [width-1:0]    x1045_in,                     
			input    [width-1:0]    x1046_in,                     
			input    [width-1:0]    x1047_in,                     
			input    [width-1:0]    x1048_in,                     
			input    [width-1:0]    x1049_in,                     
			input    [width-1:0]    x1050_in,                     
			input    [width-1:0]    x1051_in,                     
			input    [width-1:0]    x1052_in,                     
			input    [width-1:0]    x1053_in,                     
			input    [width-1:0]    x1054_in,                     
			input    [width-1:0]    x1055_in,                     
			input    [width-1:0]    x1056_in,                     
			input    [width-1:0]    x1057_in,                     
			input    [width-1:0]    x1058_in,                     
			input    [width-1:0]    x1059_in,                     
			input    [width-1:0]    x1060_in,                     
			input    [width-1:0]    x1061_in,                     
			input    [width-1:0]    x1062_in,                     
			input    [width-1:0]    x1063_in,                     
			input    [width-1:0]    x1064_in,                     
			input    [width-1:0]    x1065_in,                     
			input    [width-1:0]    x1066_in,                     
			input    [width-1:0]    x1067_in,                     
			input    [width-1:0]    x1068_in,                     
			input    [width-1:0]    x1069_in,                     
			input    [width-1:0]    x1070_in,                     
			input    [width-1:0]    x1071_in,                     
			input    [width-1:0]    x1072_in,                     
			input    [width-1:0]    x1073_in,                     
			input    [width-1:0]    x1074_in,                     
			input    [width-1:0]    x1075_in,                     
			input    [width-1:0]    x1076_in,                     
			input    [width-1:0]    x1077_in,                     
			input    [width-1:0]    x1078_in,                     
			input    [width-1:0]    x1079_in,                     
			input    [width-1:0]    x1080_in,                     
			input    [width-1:0]    x1081_in,                     
			input    [width-1:0]    x1082_in,                     
			input    [width-1:0]    x1083_in,                     
			input    [width-1:0]    x1084_in,                     
			input    [width-1:0]    x1085_in,                     
			input    [width-1:0]    x1086_in,                     
			input    [width-1:0]    x1087_in,                     
			input    [width-1:0]    x1088_in,                     
			input    [width-1:0]    x1089_in,                     
			input    [width-1:0]    x1090_in,                     
			input    [width-1:0]    x1091_in,                     
			input    [width-1:0]    x1092_in,                     
			input    [width-1:0]    x1093_in,                     
			input    [width-1:0]    x1094_in,                     
			input    [width-1:0]    x1095_in,                     
			input    [width-1:0]    x1096_in,                     
			input    [width-1:0]    x1097_in,                     
			input    [width-1:0]    x1098_in,                     
			input    [width-1:0]    x1099_in,                     
			input    [width-1:0]    x1100_in,                     
			input    [width-1:0]    x1101_in,                     
			input    [width-1:0]    x1102_in,                     
			input    [width-1:0]    x1103_in,                     
			input    [width-1:0]    x1104_in,                     
			input    [width-1:0]    x1105_in,                     
			input    [width-1:0]    x1106_in,                     
			input    [width-1:0]    x1107_in,                     
			input    [width-1:0]    x1108_in,                     
			input    [width-1:0]    x1109_in,                     
			input    [width-1:0]    x1110_in,                     
			input    [width-1:0]    x1111_in,                     
			input    [width-1:0]    x1112_in,                     
			input    [width-1:0]    x1113_in,                     
			input    [width-1:0]    x1114_in,                     
			input    [width-1:0]    x1115_in,                     
			input    [width-1:0]    x1116_in,                     
			input    [width-1:0]    x1117_in,                     
			input    [width-1:0]    x1118_in,                     
			input    [width-1:0]    x1119_in,                     
			input    [width-1:0]    x1120_in,                     
			input    [width-1:0]    x1121_in,                     
			input    [width-1:0]    x1122_in,                     
			input    [width-1:0]    x1123_in,                     
			input    [width-1:0]    x1124_in,                     
			input    [width-1:0]    x1125_in,                     
			input    [width-1:0]    x1126_in,                     
			input    [width-1:0]    x1127_in,                     
			input    [width-1:0]    x1128_in,                     
			input    [width-1:0]    x1129_in,                     
			input    [width-1:0]    x1130_in,                     
			input    [width-1:0]    x1131_in,                     
			input    [width-1:0]    x1132_in,                     
			input    [width-1:0]    x1133_in,                     
			input    [width-1:0]    x1134_in,                     
			input    [width-1:0]    x1135_in,                     
			input    [width-1:0]    x1136_in,                     
			input    [width-1:0]    x1137_in,                     
			input    [width-1:0]    x1138_in,                     
			input    [width-1:0]    x1139_in,                     
			input    [width-1:0]    x1140_in,                     
			input    [width-1:0]    x1141_in,                     
			input    [width-1:0]    x1142_in,                     
			input    [width-1:0]    x1143_in,                     
			input    [width-1:0]    x1144_in,                     
			input    [width-1:0]    x1145_in,                     
			input    [width-1:0]    x1146_in,                     
			input    [width-1:0]    x1147_in,                     
			input    [width-1:0]    x1148_in,                     
			input    [width-1:0]    x1149_in,                     
			input    [width-1:0]    x1150_in,                     
			input    [width-1:0]    x1151_in,                     
			input    [width-1:0]    x1152_in,                     
			input    [width-1:0]    x1153_in,                     
			input    [width-1:0]    x1154_in,                     
			input    [width-1:0]    x1155_in,                     
			input    [width-1:0]    x1156_in,                     
			input    [width-1:0]    x1157_in,                     
			input    [width-1:0]    x1158_in,                     
			input    [width-1:0]    x1159_in,                     
			input    [width-1:0]    x1160_in,                     
			input    [width-1:0]    x1161_in,                     
			input    [width-1:0]    x1162_in,                     
			input    [width-1:0]    x1163_in,                     
			input    [width-1:0]    x1164_in,                     
			input    [width-1:0]    x1165_in,                     
			input    [width-1:0]    x1166_in,                     
			input    [width-1:0]    x1167_in,                     
			input    [width-1:0]    x1168_in,                     
			input    [width-1:0]    x1169_in,                     
			input    [width-1:0]    x1170_in,                     
			input    [width-1:0]    x1171_in,                     
			input    [width-1:0]    x1172_in,                     
			input    [width-1:0]    x1173_in,                     
			input    [width-1:0]    x1174_in,                     
			input    [width-1:0]    x1175_in,                     
			input    [width-1:0]    x1176_in,                     
			input    [width-1:0]    x1177_in,                     
			input    [width-1:0]    x1178_in,                     
			input    [width-1:0]    x1179_in,                     
			input    [width-1:0]    x1180_in,                     
			input    [width-1:0]    x1181_in,                     
			input    [width-1:0]    x1182_in,                     
			input    [width-1:0]    x1183_in,                     
			input    [width-1:0]    x1184_in,                     
			input    [width-1:0]    x1185_in,                     
			input    [width-1:0]    x1186_in,                     
			input    [width-1:0]    x1187_in,                     
			input    [width-1:0]    x1188_in,                     
			input    [width-1:0]    x1189_in,                     
			input    [width-1:0]    x1190_in,                     
			input    [width-1:0]    x1191_in,                     
			input    [width-1:0]    x1192_in,                     
			input    [width-1:0]    x1193_in,                     
			input    [width-1:0]    x1194_in,                     
			input    [width-1:0]    x1195_in,                     
			input    [width-1:0]    x1196_in,                     
			input    [width-1:0]    x1197_in,                     
			input    [width-1:0]    x1198_in,                     
			input    [width-1:0]    x1199_in,                     
			input    [width-1:0]    x1200_in,                     
			input    [width-1:0]    x1201_in,                     
			input    [width-1:0]    x1202_in,                     
			input    [width-1:0]    x1203_in,                     
			input    [width-1:0]    x1204_in,                     
			input    [width-1:0]    x1205_in,                     
			input    [width-1:0]    x1206_in,                     
			input    [width-1:0]    x1207_in,                     
			input    [width-1:0]    x1208_in,                     
			input    [width-1:0]    x1209_in,                     
			input    [width-1:0]    x1210_in,                     
			input    [width-1:0]    x1211_in,                     
			input    [width-1:0]    x1212_in,                     
			input    [width-1:0]    x1213_in,                     
			input    [width-1:0]    x1214_in,                     
			input    [width-1:0]    x1215_in,                     
			input    [width-1:0]    x1216_in,                     
			input    [width-1:0]    x1217_in,                     
			input    [width-1:0]    x1218_in,                     
			input    [width-1:0]    x1219_in,                     
			input    [width-1:0]    x1220_in,                     
			input    [width-1:0]    x1221_in,                     
			input    [width-1:0]    x1222_in,                     
			input    [width-1:0]    x1223_in,                     
			input    [width-1:0]    x1224_in,                     
			input    [width-1:0]    x1225_in,                     
			input    [width-1:0]    x1226_in,                     
			input    [width-1:0]    x1227_in,                     
			input    [width-1:0]    x1228_in,                     
			input    [width-1:0]    x1229_in,                     
			input    [width-1:0]    x1230_in,                     
			input    [width-1:0]    x1231_in,                     
			input    [width-1:0]    x1232_in,                     
			input    [width-1:0]    x1233_in,                     
			input    [width-1:0]    x1234_in,                     
			input    [width-1:0]    x1235_in,                     
			input    [width-1:0]    x1236_in,                     
			input    [width-1:0]    x1237_in,                     
			input    [width-1:0]    x1238_in,                     
			input    [width-1:0]    x1239_in,                     
			input    [width-1:0]    x1240_in,                     
			input    [width-1:0]    x1241_in,                     
			input    [width-1:0]    x1242_in,                     
			input    [width-1:0]    x1243_in,                     
			input    [width-1:0]    x1244_in,                     
			input    [width-1:0]    x1245_in,                     
			input    [width-1:0]    x1246_in,                     
			input    [width-1:0]    x1247_in,                     
			input    [width-1:0]    x1248_in,                     
			input    [width-1:0]    x1249_in,                     
			input    [width-1:0]    x1250_in,                     
			input    [width-1:0]    x1251_in,                     
			input    [width-1:0]    x1252_in,                     
			input    [width-1:0]    x1253_in,                     
			input    [width-1:0]    x1254_in,                     
			input    [width-1:0]    x1255_in,                     
			input    [width-1:0]    x1256_in,                     
			input    [width-1:0]    x1257_in,                     
			input    [width-1:0]    x1258_in,                     
			input    [width-1:0]    x1259_in,                     
			input    [width-1:0]    x1260_in,                     
			input    [width-1:0]    x1261_in,                     
			input    [width-1:0]    x1262_in,                     
			input    [width-1:0]    x1263_in,                     
			input    [width-1:0]    x1264_in,                     
			input    [width-1:0]    x1265_in,                     
			input    [width-1:0]    x1266_in,                     
			input    [width-1:0]    x1267_in,                     
			input    [width-1:0]    x1268_in,                     
			input    [width-1:0]    x1269_in,                     
			input    [width-1:0]    x1270_in,                     
			input    [width-1:0]    x1271_in,                     
			input    [width-1:0]    x1272_in,                     
			input    [width-1:0]    x1273_in,                     
			input    [width-1:0]    x1274_in,                     
			input    [width-1:0]    x1275_in,                     
			input    [width-1:0]    x1276_in,                     
			input    [width-1:0]    x1277_in,                     
			input    [width-1:0]    x1278_in,                     
			input    [width-1:0]    x1279_in,                     
			input    [width-1:0]    x1280_in,                     
			input    [width-1:0]    x1281_in,                     
			input    [width-1:0]    x1282_in,                     
			input    [width-1:0]    x1283_in,                     
			input    [width-1:0]    x1284_in,                     
			input    [width-1:0]    x1285_in,                     
			input    [width-1:0]    x1286_in,                     
			input    [width-1:0]    x1287_in,                     
			input    [width-1:0]    x1288_in,                     
			input    [width-1:0]    x1289_in,                     
			input    [width-1:0]    x1290_in,                     
			input    [width-1:0]    x1291_in,                     
			input    [width-1:0]    x1292_in,                     
			input    [width-1:0]    x1293_in,                     
			input    [width-1:0]    x1294_in,                     
			input    [width-1:0]    x1295_in,                     
			input    [width-1:0]    x1296_in,                     
			input    [width-1:0]    x1297_in,                     
			input    [width-1:0]    x1298_in,                     
			input    [width-1:0]    x1299_in,                     
			input    [width-1:0]    x1300_in,                     
			input    [width-1:0]    x1301_in,                     
			input    [width-1:0]    x1302_in,                     
			input    [width-1:0]    x1303_in,                     
			input    [width-1:0]    x1304_in,                     
			input    [width-1:0]    x1305_in,                     
			input    [width-1:0]    x1306_in,                     
			input    [width-1:0]    x1307_in,                     
			input    [width-1:0]    x1308_in,                     
			input    [width-1:0]    x1309_in,                     
			input    [width-1:0]    x1310_in,                     
			input    [width-1:0]    x1311_in,                     
			input    [width-1:0]    x1312_in,                     
			input    [width-1:0]    x1313_in,                     
			input    [width-1:0]    x1314_in,                     
			input    [width-1:0]    x1315_in,                     
			input    [width-1:0]    x1316_in,                     
			input    [width-1:0]    x1317_in,                     
			input    [width-1:0]    x1318_in,                     
			input    [width-1:0]    x1319_in,                     
			input    [width-1:0]    x1320_in,                     
			input    [width-1:0]    x1321_in,                     
			input    [width-1:0]    x1322_in,                     
			input    [width-1:0]    x1323_in,                     
			input    [width-1:0]    x1324_in,                     
			input    [width-1:0]    x1325_in,                     
			input    [width-1:0]    x1326_in,                     
			input    [width-1:0]    x1327_in,                     
			input    [width-1:0]    x1328_in,                     
			input    [width-1:0]    x1329_in,                     
			input    [width-1:0]    x1330_in,                     
			input    [width-1:0]    x1331_in,                     
			input    [width-1:0]    x1332_in,                     
			input    [width-1:0]    x1333_in,                     
			input    [width-1:0]    x1334_in,                     
			input    [width-1:0]    x1335_in,                     
			input    [width-1:0]    x1336_in,                     
			input    [width-1:0]    x1337_in,                     
			input    [width-1:0]    x1338_in,                     
			input    [width-1:0]    x1339_in,                     
			input    [width-1:0]    x1340_in,                     
			input    [width-1:0]    x1341_in,                     
			input    [width-1:0]    x1342_in,                     
			input    [width-1:0]    x1343_in,                     
			input    [width-1:0]    x1344_in,                     
			input    [width-1:0]    x1345_in,                     
			input    [width-1:0]    x1346_in,                     
			input    [width-1:0]    x1347_in,                     
			input    [width-1:0]    x1348_in,                     
			input    [width-1:0]    x1349_in,                     
			input    [width-1:0]    x1350_in,                     
			input    [width-1:0]    x1351_in,                     
			input    [width-1:0]    x1352_in,                     
			input    [width-1:0]    x1353_in,                     
			input    [width-1:0]    x1354_in,                     
			input    [width-1:0]    x1355_in,                     
			input    [width-1:0]    x1356_in,                     
			input    [width-1:0]    x1357_in,                     
			input    [width-1:0]    x1358_in,                     
			input    [width-1:0]    x1359_in,                     
			input    [width-1:0]    x1360_in,                     
			input    [width-1:0]    x1361_in,                     
			input    [width-1:0]    x1362_in,                     
			input    [width-1:0]    x1363_in,                     
			input    [width-1:0]    x1364_in,                     
			input    [width-1:0]    x1365_in,                     
			input    [width-1:0]    x1366_in,                     
			input    [width-1:0]    x1367_in,                     
			input    [width-1:0]    x1368_in,                     
			input    [width-1:0]    x1369_in,                     
			input    [width-1:0]    x1370_in,                     
			input    [width-1:0]    x1371_in,                     
			input    [width-1:0]    x1372_in,                     
			input    [width-1:0]    x1373_in,                     
			input    [width-1:0]    x1374_in,                     
			input    [width-1:0]    x1375_in,                     
			input    [width-1:0]    x1376_in,                     
			input    [width-1:0]    x1377_in,                     
			input    [width-1:0]    x1378_in,                     
			input    [width-1:0]    x1379_in,                     
			input    [width-1:0]    x1380_in,                     
			input    [width-1:0]    x1381_in,                     
			input    [width-1:0]    x1382_in,                     
			input    [width-1:0]    x1383_in,                     
			input    [width-1:0]    x1384_in,                     
			input    [width-1:0]    x1385_in,                     
			input    [width-1:0]    x1386_in,                     
			input    [width-1:0]    x1387_in,                     
			input    [width-1:0]    x1388_in,                     
			input    [width-1:0]    x1389_in,                     
			input    [width-1:0]    x1390_in,                     
			input    [width-1:0]    x1391_in,                     
			input    [width-1:0]    x1392_in,                     
			input    [width-1:0]    x1393_in,                     
			input    [width-1:0]    x1394_in,                     
			input    [width-1:0]    x1395_in,                     
			input    [width-1:0]    x1396_in,                     
			input    [width-1:0]    x1397_in,                     
			input    [width-1:0]    x1398_in,                     
			input    [width-1:0]    x1399_in,                     
			input    [width-1:0]    x1400_in,                     
			input    [width-1:0]    x1401_in,                     
			input    [width-1:0]    x1402_in,                     
			input    [width-1:0]    x1403_in,                     
			input    [width-1:0]    x1404_in,                     
			input    [width-1:0]    x1405_in,                     
			input    [width-1:0]    x1406_in,                     
			input    [width-1:0]    x1407_in,                     
			input    [width-1:0]    x1408_in,                     
			input    [width-1:0]    x1409_in,                     
			input    [width-1:0]    x1410_in,                     
			input    [width-1:0]    x1411_in,                     
			input    [width-1:0]    x1412_in,                     
			input    [width-1:0]    x1413_in,                     
			input    [width-1:0]    x1414_in,                     
			input    [width-1:0]    x1415_in,                     
			input    [width-1:0]    x1416_in,                     
			input    [width-1:0]    x1417_in,                     
			input    [width-1:0]    x1418_in,                     
			input    [width-1:0]    x1419_in,                     
			input    [width-1:0]    x1420_in,                     
			input    [width-1:0]    x1421_in,                     
			input    [width-1:0]    x1422_in,                     
			input    [width-1:0]    x1423_in,                     
			input    [width-1:0]    x1424_in,                     
			input    [width-1:0]    x1425_in,                     
			input    [width-1:0]    x1426_in,                     
			input    [width-1:0]    x1427_in,                     
			input    [width-1:0]    x1428_in,                     
			input    [width-1:0]    x1429_in,                     
			input    [width-1:0]    x1430_in,                     
			input    [width-1:0]    x1431_in,                     
			input    [width-1:0]    x1432_in,                     
			input    [width-1:0]    x1433_in,                     
			input    [width-1:0]    x1434_in,                     
			input    [width-1:0]    x1435_in,                     
			input    [width-1:0]    x1436_in,                     
			input    [width-1:0]    x1437_in,                     
			input    [width-1:0]    x1438_in,                     
			input    [width-1:0]    x1439_in,                     
			input    [width-1:0]    x1440_in,                     
			input    [width-1:0]    x1441_in,                     
			input    [width-1:0]    x1442_in,                     
			input    [width-1:0]    x1443_in,                     
			input    [width-1:0]    x1444_in,                     
			input    [width-1:0]    x1445_in,                     
			input    [width-1:0]    x1446_in,                     
			input    [width-1:0]    x1447_in,                     
			input    [width-1:0]    x1448_in,                     
			input    [width-1:0]    x1449_in,                     
			input    [width-1:0]    x1450_in,                     
			input    [width-1:0]    x1451_in,                     
			input    [width-1:0]    x1452_in,                     
			input    [width-1:0]    x1453_in,                     
			input    [width-1:0]    x1454_in,                     
			input    [width-1:0]    x1455_in,                     
			input    [width-1:0]    x1456_in,                     
			input    [width-1:0]    x1457_in,                     
			input    [width-1:0]    x1458_in,                     
			input    [width-1:0]    x1459_in,                     
			input    [width-1:0]    x1460_in,                     
			input    [width-1:0]    x1461_in,                     
			input    [width-1:0]    x1462_in,                     
			input    [width-1:0]    x1463_in,                     
			input    [width-1:0]    x1464_in,                     
			input    [width-1:0]    x1465_in,                     
			input    [width-1:0]    x1466_in,                     
			input    [width-1:0]    x1467_in,                     
			input    [width-1:0]    x1468_in,                     
			input    [width-1:0]    x1469_in,                     
			input    [width-1:0]    x1470_in,                     
			input    [width-1:0]    x1471_in,                     
			input    [width-1:0]    x1472_in,                     
			input    [width-1:0]    x1473_in,                     
			input    [width-1:0]    x1474_in,                     
			input    [width-1:0]    x1475_in,                     
			input    [width-1:0]    x1476_in,                     
			input    [width-1:0]    x1477_in,                     
			input    [width-1:0]    x1478_in,                     
			input    [width-1:0]    x1479_in,                     
			input    [width-1:0]    x1480_in,                     
			input    [width-1:0]    x1481_in,                     
			input    [width-1:0]    x1482_in,                     
			input    [width-1:0]    x1483_in,                     
			input    [width-1:0]    x1484_in,                     
			input    [width-1:0]    x1485_in,                     
			input    [width-1:0]    x1486_in,                     
			input    [width-1:0]    x1487_in,                     
			input    [width-1:0]    x1488_in,                     
			input    [width-1:0]    x1489_in,                     
			input    [width-1:0]    x1490_in,                     
			input    [width-1:0]    x1491_in,                     
			input    [width-1:0]    x1492_in,                     
			input    [width-1:0]    x1493_in,                     
			input    [width-1:0]    x1494_in,                     
			input    [width-1:0]    x1495_in,                     
			input    [width-1:0]    x1496_in,                     
			input    [width-1:0]    x1497_in,                     
			input    [width-1:0]    x1498_in,                     
			input    [width-1:0]    x1499_in,                     
			input    [width-1:0]    x1500_in,                     
			input    [width-1:0]    x1501_in,                     
			input    [width-1:0]    x1502_in,                     
			input    [width-1:0]    x1503_in,                     
			input    [width-1:0]    x1504_in,                     
			input    [width-1:0]    x1505_in,                     
			input    [width-1:0]    x1506_in,                     
			input    [width-1:0]    x1507_in,                     
			input    [width-1:0]    x1508_in,                     
			input    [width-1:0]    x1509_in,                     
			input    [width-1:0]    x1510_in,                     
			input    [width-1:0]    x1511_in,                     
			input    [width-1:0]    x1512_in,                     
			input    [width-1:0]    x1513_in,                     
			input    [width-1:0]    x1514_in,                     
			input    [width-1:0]    x1515_in,                     
			input    [width-1:0]    x1516_in,                     
			input    [width-1:0]    x1517_in,                     
			input    [width-1:0]    x1518_in,                     
			input    [width-1:0]    x1519_in,                     
			input    [width-1:0]    x1520_in,                     
			input    [width-1:0]    x1521_in,                     
			input    [width-1:0]    x1522_in,                     
			input    [width-1:0]    x1523_in,                     
			input    [width-1:0]    x1524_in,                     
			input    [width-1:0]    x1525_in,                     
			input    [width-1:0]    x1526_in,                     
			input    [width-1:0]    x1527_in,                     
			input    [width-1:0]    x1528_in,                     
			input    [width-1:0]    x1529_in,                     
			input    [width-1:0]    x1530_in,                     
			input    [width-1:0]    x1531_in,                     
			input    [width-1:0]    x1532_in,                     
			input    [width-1:0]    x1533_in,                     
			input    [width-1:0]    x1534_in,                     
			input    [width-1:0]    x1535_in,                     
			input    [width-1:0]    x1536_in,                     
			input    [width-1:0]    x1537_in,                     
			input    [width-1:0]    x1538_in,                     
			input    [width-1:0]    x1539_in,                     
			input    [width-1:0]    x1540_in,                     
			input    [width-1:0]    x1541_in,                     
			input    [width-1:0]    x1542_in,                     
			input    [width-1:0]    x1543_in,                     
			input    [width-1:0]    x1544_in,                     
			input    [width-1:0]    x1545_in,                     
			input    [width-1:0]    x1546_in,                     
			input    [width-1:0]    x1547_in,                     
			input    [width-1:0]    x1548_in,                     
			input    [width-1:0]    x1549_in,                     
			input    [width-1:0]    x1550_in,                     
			input    [width-1:0]    x1551_in,                     
			input    [width-1:0]    x1552_in,                     
			input    [width-1:0]    x1553_in,                     
			input    [width-1:0]    x1554_in,                     
			input    [width-1:0]    x1555_in,                     
			input    [width-1:0]    x1556_in,                     
			input    [width-1:0]    x1557_in,                     
			input    [width-1:0]    x1558_in,                     
			input    [width-1:0]    x1559_in,                     
			input    [width-1:0]    x1560_in,                     
			input    [width-1:0]    x1561_in,                     
			input    [width-1:0]    x1562_in,                     
			input    [width-1:0]    x1563_in,                     
			input    [width-1:0]    x1564_in,                     
			input    [width-1:0]    x1565_in,                     
			input    [width-1:0]    x1566_in,                     
			input    [width-1:0]    x1567_in,                     
			input    [width-1:0]    x1568_in,                     
			input    [width-1:0]    x1569_in,                     
			input    [width-1:0]    x1570_in,                     
			input    [width-1:0]    x1571_in,                     
			input    [width-1:0]    x1572_in,                     
			input    [width-1:0]    x1573_in,                     
			input    [width-1:0]    x1574_in,                     
			input    [width-1:0]    x1575_in,                     
			input    [width-1:0]    x1576_in,                     
			input    [width-1:0]    x1577_in,                     
			input    [width-1:0]    x1578_in,                     
			input    [width-1:0]    x1579_in,                     
			input    [width-1:0]    x1580_in,                     
			input    [width-1:0]    x1581_in,                     
			input    [width-1:0]    x1582_in,                     
			input    [width-1:0]    x1583_in,                     
			input    [width-1:0]    x1584_in,                     
			input    [width-1:0]    x1585_in,                     
			input    [width-1:0]    x1586_in,                     
			input    [width-1:0]    x1587_in,                     
			input    [width-1:0]    x1588_in,                     
			input    [width-1:0]    x1589_in,                     
			input    [width-1:0]    x1590_in,                     
			input    [width-1:0]    x1591_in,                     
			input    [width-1:0]    x1592_in,                     
			input    [width-1:0]    x1593_in,                     
			input    [width-1:0]    x1594_in,                     
			input    [width-1:0]    x1595_in,                     
			input    [width-1:0]    x1596_in,                     
			input    [width-1:0]    x1597_in,                     
			input    [width-1:0]    x1598_in,                     
			input    [width-1:0]    x1599_in,                     
			input    [width-1:0]    x1600_in,                     
			input    [width-1:0]    x1601_in,                     
			input    [width-1:0]    x1602_in,                     
			input    [width-1:0]    x1603_in,                     
			input    [width-1:0]    x1604_in,                     
			input    [width-1:0]    x1605_in,                     
			input    [width-1:0]    x1606_in,                     
			input    [width-1:0]    x1607_in,                     
			input    [width-1:0]    x1608_in,                     
			input    [width-1:0]    x1609_in,                     
			input    [width-1:0]    x1610_in,                     
			input    [width-1:0]    x1611_in,                     
			input    [width-1:0]    x1612_in,                     
			input    [width-1:0]    x1613_in,                     
			input    [width-1:0]    x1614_in,                     
			input    [width-1:0]    x1615_in,                     
			input    [width-1:0]    x1616_in,                     
			input    [width-1:0]    x1617_in,                     
			input    [width-1:0]    x1618_in,                     
			input    [width-1:0]    x1619_in,                     
			input    [width-1:0]    x1620_in,                     
			input    [width-1:0]    x1621_in,                     
			input    [width-1:0]    x1622_in,                     
			input    [width-1:0]    x1623_in,                     
			input    [width-1:0]    x1624_in,                     
			input    [width-1:0]    x1625_in,                     
			input    [width-1:0]    x1626_in,                     
			input    [width-1:0]    x1627_in,                     
			input    [width-1:0]    x1628_in,                     
			input    [width-1:0]    x1629_in,                     
			input    [width-1:0]    x1630_in,                     
			input    [width-1:0]    x1631_in,                     
			input    [width-1:0]    x1632_in,                     
			input    [width-1:0]    x1633_in,                     
			input    [width-1:0]    x1634_in,                     
			input    [width-1:0]    x1635_in,                     
			input    [width-1:0]    x1636_in,                     
			input    [width-1:0]    x1637_in,                     
			input    [width-1:0]    x1638_in,                     
			input    [width-1:0]    x1639_in,                     
			input    [width-1:0]    x1640_in,                     
			input    [width-1:0]    x1641_in,                     
			input    [width-1:0]    x1642_in,                     
			input    [width-1:0]    x1643_in,                     
			input    [width-1:0]    x1644_in,                     
			input    [width-1:0]    x1645_in,                     
			input    [width-1:0]    x1646_in,                     
			input    [width-1:0]    x1647_in,                     
			input    [width-1:0]    x1648_in,                     
			input    [width-1:0]    x1649_in,                     
			input    [width-1:0]    x1650_in,                     
			input    [width-1:0]    x1651_in,                     
			input    [width-1:0]    x1652_in,                     
			input    [width-1:0]    x1653_in,                     
			input    [width-1:0]    x1654_in,                     
			input    [width-1:0]    x1655_in,                     
			input    [width-1:0]    x1656_in,                     
			input    [width-1:0]    x1657_in,                     
			input    [width-1:0]    x1658_in,                     
			input    [width-1:0]    x1659_in,                     
			input    [width-1:0]    x1660_in,                     
			input    [width-1:0]    x1661_in,                     
			input    [width-1:0]    x1662_in,                     
			input    [width-1:0]    x1663_in,                     
			input    [width-1:0]    x1664_in,                     
			input    [width-1:0]    x1665_in,                     
			input    [width-1:0]    x1666_in,                     
			input    [width-1:0]    x1667_in,                     
			input    [width-1:0]    x1668_in,                     
			input    [width-1:0]    x1669_in,                     
			input    [width-1:0]    x1670_in,                     
			input    [width-1:0]    x1671_in,                     
			input    [width-1:0]    x1672_in,                     
			input    [width-1:0]    x1673_in,                     
			input    [width-1:0]    x1674_in,                     
			input    [width-1:0]    x1675_in,                     
			input    [width-1:0]    x1676_in,                     
			input    [width-1:0]    x1677_in,                     
			input    [width-1:0]    x1678_in,                     
			input    [width-1:0]    x1679_in,                     
			input    [width-1:0]    x1680_in,                     
			input    [width-1:0]    x1681_in,                     
			input    [width-1:0]    x1682_in,                     
			input    [width-1:0]    x1683_in,                     
			input    [width-1:0]    x1684_in,                     
			input    [width-1:0]    x1685_in,                     
			input    [width-1:0]    x1686_in,                     
			input    [width-1:0]    x1687_in,                     
			input    [width-1:0]    x1688_in,                     
			input    [width-1:0]    x1689_in,                     
			input    [width-1:0]    x1690_in,                     
			input    [width-1:0]    x1691_in,                     
			input    [width-1:0]    x1692_in,                     
			input    [width-1:0]    x1693_in,                     
			input    [width-1:0]    x1694_in,                     
			input    [width-1:0]    x1695_in,                     
			input    [width-1:0]    x1696_in,                     
			input    [width-1:0]    x1697_in,                     
			input    [width-1:0]    x1698_in,                     
			input    [width-1:0]    x1699_in,                     
			input    [width-1:0]    x1700_in,                     
			input    [width-1:0]    x1701_in,                     
			input    [width-1:0]    x1702_in,                     
			input    [width-1:0]    x1703_in,                     
			input    [width-1:0]    x1704_in,                     
			input    [width-1:0]    x1705_in,                     
			input    [width-1:0]    x1706_in,                     
			input    [width-1:0]    x1707_in,                     
			input    [width-1:0]    x1708_in,                     
			input    [width-1:0]    x1709_in,                     
			input    [width-1:0]    x1710_in,                     
			input    [width-1:0]    x1711_in,                     
			input    [width-1:0]    x1712_in,                     
			input    [width-1:0]    x1713_in,                     
			input    [width-1:0]    x1714_in,                     
			input    [width-1:0]    x1715_in,                     
			input    [width-1:0]    x1716_in,                     
			input    [width-1:0]    x1717_in,                     
			input    [width-1:0]    x1718_in,                     
			input    [width-1:0]    x1719_in,                     
			input    [width-1:0]    x1720_in,                     
			input    [width-1:0]    x1721_in,                     
			input    [width-1:0]    x1722_in,                     
			input    [width-1:0]    x1723_in,                     
			input    [width-1:0]    x1724_in,                     
			input    [width-1:0]    x1725_in,                     
			input    [width-1:0]    x1726_in,                     
			input    [width-1:0]    x1727_in,                     
			input    [width-1:0]    x1728_in,                     
			input    [width-1:0]    x1729_in,                     
			input    [width-1:0]    x1730_in,                     
			input    [width-1:0]    x1731_in,                     
			input    [width-1:0]    x1732_in,                     
			input    [width-1:0]    x1733_in,                     
			input    [width-1:0]    x1734_in,                     
			input    [width-1:0]    x1735_in,                     
			input    [width-1:0]    x1736_in,                     
			input    [width-1:0]    x1737_in,                     
			input    [width-1:0]    x1738_in,                     
			input    [width-1:0]    x1739_in,                     
			input    [width-1:0]    x1740_in,                     
			input    [width-1:0]    x1741_in,                     
			input    [width-1:0]    x1742_in,                     
			input    [width-1:0]    x1743_in,                     
			input    [width-1:0]    x1744_in,                     
			input    [width-1:0]    x1745_in,                     
			input    [width-1:0]    x1746_in,                     
			input    [width-1:0]    x1747_in,                     
			input    [width-1:0]    x1748_in,                     
			input    [width-1:0]    x1749_in,                     
			input    [width-1:0]    x1750_in,                     
			input    [width-1:0]    x1751_in,                     
			input    [width-1:0]    x1752_in,                     
			input    [width-1:0]    x1753_in,                     
			input    [width-1:0]    x1754_in,                     
			input    [width-1:0]    x1755_in,                     
			input    [width-1:0]    x1756_in,                     
			input    [width-1:0]    x1757_in,                     
			input    [width-1:0]    x1758_in,                     
			input    [width-1:0]    x1759_in,                     
			input    [width-1:0]    x1760_in,                     
			input    [width-1:0]    x1761_in,                     
			input    [width-1:0]    x1762_in,                     
			input    [width-1:0]    x1763_in,                     
			input    [width-1:0]    x1764_in,                     
			input    [width-1:0]    x1765_in,                     
			input    [width-1:0]    x1766_in,                     
			input    [width-1:0]    x1767_in,                     
			input    [width-1:0]    x1768_in,                     
			input    [width-1:0]    x1769_in,                     
			input    [width-1:0]    x1770_in,                     
			input    [width-1:0]    x1771_in,                     
			input    [width-1:0]    x1772_in,                     
			input    [width-1:0]    x1773_in,                     
			input    [width-1:0]    x1774_in,                     
			input    [width-1:0]    x1775_in,                     
			input    [width-1:0]    x1776_in,                     
			input    [width-1:0]    x1777_in,                     
			input    [width-1:0]    x1778_in,                     
			input    [width-1:0]    x1779_in,                     
			input    [width-1:0]    x1780_in,                     
			input    [width-1:0]    x1781_in,                     
			input    [width-1:0]    x1782_in,                     
			input    [width-1:0]    x1783_in,                     
			input    [width-1:0]    x1784_in,                     
			input    [width-1:0]    x1785_in,                     
			input    [width-1:0]    x1786_in,                     
			input    [width-1:0]    x1787_in,                     
			input    [width-1:0]    x1788_in,                     
			input    [width-1:0]    x1789_in,                     
			input    [width-1:0]    x1790_in,                     
			input    [width-1:0]    x1791_in,                     
			input    [width-1:0]    x1792_in,                     
			input    [width-1:0]    x1793_in,                     
			input    [width-1:0]    x1794_in,                     
			input    [width-1:0]    x1795_in,                     
			input    [width-1:0]    x1796_in,                     
			input    [width-1:0]    x1797_in,                     
			input    [width-1:0]    x1798_in,                     
			input    [width-1:0]    x1799_in,                     
			input    [width-1:0]    x1800_in,                     
			input    [width-1:0]    x1801_in,                     
			input    [width-1:0]    x1802_in,                     
			input    [width-1:0]    x1803_in,                     
			input    [width-1:0]    x1804_in,                     
			input    [width-1:0]    x1805_in,                     
			input    [width-1:0]    x1806_in,                     
			input    [width-1:0]    x1807_in,                     
			input    [width-1:0]    x1808_in,                     
			input    [width-1:0]    x1809_in,                     
			input    [width-1:0]    x1810_in,                     
			input    [width-1:0]    x1811_in,                     
			input    [width-1:0]    x1812_in,                     
			input    [width-1:0]    x1813_in,                     
			input    [width-1:0]    x1814_in,                     
			input    [width-1:0]    x1815_in,                     
			input    [width-1:0]    x1816_in,                     
			input    [width-1:0]    x1817_in,                     
			input    [width-1:0]    x1818_in,                     
			input    [width-1:0]    x1819_in,                     
			input    [width-1:0]    x1820_in,                     
			input    [width-1:0]    x1821_in,                     
			input    [width-1:0]    x1822_in,                     
			input    [width-1:0]    x1823_in,                     
			input    [width-1:0]    x1824_in,                     
			input    [width-1:0]    x1825_in,                     
			input    [width-1:0]    x1826_in,                     
			input    [width-1:0]    x1827_in,                     
			input    [width-1:0]    x1828_in,                     
			input    [width-1:0]    x1829_in,                     
			input    [width-1:0]    x1830_in,                     
			input    [width-1:0]    x1831_in,                     
			input    [width-1:0]    x1832_in,                     
			input    [width-1:0]    x1833_in,                     
			input    [width-1:0]    x1834_in,                     
			input    [width-1:0]    x1835_in,                     
			input    [width-1:0]    x1836_in,                     
			input    [width-1:0]    x1837_in,                     
			input    [width-1:0]    x1838_in,                     
			input    [width-1:0]    x1839_in,                     
			input    [width-1:0]    x1840_in,                     
			input    [width-1:0]    x1841_in,                     
			input    [width-1:0]    x1842_in,                     
			input    [width-1:0]    x1843_in,                     
			input    [width-1:0]    x1844_in,                     
			input    [width-1:0]    x1845_in,                     
			input    [width-1:0]    x1846_in,                     
			input    [width-1:0]    x1847_in,                     
			input    [width-1:0]    x1848_in,                     
			input    [width-1:0]    x1849_in,                     
			input    [width-1:0]    x1850_in,                     
			input    [width-1:0]    x1851_in,                     
			input    [width-1:0]    x1852_in,                     
			input    [width-1:0]    x1853_in,                     
			input    [width-1:0]    x1854_in,                     
			input    [width-1:0]    x1855_in,                     
			input    [width-1:0]    x1856_in,                     
			input    [width-1:0]    x1857_in,                     
			input    [width-1:0]    x1858_in,                     
			input    [width-1:0]    x1859_in,                     
			input    [width-1:0]    x1860_in,                     
			input    [width-1:0]    x1861_in,                     
			input    [width-1:0]    x1862_in,                     
			input    [width-1:0]    x1863_in,                     
			input    [width-1:0]    x1864_in,                     
			input    [width-1:0]    x1865_in,                     
			input    [width-1:0]    x1866_in,                     
			input    [width-1:0]    x1867_in,                     
			input    [width-1:0]    x1868_in,                     
			input    [width-1:0]    x1869_in,                     
			input    [width-1:0]    x1870_in,                     
			input    [width-1:0]    x1871_in,                     
			input    [width-1:0]    x1872_in,                     
			input    [width-1:0]    x1873_in,                     
			input    [width-1:0]    x1874_in,                     
			input    [width-1:0]    x1875_in,                     
			input    [width-1:0]    x1876_in,                     
			input    [width-1:0]    x1877_in,                     
			input    [width-1:0]    x1878_in,                     
			input    [width-1:0]    x1879_in,                     
			input    [width-1:0]    x1880_in,                     
			input    [width-1:0]    x1881_in,                     
			input    [width-1:0]    x1882_in,                     
			input    [width-1:0]    x1883_in,                     
			input    [width-1:0]    x1884_in,                     
			input    [width-1:0]    x1885_in,                     
			input    [width-1:0]    x1886_in,                     
			input    [width-1:0]    x1887_in,                     
			input    [width-1:0]    x1888_in,                     
			input    [width-1:0]    x1889_in,                     
			input    [width-1:0]    x1890_in,                     
			input    [width-1:0]    x1891_in,                     
			input    [width-1:0]    x1892_in,                     
			input    [width-1:0]    x1893_in,                     
			input    [width-1:0]    x1894_in,                     
			input    [width-1:0]    x1895_in,                     
			input    [width-1:0]    x1896_in,                     
			input    [width-1:0]    x1897_in,                     
			input    [width-1:0]    x1898_in,                     
			input    [width-1:0]    x1899_in,                     
			input    [width-1:0]    x1900_in,                     
			input    [width-1:0]    x1901_in,                     
			input    [width-1:0]    x1902_in,                     
			input    [width-1:0]    x1903_in,                     
			input    [width-1:0]    x1904_in,                     
			input    [width-1:0]    x1905_in,                     
			input    [width-1:0]    x1906_in,                     
			input    [width-1:0]    x1907_in,                     
			input    [width-1:0]    x1908_in,                     
			input    [width-1:0]    x1909_in,                     
			input    [width-1:0]    x1910_in,                     
			input    [width-1:0]    x1911_in,                     
			input    [width-1:0]    x1912_in,                     
			input    [width-1:0]    x1913_in,                     
			input    [width-1:0]    x1914_in,                     
			input    [width-1:0]    x1915_in,                     
			input    [width-1:0]    x1916_in,                     
			input    [width-1:0]    x1917_in,                     
			input    [width-1:0]    x1918_in,                     
			input    [width-1:0]    x1919_in,                     
			input    [width-1:0]    x1920_in,                     
			input    [width-1:0]    x1921_in,                     
			input    [width-1:0]    x1922_in,                     
			input    [width-1:0]    x1923_in,                     
			input    [width-1:0]    x1924_in,                     
			input    [width-1:0]    x1925_in,                     
			input    [width-1:0]    x1926_in,                     
			input    [width-1:0]    x1927_in,                     
			input    [width-1:0]    x1928_in,                     
			input    [width-1:0]    x1929_in,                     
			input    [width-1:0]    x1930_in,                     
			input    [width-1:0]    x1931_in,                     
			input    [width-1:0]    x1932_in,                     
			input    [width-1:0]    x1933_in,                     
			input    [width-1:0]    x1934_in,                     
			input    [width-1:0]    x1935_in,                     
			input    [width-1:0]    x1936_in,                     
			input    [width-1:0]    x1937_in,                     
			input    [width-1:0]    x1938_in,                     
			input    [width-1:0]    x1939_in,                     
			input    [width-1:0]    x1940_in,                     
			input    [width-1:0]    x1941_in,                     
			input    [width-1:0]    x1942_in,                     
			input    [width-1:0]    x1943_in,                     
			input    [width-1:0]    x1944_in,                     
			input    [width-1:0]    x1945_in,                     
			input    [width-1:0]    x1946_in,                     
			input    [width-1:0]    x1947_in,                     
			input    [width-1:0]    x1948_in,                     
			input    [width-1:0]    x1949_in,                     
			input    [width-1:0]    x1950_in,                     
			input    [width-1:0]    x1951_in,                     
			input    [width-1:0]    x1952_in,                     
			input    [width-1:0]    x1953_in,                     
			input    [width-1:0]    x1954_in,                     
			input    [width-1:0]    x1955_in,                     
			input    [width-1:0]    x1956_in,                     
			input    [width-1:0]    x1957_in,                     
			input    [width-1:0]    x1958_in,                     
			input    [width-1:0]    x1959_in,                     
			input    [width-1:0]    x1960_in,                     
			input    [width-1:0]    x1961_in,                     
			input    [width-1:0]    x1962_in,                     
			input    [width-1:0]    x1963_in,                     
			input    [width-1:0]    x1964_in,                     
			input    [width-1:0]    x1965_in,                     
			input    [width-1:0]    x1966_in,                     
			input    [width-1:0]    x1967_in,                     
			input    [width-1:0]    x1968_in,                     
			input    [width-1:0]    x1969_in,                     
			input    [width-1:0]    x1970_in,                     
			input    [width-1:0]    x1971_in,                     
			input    [width-1:0]    x1972_in,                     
			input    [width-1:0]    x1973_in,                     
			input    [width-1:0]    x1974_in,                     
			input    [width-1:0]    x1975_in,                     
			input    [width-1:0]    x1976_in,                     
			input    [width-1:0]    x1977_in,                     
			input    [width-1:0]    x1978_in,                     
			input    [width-1:0]    x1979_in,                     
			input    [width-1:0]    x1980_in,                     
			input    [width-1:0]    x1981_in,                     
			input    [width-1:0]    x1982_in,                     
			input    [width-1:0]    x1983_in,                     
			input    [width-1:0]    x1984_in,                     
			input    [width-1:0]    x1985_in,                     
			input    [width-1:0]    x1986_in,                     
			input    [width-1:0]    x1987_in,                     
			input    [width-1:0]    x1988_in,                     
			input    [width-1:0]    x1989_in,                     
			input    [width-1:0]    x1990_in,                     
			input    [width-1:0]    x1991_in,                     
			input    [width-1:0]    x1992_in,                     
			input    [width-1:0]    x1993_in,                     
			input    [width-1:0]    x1994_in,                     
			input    [width-1:0]    x1995_in,                     
			input    [width-1:0]    x1996_in,                     
			input    [width-1:0]    x1997_in,                     
			input    [width-1:0]    x1998_in,                     
			input    [width-1:0]    x1999_in,                     
			input    [width-1:0]    x2000_in,                     
			input    [width-1:0]    x2001_in,                     
			input    [width-1:0]    x2002_in,                     
			input    [width-1:0]    x2003_in,                     
			input    [width-1:0]    x2004_in,                     
			input    [width-1:0]    x2005_in,                     
			input    [width-1:0]    x2006_in,                     
			input    [width-1:0]    x2007_in,                     
			input    [width-1:0]    x2008_in,                     
			input    [width-1:0]    x2009_in,                     
			input    [width-1:0]    x2010_in,                     
			input    [width-1:0]    x2011_in,                     
			input    [width-1:0]    x2012_in,                     
			input    [width-1:0]    x2013_in,                     
			input    [width-1:0]    x2014_in,                     
			input    [width-1:0]    x2015_in,                     
			input    [width-1:0]    x2016_in,                     
			input    [width-1:0]    x2017_in,                     
			input    [width-1:0]    x2018_in,                     
			input    [width-1:0]    x2019_in,                     
			input    [width-1:0]    x2020_in,                     
			input    [width-1:0]    x2021_in,                     
			input    [width-1:0]    x2022_in,                     
			input    [width-1:0]    x2023_in,                     
			input    [width-1:0]    x2024_in,                     
			input    [width-1:0]    x2025_in,                     
			input    [width-1:0]    x2026_in,                     
			input    [width-1:0]    x2027_in,                     
			input    [width-1:0]    x2028_in,                     
			input    [width-1:0]    x2029_in,                     
			input    [width-1:0]    x2030_in,                     
			input    [width-1:0]    x2031_in,                     
			input    [width-1:0]    x2032_in,                     
			input    [width-1:0]    x2033_in,                     
			input    [width-1:0]    x2034_in,                     
			input    [width-1:0]    x2035_in,                     
			input    [width-1:0]    x2036_in,                     
			input    [width-1:0]    x2037_in,                     
			input    [width-1:0]    x2038_in,                     
			input    [width-1:0]    x2039_in,                     
			input    [width-1:0]    x2040_in,                     
			input    [width-1:0]    x2041_in,                     
			input    [width-1:0]    x2042_in,                     
			input    [width-1:0]    x2043_in,                     
			input    [width-1:0]    x2044_in,                     
			input    [width-1:0]    x2045_in,                     
			input    [width-1:0]    x2046_in,                     
			input    [width-1:0]    x2047_in,                     
		//--- outputs
			output                  stall_out,                    
			output   [width-1:0]    x0_out,                       
			output   [width-1:0]    x1_out,                       
			output   [width-1:0]    x2_out,                       
			output   [width-1:0]    x3_out,                       
			output   [width-1:0]    x4_out,                       
			output   [width-1:0]    x5_out,                       
			output   [width-1:0]    x6_out,                       
			output   [width-1:0]    x7_out,                       
			output   [width-1:0]    x8_out,                       
			output   [width-1:0]    x9_out,                       
			output   [width-1:0]    x10_out,                      
			output   [width-1:0]    x11_out,                      
			output   [width-1:0]    x12_out,                      
			output   [width-1:0]    x13_out,                      
			output   [width-1:0]    x14_out,                      
			output   [width-1:0]    x15_out,                      
			output   [width-1:0]    x16_out,                      
			output   [width-1:0]    x17_out,                      
			output   [width-1:0]    x18_out,                      
			output   [width-1:0]    x19_out,                      
			output   [width-1:0]    x20_out,                      
			output   [width-1:0]    x21_out,                      
			output   [width-1:0]    x22_out,                      
			output   [width-1:0]    x23_out,                      
			output   [width-1:0]    x24_out,                      
			output   [width-1:0]    x25_out,                      
			output   [width-1:0]    x26_out,                      
			output   [width-1:0]    x27_out,                      
			output   [width-1:0]    x28_out,                      
			output   [width-1:0]    x29_out,                      
			output   [width-1:0]    x30_out,                      
			output   [width-1:0]    x31_out,                      
			output   [width-1:0]    x32_out,                      
			output   [width-1:0]    x33_out,                      
			output   [width-1:0]    x34_out,                      
			output   [width-1:0]    x35_out,                      
			output   [width-1:0]    x36_out,                      
			output   [width-1:0]    x37_out,                      
			output   [width-1:0]    x38_out,                      
			output   [width-1:0]    x39_out,                      
			output   [width-1:0]    x40_out,                      
			output   [width-1:0]    x41_out,                      
			output   [width-1:0]    x42_out,                      
			output   [width-1:0]    x43_out,                      
			output   [width-1:0]    x44_out,                      
			output   [width-1:0]    x45_out,                      
			output   [width-1:0]    x46_out,                      
			output   [width-1:0]    x47_out,                      
			output   [width-1:0]    x48_out,                      
			output   [width-1:0]    x49_out,                      
			output   [width-1:0]    x50_out,                      
			output   [width-1:0]    x51_out,                      
			output   [width-1:0]    x52_out,                      
			output   [width-1:0]    x53_out,                      
			output   [width-1:0]    x54_out,                      
			output   [width-1:0]    x55_out,                      
			output   [width-1:0]    x56_out,                      
			output   [width-1:0]    x57_out,                      
			output   [width-1:0]    x58_out,                      
			output   [width-1:0]    x59_out,                      
			output   [width-1:0]    x60_out,                      
			output   [width-1:0]    x61_out,                      
			output   [width-1:0]    x62_out,                      
			output   [width-1:0]    x63_out,                      
			output   [width-1:0]    x64_out,                      
			output   [width-1:0]    x65_out,                      
			output   [width-1:0]    x66_out,                      
			output   [width-1:0]    x67_out,                      
			output   [width-1:0]    x68_out,                      
			output   [width-1:0]    x69_out,                      
			output   [width-1:0]    x70_out,                      
			output   [width-1:0]    x71_out,                      
			output   [width-1:0]    x72_out,                      
			output   [width-1:0]    x73_out,                      
			output   [width-1:0]    x74_out,                      
			output   [width-1:0]    x75_out,                      
			output   [width-1:0]    x76_out,                      
			output   [width-1:0]    x77_out,                      
			output   [width-1:0]    x78_out,                      
			output   [width-1:0]    x79_out,                      
			output   [width-1:0]    x80_out,                      
			output   [width-1:0]    x81_out,                      
			output   [width-1:0]    x82_out,                      
			output   [width-1:0]    x83_out,                      
			output   [width-1:0]    x84_out,                      
			output   [width-1:0]    x85_out,                      
			output   [width-1:0]    x86_out,                      
			output   [width-1:0]    x87_out,                      
			output   [width-1:0]    x88_out,                      
			output   [width-1:0]    x89_out,                      
			output   [width-1:0]    x90_out,                      
			output   [width-1:0]    x91_out,                      
			output   [width-1:0]    x92_out,                      
			output   [width-1:0]    x93_out,                      
			output   [width-1:0]    x94_out,                      
			output   [width-1:0]    x95_out,                      
			output   [width-1:0]    x96_out,                      
			output   [width-1:0]    x97_out,                      
			output   [width-1:0]    x98_out,                      
			output   [width-1:0]    x99_out,                      
			output   [width-1:0]    x100_out,                     
			output   [width-1:0]    x101_out,                     
			output   [width-1:0]    x102_out,                     
			output   [width-1:0]    x103_out,                     
			output   [width-1:0]    x104_out,                     
			output   [width-1:0]    x105_out,                     
			output   [width-1:0]    x106_out,                     
			output   [width-1:0]    x107_out,                     
			output   [width-1:0]    x108_out,                     
			output   [width-1:0]    x109_out,                     
			output   [width-1:0]    x110_out,                     
			output   [width-1:0]    x111_out,                     
			output   [width-1:0]    x112_out,                     
			output   [width-1:0]    x113_out,                     
			output   [width-1:0]    x114_out,                     
			output   [width-1:0]    x115_out,                     
			output   [width-1:0]    x116_out,                     
			output   [width-1:0]    x117_out,                     
			output   [width-1:0]    x118_out,                     
			output   [width-1:0]    x119_out,                     
			output   [width-1:0]    x120_out,                     
			output   [width-1:0]    x121_out,                     
			output   [width-1:0]    x122_out,                     
			output   [width-1:0]    x123_out,                     
			output   [width-1:0]    x124_out,                     
			output   [width-1:0]    x125_out,                     
			output   [width-1:0]    x126_out,                     
			output   [width-1:0]    x127_out,                     
			output   [width-1:0]    x128_out,                     
			output   [width-1:0]    x129_out,                     
			output   [width-1:0]    x130_out,                     
			output   [width-1:0]    x131_out,                     
			output   [width-1:0]    x132_out,                     
			output   [width-1:0]    x133_out,                     
			output   [width-1:0]    x134_out,                     
			output   [width-1:0]    x135_out,                     
			output   [width-1:0]    x136_out,                     
			output   [width-1:0]    x137_out,                     
			output   [width-1:0]    x138_out,                     
			output   [width-1:0]    x139_out,                     
			output   [width-1:0]    x140_out,                     
			output   [width-1:0]    x141_out,                     
			output   [width-1:0]    x142_out,                     
			output   [width-1:0]    x143_out,                     
			output   [width-1:0]    x144_out,                     
			output   [width-1:0]    x145_out,                     
			output   [width-1:0]    x146_out,                     
			output   [width-1:0]    x147_out,                     
			output   [width-1:0]    x148_out,                     
			output   [width-1:0]    x149_out,                     
			output   [width-1:0]    x150_out,                     
			output   [width-1:0]    x151_out,                     
			output   [width-1:0]    x152_out,                     
			output   [width-1:0]    x153_out,                     
			output   [width-1:0]    x154_out,                     
			output   [width-1:0]    x155_out,                     
			output   [width-1:0]    x156_out,                     
			output   [width-1:0]    x157_out,                     
			output   [width-1:0]    x158_out,                     
			output   [width-1:0]    x159_out,                     
			output   [width-1:0]    x160_out,                     
			output   [width-1:0]    x161_out,                     
			output   [width-1:0]    x162_out,                     
			output   [width-1:0]    x163_out,                     
			output   [width-1:0]    x164_out,                     
			output   [width-1:0]    x165_out,                     
			output   [width-1:0]    x166_out,                     
			output   [width-1:0]    x167_out,                     
			output   [width-1:0]    x168_out,                     
			output   [width-1:0]    x169_out,                     
			output   [width-1:0]    x170_out,                     
			output   [width-1:0]    x171_out,                     
			output   [width-1:0]    x172_out,                     
			output   [width-1:0]    x173_out,                     
			output   [width-1:0]    x174_out,                     
			output   [width-1:0]    x175_out,                     
			output   [width-1:0]    x176_out,                     
			output   [width-1:0]    x177_out,                     
			output   [width-1:0]    x178_out,                     
			output   [width-1:0]    x179_out,                     
			output   [width-1:0]    x180_out,                     
			output   [width-1:0]    x181_out,                     
			output   [width-1:0]    x182_out,                     
			output   [width-1:0]    x183_out,                     
			output   [width-1:0]    x184_out,                     
			output   [width-1:0]    x185_out,                     
			output   [width-1:0]    x186_out,                     
			output   [width-1:0]    x187_out,                     
			output   [width-1:0]    x188_out,                     
			output   [width-1:0]    x189_out,                     
			output   [width-1:0]    x190_out,                     
			output   [width-1:0]    x191_out,                     
			output   [width-1:0]    x192_out,                     
			output   [width-1:0]    x193_out,                     
			output   [width-1:0]    x194_out,                     
			output   [width-1:0]    x195_out,                     
			output   [width-1:0]    x196_out,                     
			output   [width-1:0]    x197_out,                     
			output   [width-1:0]    x198_out,                     
			output   [width-1:0]    x199_out,                     
			output   [width-1:0]    x200_out,                     
			output   [width-1:0]    x201_out,                     
			output   [width-1:0]    x202_out,                     
			output   [width-1:0]    x203_out,                     
			output   [width-1:0]    x204_out,                     
			output   [width-1:0]    x205_out,                     
			output   [width-1:0]    x206_out,                     
			output   [width-1:0]    x207_out,                     
			output   [width-1:0]    x208_out,                     
			output   [width-1:0]    x209_out,                     
			output   [width-1:0]    x210_out,                     
			output   [width-1:0]    x211_out,                     
			output   [width-1:0]    x212_out,                     
			output   [width-1:0]    x213_out,                     
			output   [width-1:0]    x214_out,                     
			output   [width-1:0]    x215_out,                     
			output   [width-1:0]    x216_out,                     
			output   [width-1:0]    x217_out,                     
			output   [width-1:0]    x218_out,                     
			output   [width-1:0]    x219_out,                     
			output   [width-1:0]    x220_out,                     
			output   [width-1:0]    x221_out,                     
			output   [width-1:0]    x222_out,                     
			output   [width-1:0]    x223_out,                     
			output   [width-1:0]    x224_out,                     
			output   [width-1:0]    x225_out,                     
			output   [width-1:0]    x226_out,                     
			output   [width-1:0]    x227_out,                     
			output   [width-1:0]    x228_out,                     
			output   [width-1:0]    x229_out,                     
			output   [width-1:0]    x230_out,                     
			output   [width-1:0]    x231_out,                     
			output   [width-1:0]    x232_out,                     
			output   [width-1:0]    x233_out,                     
			output   [width-1:0]    x234_out,                     
			output   [width-1:0]    x235_out,                     
			output   [width-1:0]    x236_out,                     
			output   [width-1:0]    x237_out,                     
			output   [width-1:0]    x238_out,                     
			output   [width-1:0]    x239_out,                     
			output   [width-1:0]    x240_out,                     
			output   [width-1:0]    x241_out,                     
			output   [width-1:0]    x242_out,                     
			output   [width-1:0]    x243_out,                     
			output   [width-1:0]    x244_out,                     
			output   [width-1:0]    x245_out,                     
			output   [width-1:0]    x246_out,                     
			output   [width-1:0]    x247_out,                     
			output   [width-1:0]    x248_out,                     
			output   [width-1:0]    x249_out,                     
			output   [width-1:0]    x250_out,                     
			output   [width-1:0]    x251_out,                     
			output   [width-1:0]    x252_out,                     
			output   [width-1:0]    x253_out,                     
			output   [width-1:0]    x254_out,                     
			output   [width-1:0]    x255_out,                     
			output   [width-1:0]    x256_out,                     
			output   [width-1:0]    x257_out,                     
			output   [width-1:0]    x258_out,                     
			output   [width-1:0]    x259_out,                     
			output   [width-1:0]    x260_out,                     
			output   [width-1:0]    x261_out,                     
			output   [width-1:0]    x262_out,                     
			output   [width-1:0]    x263_out,                     
			output   [width-1:0]    x264_out,                     
			output   [width-1:0]    x265_out,                     
			output   [width-1:0]    x266_out,                     
			output   [width-1:0]    x267_out,                     
			output   [width-1:0]    x268_out,                     
			output   [width-1:0]    x269_out,                     
			output   [width-1:0]    x270_out,                     
			output   [width-1:0]    x271_out,                     
			output   [width-1:0]    x272_out,                     
			output   [width-1:0]    x273_out,                     
			output   [width-1:0]    x274_out,                     
			output   [width-1:0]    x275_out,                     
			output   [width-1:0]    x276_out,                     
			output   [width-1:0]    x277_out,                     
			output   [width-1:0]    x278_out,                     
			output   [width-1:0]    x279_out,                     
			output   [width-1:0]    x280_out,                     
			output   [width-1:0]    x281_out,                     
			output   [width-1:0]    x282_out,                     
			output   [width-1:0]    x283_out,                     
			output   [width-1:0]    x284_out,                     
			output   [width-1:0]    x285_out,                     
			output   [width-1:0]    x286_out,                     
			output   [width-1:0]    x287_out,                     
			output   [width-1:0]    x288_out,                     
			output   [width-1:0]    x289_out,                     
			output   [width-1:0]    x290_out,                     
			output   [width-1:0]    x291_out,                     
			output   [width-1:0]    x292_out,                     
			output   [width-1:0]    x293_out,                     
			output   [width-1:0]    x294_out,                     
			output   [width-1:0]    x295_out,                     
			output   [width-1:0]    x296_out,                     
			output   [width-1:0]    x297_out,                     
			output   [width-1:0]    x298_out,                     
			output   [width-1:0]    x299_out,                     
			output   [width-1:0]    x300_out,                     
			output   [width-1:0]    x301_out,                     
			output   [width-1:0]    x302_out,                     
			output   [width-1:0]    x303_out,                     
			output   [width-1:0]    x304_out,                     
			output   [width-1:0]    x305_out,                     
			output   [width-1:0]    x306_out,                     
			output   [width-1:0]    x307_out,                     
			output   [width-1:0]    x308_out,                     
			output   [width-1:0]    x309_out,                     
			output   [width-1:0]    x310_out,                     
			output   [width-1:0]    x311_out,                     
			output   [width-1:0]    x312_out,                     
			output   [width-1:0]    x313_out,                     
			output   [width-1:0]    x314_out,                     
			output   [width-1:0]    x315_out,                     
			output   [width-1:0]    x316_out,                     
			output   [width-1:0]    x317_out,                     
			output   [width-1:0]    x318_out,                     
			output   [width-1:0]    x319_out,                     
			output   [width-1:0]    x320_out,                     
			output   [width-1:0]    x321_out,                     
			output   [width-1:0]    x322_out,                     
			output   [width-1:0]    x323_out,                     
			output   [width-1:0]    x324_out,                     
			output   [width-1:0]    x325_out,                     
			output   [width-1:0]    x326_out,                     
			output   [width-1:0]    x327_out,                     
			output   [width-1:0]    x328_out,                     
			output   [width-1:0]    x329_out,                     
			output   [width-1:0]    x330_out,                     
			output   [width-1:0]    x331_out,                     
			output   [width-1:0]    x332_out,                     
			output   [width-1:0]    x333_out,                     
			output   [width-1:0]    x334_out,                     
			output   [width-1:0]    x335_out,                     
			output   [width-1:0]    x336_out,                     
			output   [width-1:0]    x337_out,                     
			output   [width-1:0]    x338_out,                     
			output   [width-1:0]    x339_out,                     
			output   [width-1:0]    x340_out,                     
			output   [width-1:0]    x341_out,                     
			output   [width-1:0]    x342_out,                     
			output   [width-1:0]    x343_out,                     
			output   [width-1:0]    x344_out,                     
			output   [width-1:0]    x345_out,                     
			output   [width-1:0]    x346_out,                     
			output   [width-1:0]    x347_out,                     
			output   [width-1:0]    x348_out,                     
			output   [width-1:0]    x349_out,                     
			output   [width-1:0]    x350_out,                     
			output   [width-1:0]    x351_out,                     
			output   [width-1:0]    x352_out,                     
			output   [width-1:0]    x353_out,                     
			output   [width-1:0]    x354_out,                     
			output   [width-1:0]    x355_out,                     
			output   [width-1:0]    x356_out,                     
			output   [width-1:0]    x357_out,                     
			output   [width-1:0]    x358_out,                     
			output   [width-1:0]    x359_out,                     
			output   [width-1:0]    x360_out,                     
			output   [width-1:0]    x361_out,                     
			output   [width-1:0]    x362_out,                     
			output   [width-1:0]    x363_out,                     
			output   [width-1:0]    x364_out,                     
			output   [width-1:0]    x365_out,                     
			output   [width-1:0]    x366_out,                     
			output   [width-1:0]    x367_out,                     
			output   [width-1:0]    x368_out,                     
			output   [width-1:0]    x369_out,                     
			output   [width-1:0]    x370_out,                     
			output   [width-1:0]    x371_out,                     
			output   [width-1:0]    x372_out,                     
			output   [width-1:0]    x373_out,                     
			output   [width-1:0]    x374_out,                     
			output   [width-1:0]    x375_out,                     
			output   [width-1:0]    x376_out,                     
			output   [width-1:0]    x377_out,                     
			output   [width-1:0]    x378_out,                     
			output   [width-1:0]    x379_out,                     
			output   [width-1:0]    x380_out,                     
			output   [width-1:0]    x381_out,                     
			output   [width-1:0]    x382_out,                     
			output   [width-1:0]    x383_out,                     
			output   [width-1:0]    x384_out,                     
			output   [width-1:0]    x385_out,                     
			output   [width-1:0]    x386_out,                     
			output   [width-1:0]    x387_out,                     
			output   [width-1:0]    x388_out,                     
			output   [width-1:0]    x389_out,                     
			output   [width-1:0]    x390_out,                     
			output   [width-1:0]    x391_out,                     
			output   [width-1:0]    x392_out,                     
			output   [width-1:0]    x393_out,                     
			output   [width-1:0]    x394_out,                     
			output   [width-1:0]    x395_out,                     
			output   [width-1:0]    x396_out,                     
			output   [width-1:0]    x397_out,                     
			output   [width-1:0]    x398_out,                     
			output   [width-1:0]    x399_out,                     
			output   [width-1:0]    x400_out,                     
			output   [width-1:0]    x401_out,                     
			output   [width-1:0]    x402_out,                     
			output   [width-1:0]    x403_out,                     
			output   [width-1:0]    x404_out,                     
			output   [width-1:0]    x405_out,                     
			output   [width-1:0]    x406_out,                     
			output   [width-1:0]    x407_out,                     
			output   [width-1:0]    x408_out,                     
			output   [width-1:0]    x409_out,                     
			output   [width-1:0]    x410_out,                     
			output   [width-1:0]    x411_out,                     
			output   [width-1:0]    x412_out,                     
			output   [width-1:0]    x413_out,                     
			output   [width-1:0]    x414_out,                     
			output   [width-1:0]    x415_out,                     
			output   [width-1:0]    x416_out,                     
			output   [width-1:0]    x417_out,                     
			output   [width-1:0]    x418_out,                     
			output   [width-1:0]    x419_out,                     
			output   [width-1:0]    x420_out,                     
			output   [width-1:0]    x421_out,                     
			output   [width-1:0]    x422_out,                     
			output   [width-1:0]    x423_out,                     
			output   [width-1:0]    x424_out,                     
			output   [width-1:0]    x425_out,                     
			output   [width-1:0]    x426_out,                     
			output   [width-1:0]    x427_out,                     
			output   [width-1:0]    x428_out,                     
			output   [width-1:0]    x429_out,                     
			output   [width-1:0]    x430_out,                     
			output   [width-1:0]    x431_out,                     
			output   [width-1:0]    x432_out,                     
			output   [width-1:0]    x433_out,                     
			output   [width-1:0]    x434_out,                     
			output   [width-1:0]    x435_out,                     
			output   [width-1:0]    x436_out,                     
			output   [width-1:0]    x437_out,                     
			output   [width-1:0]    x438_out,                     
			output   [width-1:0]    x439_out,                     
			output   [width-1:0]    x440_out,                     
			output   [width-1:0]    x441_out,                     
			output   [width-1:0]    x442_out,                     
			output   [width-1:0]    x443_out,                     
			output   [width-1:0]    x444_out,                     
			output   [width-1:0]    x445_out,                     
			output   [width-1:0]    x446_out,                     
			output   [width-1:0]    x447_out,                     
			output   [width-1:0]    x448_out,                     
			output   [width-1:0]    x449_out,                     
			output   [width-1:0]    x450_out,                     
			output   [width-1:0]    x451_out,                     
			output   [width-1:0]    x452_out,                     
			output   [width-1:0]    x453_out,                     
			output   [width-1:0]    x454_out,                     
			output   [width-1:0]    x455_out,                     
			output   [width-1:0]    x456_out,                     
			output   [width-1:0]    x457_out,                     
			output   [width-1:0]    x458_out,                     
			output   [width-1:0]    x459_out,                     
			output   [width-1:0]    x460_out,                     
			output   [width-1:0]    x461_out,                     
			output   [width-1:0]    x462_out,                     
			output   [width-1:0]    x463_out,                     
			output   [width-1:0]    x464_out,                     
			output   [width-1:0]    x465_out,                     
			output   [width-1:0]    x466_out,                     
			output   [width-1:0]    x467_out,                     
			output   [width-1:0]    x468_out,                     
			output   [width-1:0]    x469_out,                     
			output   [width-1:0]    x470_out,                     
			output   [width-1:0]    x471_out,                     
			output   [width-1:0]    x472_out,                     
			output   [width-1:0]    x473_out,                     
			output   [width-1:0]    x474_out,                     
			output   [width-1:0]    x475_out,                     
			output   [width-1:0]    x476_out,                     
			output   [width-1:0]    x477_out,                     
			output   [width-1:0]    x478_out,                     
			output   [width-1:0]    x479_out,                     
			output   [width-1:0]    x480_out,                     
			output   [width-1:0]    x481_out,                     
			output   [width-1:0]    x482_out,                     
			output   [width-1:0]    x483_out,                     
			output   [width-1:0]    x484_out,                     
			output   [width-1:0]    x485_out,                     
			output   [width-1:0]    x486_out,                     
			output   [width-1:0]    x487_out,                     
			output   [width-1:0]    x488_out,                     
			output   [width-1:0]    x489_out,                     
			output   [width-1:0]    x490_out,                     
			output   [width-1:0]    x491_out,                     
			output   [width-1:0]    x492_out,                     
			output   [width-1:0]    x493_out,                     
			output   [width-1:0]    x494_out,                     
			output   [width-1:0]    x495_out,                     
			output   [width-1:0]    x496_out,                     
			output   [width-1:0]    x497_out,                     
			output   [width-1:0]    x498_out,                     
			output   [width-1:0]    x499_out,                     
			output   [width-1:0]    x500_out,                     
			output   [width-1:0]    x501_out,                     
			output   [width-1:0]    x502_out,                     
			output   [width-1:0]    x503_out,                     
			output   [width-1:0]    x504_out,                     
			output   [width-1:0]    x505_out,                     
			output   [width-1:0]    x506_out,                     
			output   [width-1:0]    x507_out,                     
			output   [width-1:0]    x508_out,                     
			output   [width-1:0]    x509_out,                     
			output   [width-1:0]    x510_out,                     
			output   [width-1:0]    x511_out,                     
			output   [width-1:0]    x512_out,                     
			output   [width-1:0]    x513_out,                     
			output   [width-1:0]    x514_out,                     
			output   [width-1:0]    x515_out,                     
			output   [width-1:0]    x516_out,                     
			output   [width-1:0]    x517_out,                     
			output   [width-1:0]    x518_out,                     
			output   [width-1:0]    x519_out,                     
			output   [width-1:0]    x520_out,                     
			output   [width-1:0]    x521_out,                     
			output   [width-1:0]    x522_out,                     
			output   [width-1:0]    x523_out,                     
			output   [width-1:0]    x524_out,                     
			output   [width-1:0]    x525_out,                     
			output   [width-1:0]    x526_out,                     
			output   [width-1:0]    x527_out,                     
			output   [width-1:0]    x528_out,                     
			output   [width-1:0]    x529_out,                     
			output   [width-1:0]    x530_out,                     
			output   [width-1:0]    x531_out,                     
			output   [width-1:0]    x532_out,                     
			output   [width-1:0]    x533_out,                     
			output   [width-1:0]    x534_out,                     
			output   [width-1:0]    x535_out,                     
			output   [width-1:0]    x536_out,                     
			output   [width-1:0]    x537_out,                     
			output   [width-1:0]    x538_out,                     
			output   [width-1:0]    x539_out,                     
			output   [width-1:0]    x540_out,                     
			output   [width-1:0]    x541_out,                     
			output   [width-1:0]    x542_out,                     
			output   [width-1:0]    x543_out,                     
			output   [width-1:0]    x544_out,                     
			output   [width-1:0]    x545_out,                     
			output   [width-1:0]    x546_out,                     
			output   [width-1:0]    x547_out,                     
			output   [width-1:0]    x548_out,                     
			output   [width-1:0]    x549_out,                     
			output   [width-1:0]    x550_out,                     
			output   [width-1:0]    x551_out,                     
			output   [width-1:0]    x552_out,                     
			output   [width-1:0]    x553_out,                     
			output   [width-1:0]    x554_out,                     
			output   [width-1:0]    x555_out,                     
			output   [width-1:0]    x556_out,                     
			output   [width-1:0]    x557_out,                     
			output   [width-1:0]    x558_out,                     
			output   [width-1:0]    x559_out,                     
			output   [width-1:0]    x560_out,                     
			output   [width-1:0]    x561_out,                     
			output   [width-1:0]    x562_out,                     
			output   [width-1:0]    x563_out,                     
			output   [width-1:0]    x564_out,                     
			output   [width-1:0]    x565_out,                     
			output   [width-1:0]    x566_out,                     
			output   [width-1:0]    x567_out,                     
			output   [width-1:0]    x568_out,                     
			output   [width-1:0]    x569_out,                     
			output   [width-1:0]    x570_out,                     
			output   [width-1:0]    x571_out,                     
			output   [width-1:0]    x572_out,                     
			output   [width-1:0]    x573_out,                     
			output   [width-1:0]    x574_out,                     
			output   [width-1:0]    x575_out,                     
			output   [width-1:0]    x576_out,                     
			output   [width-1:0]    x577_out,                     
			output   [width-1:0]    x578_out,                     
			output   [width-1:0]    x579_out,                     
			output   [width-1:0]    x580_out,                     
			output   [width-1:0]    x581_out,                     
			output   [width-1:0]    x582_out,                     
			output   [width-1:0]    x583_out,                     
			output   [width-1:0]    x584_out,                     
			output   [width-1:0]    x585_out,                     
			output   [width-1:0]    x586_out,                     
			output   [width-1:0]    x587_out,                     
			output   [width-1:0]    x588_out,                     
			output   [width-1:0]    x589_out,                     
			output   [width-1:0]    x590_out,                     
			output   [width-1:0]    x591_out,                     
			output   [width-1:0]    x592_out,                     
			output   [width-1:0]    x593_out,                     
			output   [width-1:0]    x594_out,                     
			output   [width-1:0]    x595_out,                     
			output   [width-1:0]    x596_out,                     
			output   [width-1:0]    x597_out,                     
			output   [width-1:0]    x598_out,                     
			output   [width-1:0]    x599_out,                     
			output   [width-1:0]    x600_out,                     
			output   [width-1:0]    x601_out,                     
			output   [width-1:0]    x602_out,                     
			output   [width-1:0]    x603_out,                     
			output   [width-1:0]    x604_out,                     
			output   [width-1:0]    x605_out,                     
			output   [width-1:0]    x606_out,                     
			output   [width-1:0]    x607_out,                     
			output   [width-1:0]    x608_out,                     
			output   [width-1:0]    x609_out,                     
			output   [width-1:0]    x610_out,                     
			output   [width-1:0]    x611_out,                     
			output   [width-1:0]    x612_out,                     
			output   [width-1:0]    x613_out,                     
			output   [width-1:0]    x614_out,                     
			output   [width-1:0]    x615_out,                     
			output   [width-1:0]    x616_out,                     
			output   [width-1:0]    x617_out,                     
			output   [width-1:0]    x618_out,                     
			output   [width-1:0]    x619_out,                     
			output   [width-1:0]    x620_out,                     
			output   [width-1:0]    x621_out,                     
			output   [width-1:0]    x622_out,                     
			output   [width-1:0]    x623_out,                     
			output   [width-1:0]    x624_out,                     
			output   [width-1:0]    x625_out,                     
			output   [width-1:0]    x626_out,                     
			output   [width-1:0]    x627_out,                     
			output   [width-1:0]    x628_out,                     
			output   [width-1:0]    x629_out,                     
			output   [width-1:0]    x630_out,                     
			output   [width-1:0]    x631_out,                     
			output   [width-1:0]    x632_out,                     
			output   [width-1:0]    x633_out,                     
			output   [width-1:0]    x634_out,                     
			output   [width-1:0]    x635_out,                     
			output   [width-1:0]    x636_out,                     
			output   [width-1:0]    x637_out,                     
			output   [width-1:0]    x638_out,                     
			output   [width-1:0]    x639_out,                     
			output   [width-1:0]    x640_out,                     
			output   [width-1:0]    x641_out,                     
			output   [width-1:0]    x642_out,                     
			output   [width-1:0]    x643_out,                     
			output   [width-1:0]    x644_out,                     
			output   [width-1:0]    x645_out,                     
			output   [width-1:0]    x646_out,                     
			output   [width-1:0]    x647_out,                     
			output   [width-1:0]    x648_out,                     
			output   [width-1:0]    x649_out,                     
			output   [width-1:0]    x650_out,                     
			output   [width-1:0]    x651_out,                     
			output   [width-1:0]    x652_out,                     
			output   [width-1:0]    x653_out,                     
			output   [width-1:0]    x654_out,                     
			output   [width-1:0]    x655_out,                     
			output   [width-1:0]    x656_out,                     
			output   [width-1:0]    x657_out,                     
			output   [width-1:0]    x658_out,                     
			output   [width-1:0]    x659_out,                     
			output   [width-1:0]    x660_out,                     
			output   [width-1:0]    x661_out,                     
			output   [width-1:0]    x662_out,                     
			output   [width-1:0]    x663_out,                     
			output   [width-1:0]    x664_out,                     
			output   [width-1:0]    x665_out,                     
			output   [width-1:0]    x666_out,                     
			output   [width-1:0]    x667_out,                     
			output   [width-1:0]    x668_out,                     
			output   [width-1:0]    x669_out,                     
			output   [width-1:0]    x670_out,                     
			output   [width-1:0]    x671_out,                     
			output   [width-1:0]    x672_out,                     
			output   [width-1:0]    x673_out,                     
			output   [width-1:0]    x674_out,                     
			output   [width-1:0]    x675_out,                     
			output   [width-1:0]    x676_out,                     
			output   [width-1:0]    x677_out,                     
			output   [width-1:0]    x678_out,                     
			output   [width-1:0]    x679_out,                     
			output   [width-1:0]    x680_out,                     
			output   [width-1:0]    x681_out,                     
			output   [width-1:0]    x682_out,                     
			output   [width-1:0]    x683_out,                     
			output   [width-1:0]    x684_out,                     
			output   [width-1:0]    x685_out,                     
			output   [width-1:0]    x686_out,                     
			output   [width-1:0]    x687_out,                     
			output   [width-1:0]    x688_out,                     
			output   [width-1:0]    x689_out,                     
			output   [width-1:0]    x690_out,                     
			output   [width-1:0]    x691_out,                     
			output   [width-1:0]    x692_out,                     
			output   [width-1:0]    x693_out,                     
			output   [width-1:0]    x694_out,                     
			output   [width-1:0]    x695_out,                     
			output   [width-1:0]    x696_out,                     
			output   [width-1:0]    x697_out,                     
			output   [width-1:0]    x698_out,                     
			output   [width-1:0]    x699_out,                     
			output   [width-1:0]    x700_out,                     
			output   [width-1:0]    x701_out,                     
			output   [width-1:0]    x702_out,                     
			output   [width-1:0]    x703_out,                     
			output   [width-1:0]    x704_out,                     
			output   [width-1:0]    x705_out,                     
			output   [width-1:0]    x706_out,                     
			output   [width-1:0]    x707_out,                     
			output   [width-1:0]    x708_out,                     
			output   [width-1:0]    x709_out,                     
			output   [width-1:0]    x710_out,                     
			output   [width-1:0]    x711_out,                     
			output   [width-1:0]    x712_out,                     
			output   [width-1:0]    x713_out,                     
			output   [width-1:0]    x714_out,                     
			output   [width-1:0]    x715_out,                     
			output   [width-1:0]    x716_out,                     
			output   [width-1:0]    x717_out,                     
			output   [width-1:0]    x718_out,                     
			output   [width-1:0]    x719_out,                     
			output   [width-1:0]    x720_out,                     
			output   [width-1:0]    x721_out,                     
			output   [width-1:0]    x722_out,                     
			output   [width-1:0]    x723_out,                     
			output   [width-1:0]    x724_out,                     
			output   [width-1:0]    x725_out,                     
			output   [width-1:0]    x726_out,                     
			output   [width-1:0]    x727_out,                     
			output   [width-1:0]    x728_out,                     
			output   [width-1:0]    x729_out,                     
			output   [width-1:0]    x730_out,                     
			output   [width-1:0]    x731_out,                     
			output   [width-1:0]    x732_out,                     
			output   [width-1:0]    x733_out,                     
			output   [width-1:0]    x734_out,                     
			output   [width-1:0]    x735_out,                     
			output   [width-1:0]    x736_out,                     
			output   [width-1:0]    x737_out,                     
			output   [width-1:0]    x738_out,                     
			output   [width-1:0]    x739_out,                     
			output   [width-1:0]    x740_out,                     
			output   [width-1:0]    x741_out,                     
			output   [width-1:0]    x742_out,                     
			output   [width-1:0]    x743_out,                     
			output   [width-1:0]    x744_out,                     
			output   [width-1:0]    x745_out,                     
			output   [width-1:0]    x746_out,                     
			output   [width-1:0]    x747_out,                     
			output   [width-1:0]    x748_out,                     
			output   [width-1:0]    x749_out,                     
			output   [width-1:0]    x750_out,                     
			output   [width-1:0]    x751_out,                     
			output   [width-1:0]    x752_out,                     
			output   [width-1:0]    x753_out,                     
			output   [width-1:0]    x754_out,                     
			output   [width-1:0]    x755_out,                     
			output   [width-1:0]    x756_out,                     
			output   [width-1:0]    x757_out,                     
			output   [width-1:0]    x758_out,                     
			output   [width-1:0]    x759_out,                     
			output   [width-1:0]    x760_out,                     
			output   [width-1:0]    x761_out,                     
			output   [width-1:0]    x762_out,                     
			output   [width-1:0]    x763_out,                     
			output   [width-1:0]    x764_out,                     
			output   [width-1:0]    x765_out,                     
			output   [width-1:0]    x766_out,                     
			output   [width-1:0]    x767_out,                     
			output   [width-1:0]    x768_out,                     
			output   [width-1:0]    x769_out,                     
			output   [width-1:0]    x770_out,                     
			output   [width-1:0]    x771_out,                     
			output   [width-1:0]    x772_out,                     
			output   [width-1:0]    x773_out,                     
			output   [width-1:0]    x774_out,                     
			output   [width-1:0]    x775_out,                     
			output   [width-1:0]    x776_out,                     
			output   [width-1:0]    x777_out,                     
			output   [width-1:0]    x778_out,                     
			output   [width-1:0]    x779_out,                     
			output   [width-1:0]    x780_out,                     
			output   [width-1:0]    x781_out,                     
			output   [width-1:0]    x782_out,                     
			output   [width-1:0]    x783_out,                     
			output   [width-1:0]    x784_out,                     
			output   [width-1:0]    x785_out,                     
			output   [width-1:0]    x786_out,                     
			output   [width-1:0]    x787_out,                     
			output   [width-1:0]    x788_out,                     
			output   [width-1:0]    x789_out,                     
			output   [width-1:0]    x790_out,                     
			output   [width-1:0]    x791_out,                     
			output   [width-1:0]    x792_out,                     
			output   [width-1:0]    x793_out,                     
			output   [width-1:0]    x794_out,                     
			output   [width-1:0]    x795_out,                     
			output   [width-1:0]    x796_out,                     
			output   [width-1:0]    x797_out,                     
			output   [width-1:0]    x798_out,                     
			output   [width-1:0]    x799_out,                     
			output   [width-1:0]    x800_out,                     
			output   [width-1:0]    x801_out,                     
			output   [width-1:0]    x802_out,                     
			output   [width-1:0]    x803_out,                     
			output   [width-1:0]    x804_out,                     
			output   [width-1:0]    x805_out,                     
			output   [width-1:0]    x806_out,                     
			output   [width-1:0]    x807_out,                     
			output   [width-1:0]    x808_out,                     
			output   [width-1:0]    x809_out,                     
			output   [width-1:0]    x810_out,                     
			output   [width-1:0]    x811_out,                     
			output   [width-1:0]    x812_out,                     
			output   [width-1:0]    x813_out,                     
			output   [width-1:0]    x814_out,                     
			output   [width-1:0]    x815_out,                     
			output   [width-1:0]    x816_out,                     
			output   [width-1:0]    x817_out,                     
			output   [width-1:0]    x818_out,                     
			output   [width-1:0]    x819_out,                     
			output   [width-1:0]    x820_out,                     
			output   [width-1:0]    x821_out,                     
			output   [width-1:0]    x822_out,                     
			output   [width-1:0]    x823_out,                     
			output   [width-1:0]    x824_out,                     
			output   [width-1:0]    x825_out,                     
			output   [width-1:0]    x826_out,                     
			output   [width-1:0]    x827_out,                     
			output   [width-1:0]    x828_out,                     
			output   [width-1:0]    x829_out,                     
			output   [width-1:0]    x830_out,                     
			output   [width-1:0]    x831_out,                     
			output   [width-1:0]    x832_out,                     
			output   [width-1:0]    x833_out,                     
			output   [width-1:0]    x834_out,                     
			output   [width-1:0]    x835_out,                     
			output   [width-1:0]    x836_out,                     
			output   [width-1:0]    x837_out,                     
			output   [width-1:0]    x838_out,                     
			output   [width-1:0]    x839_out,                     
			output   [width-1:0]    x840_out,                     
			output   [width-1:0]    x841_out,                     
			output   [width-1:0]    x842_out,                     
			output   [width-1:0]    x843_out,                     
			output   [width-1:0]    x844_out,                     
			output   [width-1:0]    x845_out,                     
			output   [width-1:0]    x846_out,                     
			output   [width-1:0]    x847_out,                     
			output   [width-1:0]    x848_out,                     
			output   [width-1:0]    x849_out,                     
			output   [width-1:0]    x850_out,                     
			output   [width-1:0]    x851_out,                     
			output   [width-1:0]    x852_out,                     
			output   [width-1:0]    x853_out,                     
			output   [width-1:0]    x854_out,                     
			output   [width-1:0]    x855_out,                     
			output   [width-1:0]    x856_out,                     
			output   [width-1:0]    x857_out,                     
			output   [width-1:0]    x858_out,                     
			output   [width-1:0]    x859_out,                     
			output   [width-1:0]    x860_out,                     
			output   [width-1:0]    x861_out,                     
			output   [width-1:0]    x862_out,                     
			output   [width-1:0]    x863_out,                     
			output   [width-1:0]    x864_out,                     
			output   [width-1:0]    x865_out,                     
			output   [width-1:0]    x866_out,                     
			output   [width-1:0]    x867_out,                     
			output   [width-1:0]    x868_out,                     
			output   [width-1:0]    x869_out,                     
			output   [width-1:0]    x870_out,                     
			output   [width-1:0]    x871_out,                     
			output   [width-1:0]    x872_out,                     
			output   [width-1:0]    x873_out,                     
			output   [width-1:0]    x874_out,                     
			output   [width-1:0]    x875_out,                     
			output   [width-1:0]    x876_out,                     
			output   [width-1:0]    x877_out,                     
			output   [width-1:0]    x878_out,                     
			output   [width-1:0]    x879_out,                     
			output   [width-1:0]    x880_out,                     
			output   [width-1:0]    x881_out,                     
			output   [width-1:0]    x882_out,                     
			output   [width-1:0]    x883_out,                     
			output   [width-1:0]    x884_out,                     
			output   [width-1:0]    x885_out,                     
			output   [width-1:0]    x886_out,                     
			output   [width-1:0]    x887_out,                     
			output   [width-1:0]    x888_out,                     
			output   [width-1:0]    x889_out,                     
			output   [width-1:0]    x890_out,                     
			output   [width-1:0]    x891_out,                     
			output   [width-1:0]    x892_out,                     
			output   [width-1:0]    x893_out,                     
			output   [width-1:0]    x894_out,                     
			output   [width-1:0]    x895_out,                     
			output   [width-1:0]    x896_out,                     
			output   [width-1:0]    x897_out,                     
			output   [width-1:0]    x898_out,                     
			output   [width-1:0]    x899_out,                     
			output   [width-1:0]    x900_out,                     
			output   [width-1:0]    x901_out,                     
			output   [width-1:0]    x902_out,                     
			output   [width-1:0]    x903_out,                     
			output   [width-1:0]    x904_out,                     
			output   [width-1:0]    x905_out,                     
			output   [width-1:0]    x906_out,                     
			output   [width-1:0]    x907_out,                     
			output   [width-1:0]    x908_out,                     
			output   [width-1:0]    x909_out,                     
			output   [width-1:0]    x910_out,                     
			output   [width-1:0]    x911_out,                     
			output   [width-1:0]    x912_out,                     
			output   [width-1:0]    x913_out,                     
			output   [width-1:0]    x914_out,                     
			output   [width-1:0]    x915_out,                     
			output   [width-1:0]    x916_out,                     
			output   [width-1:0]    x917_out,                     
			output   [width-1:0]    x918_out,                     
			output   [width-1:0]    x919_out,                     
			output   [width-1:0]    x920_out,                     
			output   [width-1:0]    x921_out,                     
			output   [width-1:0]    x922_out,                     
			output   [width-1:0]    x923_out,                     
			output   [width-1:0]    x924_out,                     
			output   [width-1:0]    x925_out,                     
			output   [width-1:0]    x926_out,                     
			output   [width-1:0]    x927_out,                     
			output   [width-1:0]    x928_out,                     
			output   [width-1:0]    x929_out,                     
			output   [width-1:0]    x930_out,                     
			output   [width-1:0]    x931_out,                     
			output   [width-1:0]    x932_out,                     
			output   [width-1:0]    x933_out,                     
			output   [width-1:0]    x934_out,                     
			output   [width-1:0]    x935_out,                     
			output   [width-1:0]    x936_out,                     
			output   [width-1:0]    x937_out,                     
			output   [width-1:0]    x938_out,                     
			output   [width-1:0]    x939_out,                     
			output   [width-1:0]    x940_out,                     
			output   [width-1:0]    x941_out,                     
			output   [width-1:0]    x942_out,                     
			output   [width-1:0]    x943_out,                     
			output   [width-1:0]    x944_out,                     
			output   [width-1:0]    x945_out,                     
			output   [width-1:0]    x946_out,                     
			output   [width-1:0]    x947_out,                     
			output   [width-1:0]    x948_out,                     
			output   [width-1:0]    x949_out,                     
			output   [width-1:0]    x950_out,                     
			output   [width-1:0]    x951_out,                     
			output   [width-1:0]    x952_out,                     
			output   [width-1:0]    x953_out,                     
			output   [width-1:0]    x954_out,                     
			output   [width-1:0]    x955_out,                     
			output   [width-1:0]    x956_out,                     
			output   [width-1:0]    x957_out,                     
			output   [width-1:0]    x958_out,                     
			output   [width-1:0]    x959_out,                     
			output   [width-1:0]    x960_out,                     
			output   [width-1:0]    x961_out,                     
			output   [width-1:0]    x962_out,                     
			output   [width-1:0]    x963_out,                     
			output   [width-1:0]    x964_out,                     
			output   [width-1:0]    x965_out,                     
			output   [width-1:0]    x966_out,                     
			output   [width-1:0]    x967_out,                     
			output   [width-1:0]    x968_out,                     
			output   [width-1:0]    x969_out,                     
			output   [width-1:0]    x970_out,                     
			output   [width-1:0]    x971_out,                     
			output   [width-1:0]    x972_out,                     
			output   [width-1:0]    x973_out,                     
			output   [width-1:0]    x974_out,                     
			output   [width-1:0]    x975_out,                     
			output   [width-1:0]    x976_out,                     
			output   [width-1:0]    x977_out,                     
			output   [width-1:0]    x978_out,                     
			output   [width-1:0]    x979_out,                     
			output   [width-1:0]    x980_out,                     
			output   [width-1:0]    x981_out,                     
			output   [width-1:0]    x982_out,                     
			output   [width-1:0]    x983_out,                     
			output   [width-1:0]    x984_out,                     
			output   [width-1:0]    x985_out,                     
			output   [width-1:0]    x986_out,                     
			output   [width-1:0]    x987_out,                     
			output   [width-1:0]    x988_out,                     
			output   [width-1:0]    x989_out,                     
			output   [width-1:0]    x990_out,                     
			output   [width-1:0]    x991_out,                     
			output   [width-1:0]    x992_out,                     
			output   [width-1:0]    x993_out,                     
			output   [width-1:0]    x994_out,                     
			output   [width-1:0]    x995_out,                     
			output   [width-1:0]    x996_out,                     
			output   [width-1:0]    x997_out,                     
			output   [width-1:0]    x998_out,                     
			output   [width-1:0]    x999_out,                     
			output   [width-1:0]    x1000_out,                    
			output   [width-1:0]    x1001_out,                    
			output   [width-1:0]    x1002_out,                    
			output   [width-1:0]    x1003_out,                    
			output   [width-1:0]    x1004_out,                    
			output   [width-1:0]    x1005_out,                    
			output   [width-1:0]    x1006_out,                    
			output   [width-1:0]    x1007_out,                    
			output   [width-1:0]    x1008_out,                    
			output   [width-1:0]    x1009_out,                    
			output   [width-1:0]    x1010_out,                    
			output   [width-1:0]    x1011_out,                    
			output   [width-1:0]    x1012_out,                    
			output   [width-1:0]    x1013_out,                    
			output   [width-1:0]    x1014_out,                    
			output   [width-1:0]    x1015_out,                    
			output   [width-1:0]    x1016_out,                    
			output   [width-1:0]    x1017_out,                    
			output   [width-1:0]    x1018_out,                    
			output   [width-1:0]    x1019_out,                    
			output   [width-1:0]    x1020_out,                    
			output   [width-1:0]    x1021_out,                    
			output   [width-1:0]    x1022_out,                    
			output   [width-1:0]    x1023_out,                    
			output   [width-1:0]    x1024_out,                    
			output   [width-1:0]    x1025_out,                    
			output   [width-1:0]    x1026_out,                    
			output   [width-1:0]    x1027_out,                    
			output   [width-1:0]    x1028_out,                    
			output   [width-1:0]    x1029_out,                    
			output   [width-1:0]    x1030_out,                    
			output   [width-1:0]    x1031_out,                    
			output   [width-1:0]    x1032_out,                    
			output   [width-1:0]    x1033_out,                    
			output   [width-1:0]    x1034_out,                    
			output   [width-1:0]    x1035_out,                    
			output   [width-1:0]    x1036_out,                    
			output   [width-1:0]    x1037_out,                    
			output   [width-1:0]    x1038_out,                    
			output   [width-1:0]    x1039_out,                    
			output   [width-1:0]    x1040_out,                    
			output   [width-1:0]    x1041_out,                    
			output   [width-1:0]    x1042_out,                    
			output   [width-1:0]    x1043_out,                    
			output   [width-1:0]    x1044_out,                    
			output   [width-1:0]    x1045_out,                    
			output   [width-1:0]    x1046_out,                    
			output   [width-1:0]    x1047_out,                    
			output   [width-1:0]    x1048_out,                    
			output   [width-1:0]    x1049_out,                    
			output   [width-1:0]    x1050_out,                    
			output   [width-1:0]    x1051_out,                    
			output   [width-1:0]    x1052_out,                    
			output   [width-1:0]    x1053_out,                    
			output   [width-1:0]    x1054_out,                    
			output   [width-1:0]    x1055_out,                    
			output   [width-1:0]    x1056_out,                    
			output   [width-1:0]    x1057_out,                    
			output   [width-1:0]    x1058_out,                    
			output   [width-1:0]    x1059_out,                    
			output   [width-1:0]    x1060_out,                    
			output   [width-1:0]    x1061_out,                    
			output   [width-1:0]    x1062_out,                    
			output   [width-1:0]    x1063_out,                    
			output   [width-1:0]    x1064_out,                    
			output   [width-1:0]    x1065_out,                    
			output   [width-1:0]    x1066_out,                    
			output   [width-1:0]    x1067_out,                    
			output   [width-1:0]    x1068_out,                    
			output   [width-1:0]    x1069_out,                    
			output   [width-1:0]    x1070_out,                    
			output   [width-1:0]    x1071_out,                    
			output   [width-1:0]    x1072_out,                    
			output   [width-1:0]    x1073_out,                    
			output   [width-1:0]    x1074_out,                    
			output   [width-1:0]    x1075_out,                    
			output   [width-1:0]    x1076_out,                    
			output   [width-1:0]    x1077_out,                    
			output   [width-1:0]    x1078_out,                    
			output   [width-1:0]    x1079_out,                    
			output   [width-1:0]    x1080_out,                    
			output   [width-1:0]    x1081_out,                    
			output   [width-1:0]    x1082_out,                    
			output   [width-1:0]    x1083_out,                    
			output   [width-1:0]    x1084_out,                    
			output   [width-1:0]    x1085_out,                    
			output   [width-1:0]    x1086_out,                    
			output   [width-1:0]    x1087_out,                    
			output   [width-1:0]    x1088_out,                    
			output   [width-1:0]    x1089_out,                    
			output   [width-1:0]    x1090_out,                    
			output   [width-1:0]    x1091_out,                    
			output   [width-1:0]    x1092_out,                    
			output   [width-1:0]    x1093_out,                    
			output   [width-1:0]    x1094_out,                    
			output   [width-1:0]    x1095_out,                    
			output   [width-1:0]    x1096_out,                    
			output   [width-1:0]    x1097_out,                    
			output   [width-1:0]    x1098_out,                    
			output   [width-1:0]    x1099_out,                    
			output   [width-1:0]    x1100_out,                    
			output   [width-1:0]    x1101_out,                    
			output   [width-1:0]    x1102_out,                    
			output   [width-1:0]    x1103_out,                    
			output   [width-1:0]    x1104_out,                    
			output   [width-1:0]    x1105_out,                    
			output   [width-1:0]    x1106_out,                    
			output   [width-1:0]    x1107_out,                    
			output   [width-1:0]    x1108_out,                    
			output   [width-1:0]    x1109_out,                    
			output   [width-1:0]    x1110_out,                    
			output   [width-1:0]    x1111_out,                    
			output   [width-1:0]    x1112_out,                    
			output   [width-1:0]    x1113_out,                    
			output   [width-1:0]    x1114_out,                    
			output   [width-1:0]    x1115_out,                    
			output   [width-1:0]    x1116_out,                    
			output   [width-1:0]    x1117_out,                    
			output   [width-1:0]    x1118_out,                    
			output   [width-1:0]    x1119_out,                    
			output   [width-1:0]    x1120_out,                    
			output   [width-1:0]    x1121_out,                    
			output   [width-1:0]    x1122_out,                    
			output   [width-1:0]    x1123_out,                    
			output   [width-1:0]    x1124_out,                    
			output   [width-1:0]    x1125_out,                    
			output   [width-1:0]    x1126_out,                    
			output   [width-1:0]    x1127_out,                    
			output   [width-1:0]    x1128_out,                    
			output   [width-1:0]    x1129_out,                    
			output   [width-1:0]    x1130_out,                    
			output   [width-1:0]    x1131_out,                    
			output   [width-1:0]    x1132_out,                    
			output   [width-1:0]    x1133_out,                    
			output   [width-1:0]    x1134_out,                    
			output   [width-1:0]    x1135_out,                    
			output   [width-1:0]    x1136_out,                    
			output   [width-1:0]    x1137_out,                    
			output   [width-1:0]    x1138_out,                    
			output   [width-1:0]    x1139_out,                    
			output   [width-1:0]    x1140_out,                    
			output   [width-1:0]    x1141_out,                    
			output   [width-1:0]    x1142_out,                    
			output   [width-1:0]    x1143_out,                    
			output   [width-1:0]    x1144_out,                    
			output   [width-1:0]    x1145_out,                    
			output   [width-1:0]    x1146_out,                    
			output   [width-1:0]    x1147_out,                    
			output   [width-1:0]    x1148_out,                    
			output   [width-1:0]    x1149_out,                    
			output   [width-1:0]    x1150_out,                    
			output   [width-1:0]    x1151_out,                    
			output   [width-1:0]    x1152_out,                    
			output   [width-1:0]    x1153_out,                    
			output   [width-1:0]    x1154_out,                    
			output   [width-1:0]    x1155_out,                    
			output   [width-1:0]    x1156_out,                    
			output   [width-1:0]    x1157_out,                    
			output   [width-1:0]    x1158_out,                    
			output   [width-1:0]    x1159_out,                    
			output   [width-1:0]    x1160_out,                    
			output   [width-1:0]    x1161_out,                    
			output   [width-1:0]    x1162_out,                    
			output   [width-1:0]    x1163_out,                    
			output   [width-1:0]    x1164_out,                    
			output   [width-1:0]    x1165_out,                    
			output   [width-1:0]    x1166_out,                    
			output   [width-1:0]    x1167_out,                    
			output   [width-1:0]    x1168_out,                    
			output   [width-1:0]    x1169_out,                    
			output   [width-1:0]    x1170_out,                    
			output   [width-1:0]    x1171_out,                    
			output   [width-1:0]    x1172_out,                    
			output   [width-1:0]    x1173_out,                    
			output   [width-1:0]    x1174_out,                    
			output   [width-1:0]    x1175_out,                    
			output   [width-1:0]    x1176_out,                    
			output   [width-1:0]    x1177_out,                    
			output   [width-1:0]    x1178_out,                    
			output   [width-1:0]    x1179_out,                    
			output   [width-1:0]    x1180_out,                    
			output   [width-1:0]    x1181_out,                    
			output   [width-1:0]    x1182_out,                    
			output   [width-1:0]    x1183_out,                    
			output   [width-1:0]    x1184_out,                    
			output   [width-1:0]    x1185_out,                    
			output   [width-1:0]    x1186_out,                    
			output   [width-1:0]    x1187_out,                    
			output   [width-1:0]    x1188_out,                    
			output   [width-1:0]    x1189_out,                    
			output   [width-1:0]    x1190_out,                    
			output   [width-1:0]    x1191_out,                    
			output   [width-1:0]    x1192_out,                    
			output   [width-1:0]    x1193_out,                    
			output   [width-1:0]    x1194_out,                    
			output   [width-1:0]    x1195_out,                    
			output   [width-1:0]    x1196_out,                    
			output   [width-1:0]    x1197_out,                    
			output   [width-1:0]    x1198_out,                    
			output   [width-1:0]    x1199_out,                    
			output   [width-1:0]    x1200_out,                    
			output   [width-1:0]    x1201_out,                    
			output   [width-1:0]    x1202_out,                    
			output   [width-1:0]    x1203_out,                    
			output   [width-1:0]    x1204_out,                    
			output   [width-1:0]    x1205_out,                    
			output   [width-1:0]    x1206_out,                    
			output   [width-1:0]    x1207_out,                    
			output   [width-1:0]    x1208_out,                    
			output   [width-1:0]    x1209_out,                    
			output   [width-1:0]    x1210_out,                    
			output   [width-1:0]    x1211_out,                    
			output   [width-1:0]    x1212_out,                    
			output   [width-1:0]    x1213_out,                    
			output   [width-1:0]    x1214_out,                    
			output   [width-1:0]    x1215_out,                    
			output   [width-1:0]    x1216_out,                    
			output   [width-1:0]    x1217_out,                    
			output   [width-1:0]    x1218_out,                    
			output   [width-1:0]    x1219_out,                    
			output   [width-1:0]    x1220_out,                    
			output   [width-1:0]    x1221_out,                    
			output   [width-1:0]    x1222_out,                    
			output   [width-1:0]    x1223_out,                    
			output   [width-1:0]    x1224_out,                    
			output   [width-1:0]    x1225_out,                    
			output   [width-1:0]    x1226_out,                    
			output   [width-1:0]    x1227_out,                    
			output   [width-1:0]    x1228_out,                    
			output   [width-1:0]    x1229_out,                    
			output   [width-1:0]    x1230_out,                    
			output   [width-1:0]    x1231_out,                    
			output   [width-1:0]    x1232_out,                    
			output   [width-1:0]    x1233_out,                    
			output   [width-1:0]    x1234_out,                    
			output   [width-1:0]    x1235_out,                    
			output   [width-1:0]    x1236_out,                    
			output   [width-1:0]    x1237_out,                    
			output   [width-1:0]    x1238_out,                    
			output   [width-1:0]    x1239_out,                    
			output   [width-1:0]    x1240_out,                    
			output   [width-1:0]    x1241_out,                    
			output   [width-1:0]    x1242_out,                    
			output   [width-1:0]    x1243_out,                    
			output   [width-1:0]    x1244_out,                    
			output   [width-1:0]    x1245_out,                    
			output   [width-1:0]    x1246_out,                    
			output   [width-1:0]    x1247_out,                    
			output   [width-1:0]    x1248_out,                    
			output   [width-1:0]    x1249_out,                    
			output   [width-1:0]    x1250_out,                    
			output   [width-1:0]    x1251_out,                    
			output   [width-1:0]    x1252_out,                    
			output   [width-1:0]    x1253_out,                    
			output   [width-1:0]    x1254_out,                    
			output   [width-1:0]    x1255_out,                    
			output   [width-1:0]    x1256_out,                    
			output   [width-1:0]    x1257_out,                    
			output   [width-1:0]    x1258_out,                    
			output   [width-1:0]    x1259_out,                    
			output   [width-1:0]    x1260_out,                    
			output   [width-1:0]    x1261_out,                    
			output   [width-1:0]    x1262_out,                    
			output   [width-1:0]    x1263_out,                    
			output   [width-1:0]    x1264_out,                    
			output   [width-1:0]    x1265_out,                    
			output   [width-1:0]    x1266_out,                    
			output   [width-1:0]    x1267_out,                    
			output   [width-1:0]    x1268_out,                    
			output   [width-1:0]    x1269_out,                    
			output   [width-1:0]    x1270_out,                    
			output   [width-1:0]    x1271_out,                    
			output   [width-1:0]    x1272_out,                    
			output   [width-1:0]    x1273_out,                    
			output   [width-1:0]    x1274_out,                    
			output   [width-1:0]    x1275_out,                    
			output   [width-1:0]    x1276_out,                    
			output   [width-1:0]    x1277_out,                    
			output   [width-1:0]    x1278_out,                    
			output   [width-1:0]    x1279_out,                    
			output   [width-1:0]    x1280_out,                    
			output   [width-1:0]    x1281_out,                    
			output   [width-1:0]    x1282_out,                    
			output   [width-1:0]    x1283_out,                    
			output   [width-1:0]    x1284_out,                    
			output   [width-1:0]    x1285_out,                    
			output   [width-1:0]    x1286_out,                    
			output   [width-1:0]    x1287_out,                    
			output   [width-1:0]    x1288_out,                    
			output   [width-1:0]    x1289_out,                    
			output   [width-1:0]    x1290_out,                    
			output   [width-1:0]    x1291_out,                    
			output   [width-1:0]    x1292_out,                    
			output   [width-1:0]    x1293_out,                    
			output   [width-1:0]    x1294_out,                    
			output   [width-1:0]    x1295_out,                    
			output   [width-1:0]    x1296_out,                    
			output   [width-1:0]    x1297_out,                    
			output   [width-1:0]    x1298_out,                    
			output   [width-1:0]    x1299_out,                    
			output   [width-1:0]    x1300_out,                    
			output   [width-1:0]    x1301_out,                    
			output   [width-1:0]    x1302_out,                    
			output   [width-1:0]    x1303_out,                    
			output   [width-1:0]    x1304_out,                    
			output   [width-1:0]    x1305_out,                    
			output   [width-1:0]    x1306_out,                    
			output   [width-1:0]    x1307_out,                    
			output   [width-1:0]    x1308_out,                    
			output   [width-1:0]    x1309_out,                    
			output   [width-1:0]    x1310_out,                    
			output   [width-1:0]    x1311_out,                    
			output   [width-1:0]    x1312_out,                    
			output   [width-1:0]    x1313_out,                    
			output   [width-1:0]    x1314_out,                    
			output   [width-1:0]    x1315_out,                    
			output   [width-1:0]    x1316_out,                    
			output   [width-1:0]    x1317_out,                    
			output   [width-1:0]    x1318_out,                    
			output   [width-1:0]    x1319_out,                    
			output   [width-1:0]    x1320_out,                    
			output   [width-1:0]    x1321_out,                    
			output   [width-1:0]    x1322_out,                    
			output   [width-1:0]    x1323_out,                    
			output   [width-1:0]    x1324_out,                    
			output   [width-1:0]    x1325_out,                    
			output   [width-1:0]    x1326_out,                    
			output   [width-1:0]    x1327_out,                    
			output   [width-1:0]    x1328_out,                    
			output   [width-1:0]    x1329_out,                    
			output   [width-1:0]    x1330_out,                    
			output   [width-1:0]    x1331_out,                    
			output   [width-1:0]    x1332_out,                    
			output   [width-1:0]    x1333_out,                    
			output   [width-1:0]    x1334_out,                    
			output   [width-1:0]    x1335_out,                    
			output   [width-1:0]    x1336_out,                    
			output   [width-1:0]    x1337_out,                    
			output   [width-1:0]    x1338_out,                    
			output   [width-1:0]    x1339_out,                    
			output   [width-1:0]    x1340_out,                    
			output   [width-1:0]    x1341_out,                    
			output   [width-1:0]    x1342_out,                    
			output   [width-1:0]    x1343_out,                    
			output   [width-1:0]    x1344_out,                    
			output   [width-1:0]    x1345_out,                    
			output   [width-1:0]    x1346_out,                    
			output   [width-1:0]    x1347_out,                    
			output   [width-1:0]    x1348_out,                    
			output   [width-1:0]    x1349_out,                    
			output   [width-1:0]    x1350_out,                    
			output   [width-1:0]    x1351_out,                    
			output   [width-1:0]    x1352_out,                    
			output   [width-1:0]    x1353_out,                    
			output   [width-1:0]    x1354_out,                    
			output   [width-1:0]    x1355_out,                    
			output   [width-1:0]    x1356_out,                    
			output   [width-1:0]    x1357_out,                    
			output   [width-1:0]    x1358_out,                    
			output   [width-1:0]    x1359_out,                    
			output   [width-1:0]    x1360_out,                    
			output   [width-1:0]    x1361_out,                    
			output   [width-1:0]    x1362_out,                    
			output   [width-1:0]    x1363_out,                    
			output   [width-1:0]    x1364_out,                    
			output   [width-1:0]    x1365_out,                    
			output   [width-1:0]    x1366_out,                    
			output   [width-1:0]    x1367_out,                    
			output   [width-1:0]    x1368_out,                    
			output   [width-1:0]    x1369_out,                    
			output   [width-1:0]    x1370_out,                    
			output   [width-1:0]    x1371_out,                    
			output   [width-1:0]    x1372_out,                    
			output   [width-1:0]    x1373_out,                    
			output   [width-1:0]    x1374_out,                    
			output   [width-1:0]    x1375_out,                    
			output   [width-1:0]    x1376_out,                    
			output   [width-1:0]    x1377_out,                    
			output   [width-1:0]    x1378_out,                    
			output   [width-1:0]    x1379_out,                    
			output   [width-1:0]    x1380_out,                    
			output   [width-1:0]    x1381_out,                    
			output   [width-1:0]    x1382_out,                    
			output   [width-1:0]    x1383_out,                    
			output   [width-1:0]    x1384_out,                    
			output   [width-1:0]    x1385_out,                    
			output   [width-1:0]    x1386_out,                    
			output   [width-1:0]    x1387_out,                    
			output   [width-1:0]    x1388_out,                    
			output   [width-1:0]    x1389_out,                    
			output   [width-1:0]    x1390_out,                    
			output   [width-1:0]    x1391_out,                    
			output   [width-1:0]    x1392_out,                    
			output   [width-1:0]    x1393_out,                    
			output   [width-1:0]    x1394_out,                    
			output   [width-1:0]    x1395_out,                    
			output   [width-1:0]    x1396_out,                    
			output   [width-1:0]    x1397_out,                    
			output   [width-1:0]    x1398_out,                    
			output   [width-1:0]    x1399_out,                    
			output   [width-1:0]    x1400_out,                    
			output   [width-1:0]    x1401_out,                    
			output   [width-1:0]    x1402_out,                    
			output   [width-1:0]    x1403_out,                    
			output   [width-1:0]    x1404_out,                    
			output   [width-1:0]    x1405_out,                    
			output   [width-1:0]    x1406_out,                    
			output   [width-1:0]    x1407_out,                    
			output   [width-1:0]    x1408_out,                    
			output   [width-1:0]    x1409_out,                    
			output   [width-1:0]    x1410_out,                    
			output   [width-1:0]    x1411_out,                    
			output   [width-1:0]    x1412_out,                    
			output   [width-1:0]    x1413_out,                    
			output   [width-1:0]    x1414_out,                    
			output   [width-1:0]    x1415_out,                    
			output   [width-1:0]    x1416_out,                    
			output   [width-1:0]    x1417_out,                    
			output   [width-1:0]    x1418_out,                    
			output   [width-1:0]    x1419_out,                    
			output   [width-1:0]    x1420_out,                    
			output   [width-1:0]    x1421_out,                    
			output   [width-1:0]    x1422_out,                    
			output   [width-1:0]    x1423_out,                    
			output   [width-1:0]    x1424_out,                    
			output   [width-1:0]    x1425_out,                    
			output   [width-1:0]    x1426_out,                    
			output   [width-1:0]    x1427_out,                    
			output   [width-1:0]    x1428_out,                    
			output   [width-1:0]    x1429_out,                    
			output   [width-1:0]    x1430_out,                    
			output   [width-1:0]    x1431_out,                    
			output   [width-1:0]    x1432_out,                    
			output   [width-1:0]    x1433_out,                    
			output   [width-1:0]    x1434_out,                    
			output   [width-1:0]    x1435_out,                    
			output   [width-1:0]    x1436_out,                    
			output   [width-1:0]    x1437_out,                    
			output   [width-1:0]    x1438_out,                    
			output   [width-1:0]    x1439_out,                    
			output   [width-1:0]    x1440_out,                    
			output   [width-1:0]    x1441_out,                    
			output   [width-1:0]    x1442_out,                    
			output   [width-1:0]    x1443_out,                    
			output   [width-1:0]    x1444_out,                    
			output   [width-1:0]    x1445_out,                    
			output   [width-1:0]    x1446_out,                    
			output   [width-1:0]    x1447_out,                    
			output   [width-1:0]    x1448_out,                    
			output   [width-1:0]    x1449_out,                    
			output   [width-1:0]    x1450_out,                    
			output   [width-1:0]    x1451_out,                    
			output   [width-1:0]    x1452_out,                    
			output   [width-1:0]    x1453_out,                    
			output   [width-1:0]    x1454_out,                    
			output   [width-1:0]    x1455_out,                    
			output   [width-1:0]    x1456_out,                    
			output   [width-1:0]    x1457_out,                    
			output   [width-1:0]    x1458_out,                    
			output   [width-1:0]    x1459_out,                    
			output   [width-1:0]    x1460_out,                    
			output   [width-1:0]    x1461_out,                    
			output   [width-1:0]    x1462_out,                    
			output   [width-1:0]    x1463_out,                    
			output   [width-1:0]    x1464_out,                    
			output   [width-1:0]    x1465_out,                    
			output   [width-1:0]    x1466_out,                    
			output   [width-1:0]    x1467_out,                    
			output   [width-1:0]    x1468_out,                    
			output   [width-1:0]    x1469_out,                    
			output   [width-1:0]    x1470_out,                    
			output   [width-1:0]    x1471_out,                    
			output   [width-1:0]    x1472_out,                    
			output   [width-1:0]    x1473_out,                    
			output   [width-1:0]    x1474_out,                    
			output   [width-1:0]    x1475_out,                    
			output   [width-1:0]    x1476_out,                    
			output   [width-1:0]    x1477_out,                    
			output   [width-1:0]    x1478_out,                    
			output   [width-1:0]    x1479_out,                    
			output   [width-1:0]    x1480_out,                    
			output   [width-1:0]    x1481_out,                    
			output   [width-1:0]    x1482_out,                    
			output   [width-1:0]    x1483_out,                    
			output   [width-1:0]    x1484_out,                    
			output   [width-1:0]    x1485_out,                    
			output   [width-1:0]    x1486_out,                    
			output   [width-1:0]    x1487_out,                    
			output   [width-1:0]    x1488_out,                    
			output   [width-1:0]    x1489_out,                    
			output   [width-1:0]    x1490_out,                    
			output   [width-1:0]    x1491_out,                    
			output   [width-1:0]    x1492_out,                    
			output   [width-1:0]    x1493_out,                    
			output   [width-1:0]    x1494_out,                    
			output   [width-1:0]    x1495_out,                    
			output   [width-1:0]    x1496_out,                    
			output   [width-1:0]    x1497_out,                    
			output   [width-1:0]    x1498_out,                    
			output   [width-1:0]    x1499_out,                    
			output   [width-1:0]    x1500_out,                    
			output   [width-1:0]    x1501_out,                    
			output   [width-1:0]    x1502_out,                    
			output   [width-1:0]    x1503_out,                    
			output   [width-1:0]    x1504_out,                    
			output   [width-1:0]    x1505_out,                    
			output   [width-1:0]    x1506_out,                    
			output   [width-1:0]    x1507_out,                    
			output   [width-1:0]    x1508_out,                    
			output   [width-1:0]    x1509_out,                    
			output   [width-1:0]    x1510_out,                    
			output   [width-1:0]    x1511_out,                    
			output   [width-1:0]    x1512_out,                    
			output   [width-1:0]    x1513_out,                    
			output   [width-1:0]    x1514_out,                    
			output   [width-1:0]    x1515_out,                    
			output   [width-1:0]    x1516_out,                    
			output   [width-1:0]    x1517_out,                    
			output   [width-1:0]    x1518_out,                    
			output   [width-1:0]    x1519_out,                    
			output   [width-1:0]    x1520_out,                    
			output   [width-1:0]    x1521_out,                    
			output   [width-1:0]    x1522_out,                    
			output   [width-1:0]    x1523_out,                    
			output   [width-1:0]    x1524_out,                    
			output   [width-1:0]    x1525_out,                    
			output   [width-1:0]    x1526_out,                    
			output   [width-1:0]    x1527_out,                    
			output   [width-1:0]    x1528_out,                    
			output   [width-1:0]    x1529_out,                    
			output   [width-1:0]    x1530_out,                    
			output   [width-1:0]    x1531_out,                    
			output   [width-1:0]    x1532_out,                    
			output   [width-1:0]    x1533_out,                    
			output   [width-1:0]    x1534_out,                    
			output   [width-1:0]    x1535_out,                    
			output   [width-1:0]    x1536_out,                    
			output   [width-1:0]    x1537_out,                    
			output   [width-1:0]    x1538_out,                    
			output   [width-1:0]    x1539_out,                    
			output   [width-1:0]    x1540_out,                    
			output   [width-1:0]    x1541_out,                    
			output   [width-1:0]    x1542_out,                    
			output   [width-1:0]    x1543_out,                    
			output   [width-1:0]    x1544_out,                    
			output   [width-1:0]    x1545_out,                    
			output   [width-1:0]    x1546_out,                    
			output   [width-1:0]    x1547_out,                    
			output   [width-1:0]    x1548_out,                    
			output   [width-1:0]    x1549_out,                    
			output   [width-1:0]    x1550_out,                    
			output   [width-1:0]    x1551_out,                    
			output   [width-1:0]    x1552_out,                    
			output   [width-1:0]    x1553_out,                    
			output   [width-1:0]    x1554_out,                    
			output   [width-1:0]    x1555_out,                    
			output   [width-1:0]    x1556_out,                    
			output   [width-1:0]    x1557_out,                    
			output   [width-1:0]    x1558_out,                    
			output   [width-1:0]    x1559_out,                    
			output   [width-1:0]    x1560_out,                    
			output   [width-1:0]    x1561_out,                    
			output   [width-1:0]    x1562_out,                    
			output   [width-1:0]    x1563_out,                    
			output   [width-1:0]    x1564_out,                    
			output   [width-1:0]    x1565_out,                    
			output   [width-1:0]    x1566_out,                    
			output   [width-1:0]    x1567_out,                    
			output   [width-1:0]    x1568_out,                    
			output   [width-1:0]    x1569_out,                    
			output   [width-1:0]    x1570_out,                    
			output   [width-1:0]    x1571_out,                    
			output   [width-1:0]    x1572_out,                    
			output   [width-1:0]    x1573_out,                    
			output   [width-1:0]    x1574_out,                    
			output   [width-1:0]    x1575_out,                    
			output   [width-1:0]    x1576_out,                    
			output   [width-1:0]    x1577_out,                    
			output   [width-1:0]    x1578_out,                    
			output   [width-1:0]    x1579_out,                    
			output   [width-1:0]    x1580_out,                    
			output   [width-1:0]    x1581_out,                    
			output   [width-1:0]    x1582_out,                    
			output   [width-1:0]    x1583_out,                    
			output   [width-1:0]    x1584_out,                    
			output   [width-1:0]    x1585_out,                    
			output   [width-1:0]    x1586_out,                    
			output   [width-1:0]    x1587_out,                    
			output   [width-1:0]    x1588_out,                    
			output   [width-1:0]    x1589_out,                    
			output   [width-1:0]    x1590_out,                    
			output   [width-1:0]    x1591_out,                    
			output   [width-1:0]    x1592_out,                    
			output   [width-1:0]    x1593_out,                    
			output   [width-1:0]    x1594_out,                    
			output   [width-1:0]    x1595_out,                    
			output   [width-1:0]    x1596_out,                    
			output   [width-1:0]    x1597_out,                    
			output   [width-1:0]    x1598_out,                    
			output   [width-1:0]    x1599_out,                    
			output   [width-1:0]    x1600_out,                    
			output   [width-1:0]    x1601_out,                    
			output   [width-1:0]    x1602_out,                    
			output   [width-1:0]    x1603_out,                    
			output   [width-1:0]    x1604_out,                    
			output   [width-1:0]    x1605_out,                    
			output   [width-1:0]    x1606_out,                    
			output   [width-1:0]    x1607_out,                    
			output   [width-1:0]    x1608_out,                    
			output   [width-1:0]    x1609_out,                    
			output   [width-1:0]    x1610_out,                    
			output   [width-1:0]    x1611_out,                    
			output   [width-1:0]    x1612_out,                    
			output   [width-1:0]    x1613_out,                    
			output   [width-1:0]    x1614_out,                    
			output   [width-1:0]    x1615_out,                    
			output   [width-1:0]    x1616_out,                    
			output   [width-1:0]    x1617_out,                    
			output   [width-1:0]    x1618_out,                    
			output   [width-1:0]    x1619_out,                    
			output   [width-1:0]    x1620_out,                    
			output   [width-1:0]    x1621_out,                    
			output   [width-1:0]    x1622_out,                    
			output   [width-1:0]    x1623_out,                    
			output   [width-1:0]    x1624_out,                    
			output   [width-1:0]    x1625_out,                    
			output   [width-1:0]    x1626_out,                    
			output   [width-1:0]    x1627_out,                    
			output   [width-1:0]    x1628_out,                    
			output   [width-1:0]    x1629_out,                    
			output   [width-1:0]    x1630_out,                    
			output   [width-1:0]    x1631_out,                    
			output   [width-1:0]    x1632_out,                    
			output   [width-1:0]    x1633_out,                    
			output   [width-1:0]    x1634_out,                    
			output   [width-1:0]    x1635_out,                    
			output   [width-1:0]    x1636_out,                    
			output   [width-1:0]    x1637_out,                    
			output   [width-1:0]    x1638_out,                    
			output   [width-1:0]    x1639_out,                    
			output   [width-1:0]    x1640_out,                    
			output   [width-1:0]    x1641_out,                    
			output   [width-1:0]    x1642_out,                    
			output   [width-1:0]    x1643_out,                    
			output   [width-1:0]    x1644_out,                    
			output   [width-1:0]    x1645_out,                    
			output   [width-1:0]    x1646_out,                    
			output   [width-1:0]    x1647_out,                    
			output   [width-1:0]    x1648_out,                    
			output   [width-1:0]    x1649_out,                    
			output   [width-1:0]    x1650_out,                    
			output   [width-1:0]    x1651_out,                    
			output   [width-1:0]    x1652_out,                    
			output   [width-1:0]    x1653_out,                    
			output   [width-1:0]    x1654_out,                    
			output   [width-1:0]    x1655_out,                    
			output   [width-1:0]    x1656_out,                    
			output   [width-1:0]    x1657_out,                    
			output   [width-1:0]    x1658_out,                    
			output   [width-1:0]    x1659_out,                    
			output   [width-1:0]    x1660_out,                    
			output   [width-1:0]    x1661_out,                    
			output   [width-1:0]    x1662_out,                    
			output   [width-1:0]    x1663_out,                    
			output   [width-1:0]    x1664_out,                    
			output   [width-1:0]    x1665_out,                    
			output   [width-1:0]    x1666_out,                    
			output   [width-1:0]    x1667_out,                    
			output   [width-1:0]    x1668_out,                    
			output   [width-1:0]    x1669_out,                    
			output   [width-1:0]    x1670_out,                    
			output   [width-1:0]    x1671_out,                    
			output   [width-1:0]    x1672_out,                    
			output   [width-1:0]    x1673_out,                    
			output   [width-1:0]    x1674_out,                    
			output   [width-1:0]    x1675_out,                    
			output   [width-1:0]    x1676_out,                    
			output   [width-1:0]    x1677_out,                    
			output   [width-1:0]    x1678_out,                    
			output   [width-1:0]    x1679_out,                    
			output   [width-1:0]    x1680_out,                    
			output   [width-1:0]    x1681_out,                    
			output   [width-1:0]    x1682_out,                    
			output   [width-1:0]    x1683_out,                    
			output   [width-1:0]    x1684_out,                    
			output   [width-1:0]    x1685_out,                    
			output   [width-1:0]    x1686_out,                    
			output   [width-1:0]    x1687_out,                    
			output   [width-1:0]    x1688_out,                    
			output   [width-1:0]    x1689_out,                    
			output   [width-1:0]    x1690_out,                    
			output   [width-1:0]    x1691_out,                    
			output   [width-1:0]    x1692_out,                    
			output   [width-1:0]    x1693_out,                    
			output   [width-1:0]    x1694_out,                    
			output   [width-1:0]    x1695_out,                    
			output   [width-1:0]    x1696_out,                    
			output   [width-1:0]    x1697_out,                    
			output   [width-1:0]    x1698_out,                    
			output   [width-1:0]    x1699_out,                    
			output   [width-1:0]    x1700_out,                    
			output   [width-1:0]    x1701_out,                    
			output   [width-1:0]    x1702_out,                    
			output   [width-1:0]    x1703_out,                    
			output   [width-1:0]    x1704_out,                    
			output   [width-1:0]    x1705_out,                    
			output   [width-1:0]    x1706_out,                    
			output   [width-1:0]    x1707_out,                    
			output   [width-1:0]    x1708_out,                    
			output   [width-1:0]    x1709_out,                    
			output   [width-1:0]    x1710_out,                    
			output   [width-1:0]    x1711_out,                    
			output   [width-1:0]    x1712_out,                    
			output   [width-1:0]    x1713_out,                    
			output   [width-1:0]    x1714_out,                    
			output   [width-1:0]    x1715_out,                    
			output   [width-1:0]    x1716_out,                    
			output   [width-1:0]    x1717_out,                    
			output   [width-1:0]    x1718_out,                    
			output   [width-1:0]    x1719_out,                    
			output   [width-1:0]    x1720_out,                    
			output   [width-1:0]    x1721_out,                    
			output   [width-1:0]    x1722_out,                    
			output   [width-1:0]    x1723_out,                    
			output   [width-1:0]    x1724_out,                    
			output   [width-1:0]    x1725_out,                    
			output   [width-1:0]    x1726_out,                    
			output   [width-1:0]    x1727_out,                    
			output   [width-1:0]    x1728_out,                    
			output   [width-1:0]    x1729_out,                    
			output   [width-1:0]    x1730_out,                    
			output   [width-1:0]    x1731_out,                    
			output   [width-1:0]    x1732_out,                    
			output   [width-1:0]    x1733_out,                    
			output   [width-1:0]    x1734_out,                    
			output   [width-1:0]    x1735_out,                    
			output   [width-1:0]    x1736_out,                    
			output   [width-1:0]    x1737_out,                    
			output   [width-1:0]    x1738_out,                    
			output   [width-1:0]    x1739_out,                    
			output   [width-1:0]    x1740_out,                    
			output   [width-1:0]    x1741_out,                    
			output   [width-1:0]    x1742_out,                    
			output   [width-1:0]    x1743_out,                    
			output   [width-1:0]    x1744_out,                    
			output   [width-1:0]    x1745_out,                    
			output   [width-1:0]    x1746_out,                    
			output   [width-1:0]    x1747_out,                    
			output   [width-1:0]    x1748_out,                    
			output   [width-1:0]    x1749_out,                    
			output   [width-1:0]    x1750_out,                    
			output   [width-1:0]    x1751_out,                    
			output   [width-1:0]    x1752_out,                    
			output   [width-1:0]    x1753_out,                    
			output   [width-1:0]    x1754_out,                    
			output   [width-1:0]    x1755_out,                    
			output   [width-1:0]    x1756_out,                    
			output   [width-1:0]    x1757_out,                    
			output   [width-1:0]    x1758_out,                    
			output   [width-1:0]    x1759_out,                    
			output   [width-1:0]    x1760_out,                    
			output   [width-1:0]    x1761_out,                    
			output   [width-1:0]    x1762_out,                    
			output   [width-1:0]    x1763_out,                    
			output   [width-1:0]    x1764_out,                    
			output   [width-1:0]    x1765_out,                    
			output   [width-1:0]    x1766_out,                    
			output   [width-1:0]    x1767_out,                    
			output   [width-1:0]    x1768_out,                    
			output   [width-1:0]    x1769_out,                    
			output   [width-1:0]    x1770_out,                    
			output   [width-1:0]    x1771_out,                    
			output   [width-1:0]    x1772_out,                    
			output   [width-1:0]    x1773_out,                    
			output   [width-1:0]    x1774_out,                    
			output   [width-1:0]    x1775_out,                    
			output   [width-1:0]    x1776_out,                    
			output   [width-1:0]    x1777_out,                    
			output   [width-1:0]    x1778_out,                    
			output   [width-1:0]    x1779_out,                    
			output   [width-1:0]    x1780_out,                    
			output   [width-1:0]    x1781_out,                    
			output   [width-1:0]    x1782_out,                    
			output   [width-1:0]    x1783_out,                    
			output   [width-1:0]    x1784_out,                    
			output   [width-1:0]    x1785_out,                    
			output   [width-1:0]    x1786_out,                    
			output   [width-1:0]    x1787_out,                    
			output   [width-1:0]    x1788_out,                    
			output   [width-1:0]    x1789_out,                    
			output   [width-1:0]    x1790_out,                    
			output   [width-1:0]    x1791_out,                    
			output   [width-1:0]    x1792_out,                    
			output   [width-1:0]    x1793_out,                    
			output   [width-1:0]    x1794_out,                    
			output   [width-1:0]    x1795_out,                    
			output   [width-1:0]    x1796_out,                    
			output   [width-1:0]    x1797_out,                    
			output   [width-1:0]    x1798_out,                    
			output   [width-1:0]    x1799_out,                    
			output   [width-1:0]    x1800_out,                    
			output   [width-1:0]    x1801_out,                    
			output   [width-1:0]    x1802_out,                    
			output   [width-1:0]    x1803_out,                    
			output   [width-1:0]    x1804_out,                    
			output   [width-1:0]    x1805_out,                    
			output   [width-1:0]    x1806_out,                    
			output   [width-1:0]    x1807_out,                    
			output   [width-1:0]    x1808_out,                    
			output   [width-1:0]    x1809_out,                    
			output   [width-1:0]    x1810_out,                    
			output   [width-1:0]    x1811_out,                    
			output   [width-1:0]    x1812_out,                    
			output   [width-1:0]    x1813_out,                    
			output   [width-1:0]    x1814_out,                    
			output   [width-1:0]    x1815_out,                    
			output   [width-1:0]    x1816_out,                    
			output   [width-1:0]    x1817_out,                    
			output   [width-1:0]    x1818_out,                    
			output   [width-1:0]    x1819_out,                    
			output   [width-1:0]    x1820_out,                    
			output   [width-1:0]    x1821_out,                    
			output   [width-1:0]    x1822_out,                    
			output   [width-1:0]    x1823_out,                    
			output   [width-1:0]    x1824_out,                    
			output   [width-1:0]    x1825_out,                    
			output   [width-1:0]    x1826_out,                    
			output   [width-1:0]    x1827_out,                    
			output   [width-1:0]    x1828_out,                    
			output   [width-1:0]    x1829_out,                    
			output   [width-1:0]    x1830_out,                    
			output   [width-1:0]    x1831_out,                    
			output   [width-1:0]    x1832_out,                    
			output   [width-1:0]    x1833_out,                    
			output   [width-1:0]    x1834_out,                    
			output   [width-1:0]    x1835_out,                    
			output   [width-1:0]    x1836_out,                    
			output   [width-1:0]    x1837_out,                    
			output   [width-1:0]    x1838_out,                    
			output   [width-1:0]    x1839_out,                    
			output   [width-1:0]    x1840_out,                    
			output   [width-1:0]    x1841_out,                    
			output   [width-1:0]    x1842_out,                    
			output   [width-1:0]    x1843_out,                    
			output   [width-1:0]    x1844_out,                    
			output   [width-1:0]    x1845_out,                    
			output   [width-1:0]    x1846_out,                    
			output   [width-1:0]    x1847_out,                    
			output   [width-1:0]    x1848_out,                    
			output   [width-1:0]    x1849_out,                    
			output   [width-1:0]    x1850_out,                    
			output   [width-1:0]    x1851_out,                    
			output   [width-1:0]    x1852_out,                    
			output   [width-1:0]    x1853_out,                    
			output   [width-1:0]    x1854_out,                    
			output   [width-1:0]    x1855_out,                    
			output   [width-1:0]    x1856_out,                    
			output   [width-1:0]    x1857_out,                    
			output   [width-1:0]    x1858_out,                    
			output   [width-1:0]    x1859_out,                    
			output   [width-1:0]    x1860_out,                    
			output   [width-1:0]    x1861_out,                    
			output   [width-1:0]    x1862_out,                    
			output   [width-1:0]    x1863_out,                    
			output   [width-1:0]    x1864_out,                    
			output   [width-1:0]    x1865_out,                    
			output   [width-1:0]    x1866_out,                    
			output   [width-1:0]    x1867_out,                    
			output   [width-1:0]    x1868_out,                    
			output   [width-1:0]    x1869_out,                    
			output   [width-1:0]    x1870_out,                    
			output   [width-1:0]    x1871_out,                    
			output   [width-1:0]    x1872_out,                    
			output   [width-1:0]    x1873_out,                    
			output   [width-1:0]    x1874_out,                    
			output   [width-1:0]    x1875_out,                    
			output   [width-1:0]    x1876_out,                    
			output   [width-1:0]    x1877_out,                    
			output   [width-1:0]    x1878_out,                    
			output   [width-1:0]    x1879_out,                    
			output   [width-1:0]    x1880_out,                    
			output   [width-1:0]    x1881_out,                    
			output   [width-1:0]    x1882_out,                    
			output   [width-1:0]    x1883_out,                    
			output   [width-1:0]    x1884_out,                    
			output   [width-1:0]    x1885_out,                    
			output   [width-1:0]    x1886_out,                    
			output   [width-1:0]    x1887_out,                    
			output   [width-1:0]    x1888_out,                    
			output   [width-1:0]    x1889_out,                    
			output   [width-1:0]    x1890_out,                    
			output   [width-1:0]    x1891_out,                    
			output   [width-1:0]    x1892_out,                    
			output   [width-1:0]    x1893_out,                    
			output   [width-1:0]    x1894_out,                    
			output   [width-1:0]    x1895_out,                    
			output   [width-1:0]    x1896_out,                    
			output   [width-1:0]    x1897_out,                    
			output   [width-1:0]    x1898_out,                    
			output   [width-1:0]    x1899_out,                    
			output   [width-1:0]    x1900_out,                    
			output   [width-1:0]    x1901_out,                    
			output   [width-1:0]    x1902_out,                    
			output   [width-1:0]    x1903_out,                    
			output   [width-1:0]    x1904_out,                    
			output   [width-1:0]    x1905_out,                    
			output   [width-1:0]    x1906_out,                    
			output   [width-1:0]    x1907_out,                    
			output   [width-1:0]    x1908_out,                    
			output   [width-1:0]    x1909_out,                    
			output   [width-1:0]    x1910_out,                    
			output   [width-1:0]    x1911_out,                    
			output   [width-1:0]    x1912_out,                    
			output   [width-1:0]    x1913_out,                    
			output   [width-1:0]    x1914_out,                    
			output   [width-1:0]    x1915_out,                    
			output   [width-1:0]    x1916_out,                    
			output   [width-1:0]    x1917_out,                    
			output   [width-1:0]    x1918_out,                    
			output   [width-1:0]    x1919_out,                    
			output   [width-1:0]    x1920_out,                    
			output   [width-1:0]    x1921_out,                    
			output   [width-1:0]    x1922_out,                    
			output   [width-1:0]    x1923_out,                    
			output   [width-1:0]    x1924_out,                    
			output   [width-1:0]    x1925_out,                    
			output   [width-1:0]    x1926_out,                    
			output   [width-1:0]    x1927_out,                    
			output   [width-1:0]    x1928_out,                    
			output   [width-1:0]    x1929_out,                    
			output   [width-1:0]    x1930_out,                    
			output   [width-1:0]    x1931_out,                    
			output   [width-1:0]    x1932_out,                    
			output   [width-1:0]    x1933_out,                    
			output   [width-1:0]    x1934_out,                    
			output   [width-1:0]    x1935_out,                    
			output   [width-1:0]    x1936_out,                    
			output   [width-1:0]    x1937_out,                    
			output   [width-1:0]    x1938_out,                    
			output   [width-1:0]    x1939_out,                    
			output   [width-1:0]    x1940_out,                    
			output   [width-1:0]    x1941_out,                    
			output   [width-1:0]    x1942_out,                    
			output   [width-1:0]    x1943_out,                    
			output   [width-1:0]    x1944_out,                    
			output   [width-1:0]    x1945_out,                    
			output   [width-1:0]    x1946_out,                    
			output   [width-1:0]    x1947_out,                    
			output   [width-1:0]    x1948_out,                    
			output   [width-1:0]    x1949_out,                    
			output   [width-1:0]    x1950_out,                    
			output   [width-1:0]    x1951_out,                    
			output   [width-1:0]    x1952_out,                    
			output   [width-1:0]    x1953_out,                    
			output   [width-1:0]    x1954_out,                    
			output   [width-1:0]    x1955_out,                    
			output   [width-1:0]    x1956_out,                    
			output   [width-1:0]    x1957_out,                    
			output   [width-1:0]    x1958_out,                    
			output   [width-1:0]    x1959_out,                    
			output   [width-1:0]    x1960_out,                    
			output   [width-1:0]    x1961_out,                    
			output   [width-1:0]    x1962_out,                    
			output   [width-1:0]    x1963_out,                    
			output   [width-1:0]    x1964_out,                    
			output   [width-1:0]    x1965_out,                    
			output   [width-1:0]    x1966_out,                    
			output   [width-1:0]    x1967_out,                    
			output   [width-1:0]    x1968_out,                    
			output   [width-1:0]    x1969_out,                    
			output   [width-1:0]    x1970_out,                    
			output   [width-1:0]    x1971_out,                    
			output   [width-1:0]    x1972_out,                    
			output   [width-1:0]    x1973_out,                    
			output   [width-1:0]    x1974_out,                    
			output   [width-1:0]    x1975_out,                    
			output   [width-1:0]    x1976_out,                    
			output   [width-1:0]    x1977_out,                    
			output   [width-1:0]    x1978_out,                    
			output   [width-1:0]    x1979_out,                    
			output   [width-1:0]    x1980_out,                    
			output   [width-1:0]    x1981_out,                    
			output   [width-1:0]    x1982_out,                    
			output   [width-1:0]    x1983_out,                    
			output   [width-1:0]    x1984_out,                    
			output   [width-1:0]    x1985_out,                    
			output   [width-1:0]    x1986_out,                    
			output   [width-1:0]    x1987_out,                    
			output   [width-1:0]    x1988_out,                    
			output   [width-1:0]    x1989_out,                    
			output   [width-1:0]    x1990_out,                    
			output   [width-1:0]    x1991_out,                    
			output   [width-1:0]    x1992_out,                    
			output   [width-1:0]    x1993_out,                    
			output   [width-1:0]    x1994_out,                    
			output   [width-1:0]    x1995_out,                    
			output   [width-1:0]    x1996_out,                    
			output   [width-1:0]    x1997_out,                    
			output   [width-1:0]    x1998_out,                    
			output   [width-1:0]    x1999_out,                    
			output   [width-1:0]    x2000_out,                    
			output   [width-1:0]    x2001_out,                    
			output   [width-1:0]    x2002_out,                    
			output   [width-1:0]    x2003_out,                    
			output   [width-1:0]    x2004_out,                    
			output   [width-1:0]    x2005_out,                    
			output   [width-1:0]    x2006_out,                    
			output   [width-1:0]    x2007_out,                    
			output   [width-1:0]    x2008_out,                    
			output   [width-1:0]    x2009_out,                    
			output   [width-1:0]    x2010_out,                    
			output   [width-1:0]    x2011_out,                    
			output   [width-1:0]    x2012_out,                    
			output   [width-1:0]    x2013_out,                    
			output   [width-1:0]    x2014_out,                    
			output   [width-1:0]    x2015_out,                    
			output   [width-1:0]    x2016_out,                    
			output   [width-1:0]    x2017_out,                    
			output   [width-1:0]    x2018_out,                    
			output   [width-1:0]    x2019_out,                    
			output   [width-1:0]    x2020_out,                    
			output   [width-1:0]    x2021_out,                    
			output   [width-1:0]    x2022_out,                    
			output   [width-1:0]    x2023_out,                    
			output   [width-1:0]    x2024_out,                    
			output   [width-1:0]    x2025_out,                    
			output   [width-1:0]    x2026_out,                    
			output   [width-1:0]    x2027_out,                    
			output   [width-1:0]    x2028_out,                    
			output   [width-1:0]    x2029_out,                    
			output   [width-1:0]    x2030_out,                    
			output   [width-1:0]    x2031_out,                    
			output   [width-1:0]    x2032_out,                    
			output   [width-1:0]    x2033_out,                    
			output   [width-1:0]    x2034_out,                    
			output   [width-1:0]    x2035_out,                    
			output   [width-1:0]    x2036_out,                    
			output   [width-1:0]    x2037_out,                    
			output   [width-1:0]    x2038_out,                    
			output   [width-1:0]    x2039_out,                    
			output   [width-1:0]    x2040_out,                    
			output   [width-1:0]    x2041_out,                    
			output   [width-1:0]    x2042_out,                    
			output   [width-1:0]    x2043_out,                    
			output   [width-1:0]    x2044_out,                    
			output   [width-1:0]    x2045_out,                    
			output   [width-1:0]    x2046_out,                    
			output   [width-1:0]    x2047_out                     
);

		//--- signal definition
			wire  [width-1:0]        coef[size-1:0];

			reg   [width-1:0]        a0_wr[size-1:0];
			wire  [width-1:0]        a1_wr[size-1:0];
			wire  [width-1:0]        a2_wr[size-1:0];
			wire  [width-1:0]        a3_wr[size-1:0];
			wire  [width-1:0]        a4_wr[size-1:0];
			wire  [width-1:0]        a5_wr[size-1:0];
			wire  [width-1:0]        a6_wr[size-1:0];
			wire  [width-1:0]        a7_wr[size-1:0];
			wire  [width-1:0]        a8_wr[size-1:0];
			wire  [width-1:0]        a9_wr[size-1:0];
			wire  [width-1:0]        a10_wr[size-1:0];
			wire  [width-1:0]        a11_wr[size-1:0];
			wire                     comb_stall;

		//--- cofficient assignment
			assign coef[0] =    {12'b011111111111, 12'b000000000000};
			assign coef[1] =    {12'b011111111111, 12'b111111111010};
			assign coef[2] =    {12'b011111111111, 12'b111111110011};
			assign coef[3] =    {12'b011111111111, 12'b111111101101};
			assign coef[4] =    {12'b011111111111, 12'b111111100111};
			assign coef[5] =    {12'b011111111111, 12'b111111100001};
			assign coef[6] =    {12'b011111111111, 12'b111111011010};
			assign coef[7] =    {12'b011111111111, 12'b111111010100};
			assign coef[8] =    {12'b011111111110, 12'b111111001110};
			assign coef[9] =    {12'b011111111110, 12'b111111000111};
			assign coef[10] =   {12'b011111111110, 12'b111111000001};
			assign coef[11] =   {12'b011111111110, 12'b111110111011};
			assign coef[12] =   {12'b011111111110, 12'b111110110101};
			assign coef[13] =   {12'b011111111101, 12'b111110101110};
			assign coef[14] =   {12'b011111111101, 12'b111110101000};
			assign coef[15] =   {12'b011111111101, 12'b111110100010};
			assign coef[16] =   {12'b011111111101, 12'b111110011100};
			assign coef[17] =   {12'b011111111100, 12'b111110010101};
			assign coef[18] =   {12'b011111111100, 12'b111110001111};
			assign coef[19] =   {12'b011111111100, 12'b111110001001};
			assign coef[20] =   {12'b011111111011, 12'b111110000010};
			assign coef[21] =   {12'b011111111011, 12'b111101111100};
			assign coef[22] =   {12'b011111111010, 12'b111101110110};
			assign coef[23] =   {12'b011111111010, 12'b111101110000};
			assign coef[24] =   {12'b011111111010, 12'b111101101001};
			assign coef[25] =   {12'b011111111001, 12'b111101100011};
			assign coef[26] =   {12'b011111111001, 12'b111101011101};
			assign coef[27] =   {12'b011111111000, 12'b111101010111};
			assign coef[28] =   {12'b011111111000, 12'b111101010000};
			assign coef[29] =   {12'b011111110111, 12'b111101001010};
			assign coef[30] =   {12'b011111110110, 12'b111101000100};
			assign coef[31] =   {12'b011111110110, 12'b111100111110};
			assign coef[32] =   {12'b011111110101, 12'b111100110111};
			assign coef[33] =   {12'b011111110101, 12'b111100110001};
			assign coef[34] =   {12'b011111110100, 12'b111100101011};
			assign coef[35] =   {12'b011111110011, 12'b111100100101};
			assign coef[36] =   {12'b011111110011, 12'b111100011110};
			assign coef[37] =   {12'b011111110010, 12'b111100011000};
			assign coef[38] =   {12'b011111110001, 12'b111100010010};
			assign coef[39] =   {12'b011111110000, 12'b111100001100};
			assign coef[40] =   {12'b011111110000, 12'b111100000101};
			assign coef[41] =   {12'b011111101111, 12'b111011111111};
			assign coef[42] =   {12'b011111101110, 12'b111011111001};
			assign coef[43] =   {12'b011111101101, 12'b111011110011};
			assign coef[44] =   {12'b011111101100, 12'b111011101100};
			assign coef[45] =   {12'b011111101100, 12'b111011100110};
			assign coef[46] =   {12'b011111101011, 12'b111011100000};
			assign coef[47] =   {12'b011111101010, 12'b111011011010};
			assign coef[48] =   {12'b011111101001, 12'b111011010100};
			assign coef[49] =   {12'b011111101000, 12'b111011001101};
			assign coef[50] =   {12'b011111100111, 12'b111011000111};
			assign coef[51] =   {12'b011111100110, 12'b111011000001};
			assign coef[52] =   {12'b011111100101, 12'b111010111011};
			assign coef[53] =   {12'b011111100100, 12'b111010110101};
			assign coef[54] =   {12'b011111100011, 12'b111010101110};
			assign coef[55] =   {12'b011111100010, 12'b111010101000};
			assign coef[56] =   {12'b011111100001, 12'b111010100010};
			assign coef[57] =   {12'b011111100000, 12'b111010011100};
			assign coef[58] =   {12'b011111011111, 12'b111010010110};
			assign coef[59] =   {12'b011111011110, 12'b111010001111};
			assign coef[60] =   {12'b011111011100, 12'b111010001001};
			assign coef[61] =   {12'b011111011011, 12'b111010000011};
			assign coef[62] =   {12'b011111011010, 12'b111001111101};
			assign coef[63] =   {12'b011111011001, 12'b111001110111};
			assign coef[64] =   {12'b011111011000, 12'b111001110001};
			assign coef[65] =   {12'b011111010110, 12'b111001101010};
			assign coef[66] =   {12'b011111010101, 12'b111001100100};
			assign coef[67] =   {12'b011111010100, 12'b111001011110};
			assign coef[68] =   {12'b011111010011, 12'b111001011000};
			assign coef[69] =   {12'b011111010001, 12'b111001010010};
			assign coef[70] =   {12'b011111010000, 12'b111001001100};
			assign coef[71] =   {12'b011111001111, 12'b111001000110};
			assign coef[72] =   {12'b011111001101, 12'b111000111111};
			assign coef[73] =   {12'b011111001100, 12'b111000111001};
			assign coef[74] =   {12'b011111001011, 12'b111000110011};
			assign coef[75] =   {12'b011111001001, 12'b111000101101};
			assign coef[76] =   {12'b011111001000, 12'b111000100111};
			assign coef[77] =   {12'b011111000110, 12'b111000100001};
			assign coef[78] =   {12'b011111000101, 12'b111000011011};
			assign coef[79] =   {12'b011111000011, 12'b111000010101};
			assign coef[80] =   {12'b011111000010, 12'b111000001111};
			assign coef[81] =   {12'b011111000000, 12'b111000001000};
			assign coef[82] =   {12'b011110111111, 12'b111000000010};
			assign coef[83] =   {12'b011110111101, 12'b110111111100};
			assign coef[84] =   {12'b011110111011, 12'b110111110110};
			assign coef[85] =   {12'b011110111010, 12'b110111110000};
			assign coef[86] =   {12'b011110111000, 12'b110111101010};
			assign coef[87] =   {12'b011110110111, 12'b110111100100};
			assign coef[88] =   {12'b011110110101, 12'b110111011110};
			assign coef[89] =   {12'b011110110011, 12'b110111011000};
			assign coef[90] =   {12'b011110110010, 12'b110111010010};
			assign coef[91] =   {12'b011110110000, 12'b110111001100};
			assign coef[92] =   {12'b011110101110, 12'b110111000110};
			assign coef[93] =   {12'b011110101100, 12'b110111000000};
			assign coef[94] =   {12'b011110101011, 12'b110110111010};
			assign coef[95] =   {12'b011110101001, 12'b110110110100};
			assign coef[96] =   {12'b011110100111, 12'b110110101110};
			assign coef[97] =   {12'b011110100101, 12'b110110101000};
			assign coef[98] =   {12'b011110100011, 12'b110110100010};
			assign coef[99] =   {12'b011110100001, 12'b110110011100};
			assign coef[100] =  {12'b011110011111, 12'b110110010110};
			assign coef[101] =  {12'b011110011110, 12'b110110010000};
			assign coef[102] =  {12'b011110011100, 12'b110110001010};
			assign coef[103] =  {12'b011110011010, 12'b110110000100};
			assign coef[104] =  {12'b011110011000, 12'b110101111110};
			assign coef[105] =  {12'b011110010110, 12'b110101111000};
			assign coef[106] =  {12'b011110010100, 12'b110101110010};
			assign coef[107] =  {12'b011110010010, 12'b110101101100};
			assign coef[108] =  {12'b011110010000, 12'b110101100110};
			assign coef[109] =  {12'b011110001110, 12'b110101100000};
			assign coef[110] =  {12'b011110001100, 12'b110101011010};
			assign coef[111] =  {12'b011110001001, 12'b110101010100};
			assign coef[112] =  {12'b011110000111, 12'b110101001110};
			assign coef[113] =  {12'b011110000101, 12'b110101001000};
			assign coef[114] =  {12'b011110000011, 12'b110101000011};
			assign coef[115] =  {12'b011110000001, 12'b110100111101};
			assign coef[116] =  {12'b011101111111, 12'b110100110111};
			assign coef[117] =  {12'b011101111101, 12'b110100110001};
			assign coef[118] =  {12'b011101111010, 12'b110100101011};
			assign coef[119] =  {12'b011101111000, 12'b110100100101};
			assign coef[120] =  {12'b011101110110, 12'b110100011111};
			assign coef[121] =  {12'b011101110100, 12'b110100011001};
			assign coef[122] =  {12'b011101110001, 12'b110100010100};
			assign coef[123] =  {12'b011101101111, 12'b110100001110};
			assign coef[124] =  {12'b011101101101, 12'b110100001000};
			assign coef[125] =  {12'b011101101010, 12'b110100000010};
			assign coef[126] =  {12'b011101101000, 12'b110011111100};
			assign coef[127] =  {12'b011101100110, 12'b110011110110};
			assign coef[128] =  {12'b011101100011, 12'b110011110001};
			assign coef[129] =  {12'b011101100001, 12'b110011101011};
			assign coef[130] =  {12'b011101011110, 12'b110011100101};
			assign coef[131] =  {12'b011101011100, 12'b110011011111};
			assign coef[132] =  {12'b011101011001, 12'b110011011001};
			assign coef[133] =  {12'b011101010111, 12'b110011010100};
			assign coef[134] =  {12'b011101010100, 12'b110011001110};
			assign coef[135] =  {12'b011101010010, 12'b110011001000};
			assign coef[136] =  {12'b011101001111, 12'b110011000010};
			assign coef[137] =  {12'b011101001101, 12'b110010111101};
			assign coef[138] =  {12'b011101001010, 12'b110010110111};
			assign coef[139] =  {12'b011101001000, 12'b110010110001};
			assign coef[140] =  {12'b011101000101, 12'b110010101100};
			assign coef[141] =  {12'b011101000010, 12'b110010100110};
			assign coef[142] =  {12'b011101000000, 12'b110010100000};
			assign coef[143] =  {12'b011100111101, 12'b110010011010};
			assign coef[144] =  {12'b011100111011, 12'b110010010101};
			assign coef[145] =  {12'b011100111000, 12'b110010001111};
			assign coef[146] =  {12'b011100110101, 12'b110010001001};
			assign coef[147] =  {12'b011100110010, 12'b110010000100};
			assign coef[148] =  {12'b011100110000, 12'b110001111110};
			assign coef[149] =  {12'b011100101101, 12'b110001111000};
			assign coef[150] =  {12'b011100101010, 12'b110001110011};
			assign coef[151] =  {12'b011100100111, 12'b110001101101};
			assign coef[152] =  {12'b011100100100, 12'b110001101000};
			assign coef[153] =  {12'b011100100010, 12'b110001100010};
			assign coef[154] =  {12'b011100011111, 12'b110001011100};
			assign coef[155] =  {12'b011100011100, 12'b110001010111};
			assign coef[156] =  {12'b011100011001, 12'b110001010001};
			assign coef[157] =  {12'b011100010110, 12'b110001001100};
			assign coef[158] =  {12'b011100010011, 12'b110001000110};
			assign coef[159] =  {12'b011100010000, 12'b110001000001};
			assign coef[160] =  {12'b011100001101, 12'b110000111011};
			assign coef[161] =  {12'b011100001010, 12'b110000110101};
			assign coef[162] =  {12'b011100000111, 12'b110000110000};
			assign coef[163] =  {12'b011100000100, 12'b110000101010};
			assign coef[164] =  {12'b011100000001, 12'b110000100101};
			assign coef[165] =  {12'b011011111110, 12'b110000011111};
			assign coef[166] =  {12'b011011111011, 12'b110000011010};
			assign coef[167] =  {12'b011011111000, 12'b110000010100};
			assign coef[168] =  {12'b011011110101, 12'b110000001111};
			assign coef[169] =  {12'b011011110010, 12'b110000001010};
			assign coef[170] =  {12'b011011101111, 12'b110000000100};
			assign coef[171] =  {12'b011011101100, 12'b101111111111};
			assign coef[172] =  {12'b011011101001, 12'b101111111001};
			assign coef[173] =  {12'b011011100101, 12'b101111110100};
			assign coef[174] =  {12'b011011100010, 12'b101111101110};
			assign coef[175] =  {12'b011011011111, 12'b101111101001};
			assign coef[176] =  {12'b011011011100, 12'b101111100100};
			assign coef[177] =  {12'b011011011001, 12'b101111011110};
			assign coef[178] =  {12'b011011010101, 12'b101111011001};
			assign coef[179] =  {12'b011011010010, 12'b101111010011};
			assign coef[180] =  {12'b011011001111, 12'b101111001110};
			assign coef[181] =  {12'b011011001011, 12'b101111001001};
			assign coef[182] =  {12'b011011001000, 12'b101111000011};
			assign coef[183] =  {12'b011011000101, 12'b101110111110};
			assign coef[184] =  {12'b011011000001, 12'b101110111001};
			assign coef[185] =  {12'b011010111110, 12'b101110110100};
			assign coef[186] =  {12'b011010111011, 12'b101110101110};
			assign coef[187] =  {12'b011010110111, 12'b101110101001};
			assign coef[188] =  {12'b011010110100, 12'b101110100100};
			assign coef[189] =  {12'b011010110000, 12'b101110011110};
			assign coef[190] =  {12'b011010101101, 12'b101110011001};
			assign coef[191] =  {12'b011010101010, 12'b101110010100};
			assign coef[192] =  {12'b011010100110, 12'b101110001111};
			assign coef[193] =  {12'b011010100011, 12'b101110001001};
			assign coef[194] =  {12'b011010011111, 12'b101110000100};
			assign coef[195] =  {12'b011010011100, 12'b101101111111};
			assign coef[196] =  {12'b011010011000, 12'b101101111010};
			assign coef[197] =  {12'b011010010100, 12'b101101110101};
			assign coef[198] =  {12'b011010010001, 12'b101101110000};
			assign coef[199] =  {12'b011010001101, 12'b101101101010};
			assign coef[200] =  {12'b011010001010, 12'b101101100101};
			assign coef[201] =  {12'b011010000110, 12'b101101100000};
			assign coef[202] =  {12'b011010000010, 12'b101101011011};
			assign coef[203] =  {12'b011001111111, 12'b101101010110};
			assign coef[204] =  {12'b011001111011, 12'b101101010001};
			assign coef[205] =  {12'b011001110111, 12'b101101001100};
			assign coef[206] =  {12'b011001110100, 12'b101101000111};
			assign coef[207] =  {12'b011001110000, 12'b101101000010};
			assign coef[208] =  {12'b011001101100, 12'b101100111101};
			assign coef[209] =  {12'b011001101000, 12'b101100111000};
			assign coef[210] =  {12'b011001100101, 12'b101100110010};
			assign coef[211] =  {12'b011001100001, 12'b101100101101};
			assign coef[212] =  {12'b011001011101, 12'b101100101000};
			assign coef[213] =  {12'b011001011001, 12'b101100100011};
			assign coef[214] =  {12'b011001010101, 12'b101100011110};
			assign coef[215] =  {12'b011001010010, 12'b101100011010};
			assign coef[216] =  {12'b011001001110, 12'b101100010101};
			assign coef[217] =  {12'b011001001010, 12'b101100010000};
			assign coef[218] =  {12'b011001000110, 12'b101100001011};
			assign coef[219] =  {12'b011001000010, 12'b101100000110};
			assign coef[220] =  {12'b011000111110, 12'b101100000001};
			assign coef[221] =  {12'b011000111010, 12'b101011111100};
			assign coef[222] =  {12'b011000110110, 12'b101011110111};
			assign coef[223] =  {12'b011000110010, 12'b101011110010};
			assign coef[224] =  {12'b011000101110, 12'b101011101101};
			assign coef[225] =  {12'b011000101010, 12'b101011101000};
			assign coef[226] =  {12'b011000100110, 12'b101011100100};
			assign coef[227] =  {12'b011000100010, 12'b101011011111};
			assign coef[228] =  {12'b011000011110, 12'b101011011010};
			assign coef[229] =  {12'b011000011010, 12'b101011010101};
			assign coef[230] =  {12'b011000010110, 12'b101011010000};
			assign coef[231] =  {12'b011000010010, 12'b101011001100};
			assign coef[232] =  {12'b011000001110, 12'b101011000111};
			assign coef[233] =  {12'b011000001010, 12'b101011000010};
			assign coef[234] =  {12'b011000000110, 12'b101010111101};
			assign coef[235] =  {12'b011000000010, 12'b101010111001};
			assign coef[236] =  {12'b010111111110, 12'b101010110100};
			assign coef[237] =  {12'b010111111001, 12'b101010101111};
			assign coef[238] =  {12'b010111110101, 12'b101010101011};
			assign coef[239] =  {12'b010111110001, 12'b101010100110};
			assign coef[240] =  {12'b010111101101, 12'b101010100001};
			assign coef[241] =  {12'b010111101001, 12'b101010011101};
			assign coef[242] =  {12'b010111100100, 12'b101010011000};
			assign coef[243] =  {12'b010111100000, 12'b101010010011};
			assign coef[244] =  {12'b010111011100, 12'b101010001111};
			assign coef[245] =  {12'b010111011000, 12'b101010001010};
			assign coef[246] =  {12'b010111010011, 12'b101010000110};
			assign coef[247] =  {12'b010111001111, 12'b101010000001};
			assign coef[248] =  {12'b010111001011, 12'b101001111100};
			assign coef[249] =  {12'b010111000110, 12'b101001111000};
			assign coef[250] =  {12'b010111000010, 12'b101001110011};
			assign coef[251] =  {12'b010110111110, 12'b101001101111};
			assign coef[252] =  {12'b010110111001, 12'b101001101010};
			assign coef[253] =  {12'b010110110101, 12'b101001100110};
			assign coef[254] =  {12'b010110110000, 12'b101001100001};
			assign coef[255] =  {12'b010110101100, 12'b101001011101};
			assign coef[256] =  {12'b010110100111, 12'b101001011001};
			assign coef[257] =  {12'b010110100011, 12'b101001010100};
			assign coef[258] =  {12'b010110011111, 12'b101001010000};
			assign coef[259] =  {12'b010110011010, 12'b101001001011};
			assign coef[260] =  {12'b010110010110, 12'b101001000111};
			assign coef[261] =  {12'b010110010001, 12'b101001000010};
			assign coef[262] =  {12'b010110001101, 12'b101000111110};
			assign coef[263] =  {12'b010110001000, 12'b101000111010};
			assign coef[264] =  {12'b010110000100, 12'b101000110101};
			assign coef[265] =  {12'b010101111111, 12'b101000110001};
			assign coef[266] =  {12'b010101111010, 12'b101000101101};
			assign coef[267] =  {12'b010101110110, 12'b101000101000};
			assign coef[268] =  {12'b010101110001, 12'b101000100100};
			assign coef[269] =  {12'b010101101101, 12'b101000100000};
			assign coef[270] =  {12'b010101101000, 12'b101000011100};
			assign coef[271] =  {12'b010101100011, 12'b101000010111};
			assign coef[272] =  {12'b010101011111, 12'b101000010011};
			assign coef[273] =  {12'b010101011010, 12'b101000001111};
			assign coef[274] =  {12'b010101010101, 12'b101000001011};
			assign coef[275] =  {12'b010101010001, 12'b101000000111};
			assign coef[276] =  {12'b010101001100, 12'b101000000010};
			assign coef[277] =  {12'b010101000111, 12'b100111111110};
			assign coef[278] =  {12'b010101000011, 12'b100111111010};
			assign coef[279] =  {12'b010100111110, 12'b100111110110};
			assign coef[280] =  {12'b010100111001, 12'b100111110010};
			assign coef[281] =  {12'b010100110100, 12'b100111101110};
			assign coef[282] =  {12'b010100110000, 12'b100111101010};
			assign coef[283] =  {12'b010100101011, 12'b100111100110};
			assign coef[284] =  {12'b010100100110, 12'b100111100010};
			assign coef[285] =  {12'b010100100001, 12'b100111011110};
			assign coef[286] =  {12'b010100011100, 12'b100111011010};
			assign coef[287] =  {12'b010100011000, 12'b100111010110};
			assign coef[288] =  {12'b010100010011, 12'b100111010010};
			assign coef[289] =  {12'b010100001110, 12'b100111001110};
			assign coef[290] =  {12'b010100001001, 12'b100111001010};
			assign coef[291] =  {12'b010100000100, 12'b100111000110};
			assign coef[292] =  {12'b010011111111, 12'b100111000010};
			assign coef[293] =  {12'b010011111010, 12'b100110111110};
			assign coef[294] =  {12'b010011110101, 12'b100110111010};
			assign coef[295] =  {12'b010011110000, 12'b100110110110};
			assign coef[296] =  {12'b010011101011, 12'b100110110010};
			assign coef[297] =  {12'b010011100110, 12'b100110101110};
			assign coef[298] =  {12'b010011100010, 12'b100110101011};
			assign coef[299] =  {12'b010011011101, 12'b100110100111};
			assign coef[300] =  {12'b010011011000, 12'b100110100011};
			assign coef[301] =  {12'b010011010011, 12'b100110011111};
			assign coef[302] =  {12'b010011001110, 12'b100110011011};
			assign coef[303] =  {12'b010011001000, 12'b100110011000};
			assign coef[304] =  {12'b010011000011, 12'b100110010100};
			assign coef[305] =  {12'b010010111110, 12'b100110010000};
			assign coef[306] =  {12'b010010111001, 12'b100110001100};
			assign coef[307] =  {12'b010010110100, 12'b100110001001};
			assign coef[308] =  {12'b010010101111, 12'b100110000101};
			assign coef[309] =  {12'b010010101010, 12'b100110000001};
			assign coef[310] =  {12'b010010100101, 12'b100101111110};
			assign coef[311] =  {12'b010010100000, 12'b100101111010};
			assign coef[312] =  {12'b010010011011, 12'b100101110110};
			assign coef[313] =  {12'b010010010110, 12'b100101110011};
			assign coef[314] =  {12'b010010010000, 12'b100101101111};
			assign coef[315] =  {12'b010010001011, 12'b100101101100};
			assign coef[316] =  {12'b010010000110, 12'b100101101000};
			assign coef[317] =  {12'b010010000001, 12'b100101100100};
			assign coef[318] =  {12'b010001111100, 12'b100101100001};
			assign coef[319] =  {12'b010001110111, 12'b100101011101};
			assign coef[320] =  {12'b010001110001, 12'b100101011010};
			assign coef[321] =  {12'b010001101100, 12'b100101010110};
			assign coef[322] =  {12'b010001100111, 12'b100101010011};
			assign coef[323] =  {12'b010001100010, 12'b100101010000};
			assign coef[324] =  {12'b010001011100, 12'b100101001100};
			assign coef[325] =  {12'b010001010111, 12'b100101001001};
			assign coef[326] =  {12'b010001010010, 12'b100101000101};
			assign coef[327] =  {12'b010001001100, 12'b100101000010};
			assign coef[328] =  {12'b010001000111, 12'b100100111111};
			assign coef[329] =  {12'b010001000010, 12'b100100111011};
			assign coef[330] =  {12'b010000111101, 12'b100100111000};
			assign coef[331] =  {12'b010000110111, 12'b100100110101};
			assign coef[332] =  {12'b010000110010, 12'b100100110001};
			assign coef[333] =  {12'b010000101101, 12'b100100101110};
			assign coef[334] =  {12'b010000100111, 12'b100100101011};
			assign coef[335] =  {12'b010000100010, 12'b100100100111};
			assign coef[336] =  {12'b010000011100, 12'b100100100100};
			assign coef[337] =  {12'b010000010111, 12'b100100100001};
			assign coef[338] =  {12'b010000010010, 12'b100100011110};
			assign coef[339] =  {12'b010000001100, 12'b100100011011};
			assign coef[340] =  {12'b010000000111, 12'b100100010111};
			assign coef[341] =  {12'b010000000001, 12'b100100010100};
			assign coef[342] =  {12'b001111111100, 12'b100100010001};
			assign coef[343] =  {12'b001111110110, 12'b100100001110};
			assign coef[344] =  {12'b001111110001, 12'b100100001011};
			assign coef[345] =  {12'b001111101100, 12'b100100001000};
			assign coef[346] =  {12'b001111100110, 12'b100100000101};
			assign coef[347] =  {12'b001111100001, 12'b100100000010};
			assign coef[348] =  {12'b001111011011, 12'b100011111111};
			assign coef[349] =  {12'b001111010110, 12'b100011111100};
			assign coef[350] =  {12'b001111010000, 12'b100011111001};
			assign coef[351] =  {12'b001111001011, 12'b100011110110};
			assign coef[352] =  {12'b001111000101, 12'b100011110011};
			assign coef[353] =  {12'b001110111111, 12'b100011110000};
			assign coef[354] =  {12'b001110111010, 12'b100011101101};
			assign coef[355] =  {12'b001110110100, 12'b100011101010};
			assign coef[356] =  {12'b001110101111, 12'b100011100111};
			assign coef[357] =  {12'b001110101001, 12'b100011100100};
			assign coef[358] =  {12'b001110100100, 12'b100011100001};
			assign coef[359] =  {12'b001110011110, 12'b100011011110};
			assign coef[360] =  {12'b001110011000, 12'b100011011100};
			assign coef[361] =  {12'b001110010011, 12'b100011011001};
			assign coef[362] =  {12'b001110001101, 12'b100011010110};
			assign coef[363] =  {12'b001110001000, 12'b100011010011};
			assign coef[364] =  {12'b001110000010, 12'b100011010000};
			assign coef[365] =  {12'b001101111100, 12'b100011001110};
			assign coef[366] =  {12'b001101110111, 12'b100011001011};
			assign coef[367] =  {12'b001101110001, 12'b100011001000};
			assign coef[368] =  {12'b001101101011, 12'b100011000101};
			assign coef[369] =  {12'b001101100110, 12'b100011000011};
			assign coef[370] =  {12'b001101100000, 12'b100011000000};
			assign coef[371] =  {12'b001101011010, 12'b100010111110};
			assign coef[372] =  {12'b001101010100, 12'b100010111011};
			assign coef[373] =  {12'b001101001111, 12'b100010111000};
			assign coef[374] =  {12'b001101001001, 12'b100010110110};
			assign coef[375] =  {12'b001101000011, 12'b100010110011};
			assign coef[376] =  {12'b001100111110, 12'b100010110001};
			assign coef[377] =  {12'b001100111000, 12'b100010101110};
			assign coef[378] =  {12'b001100110010, 12'b100010101100};
			assign coef[379] =  {12'b001100101100, 12'b100010101001};
			assign coef[380] =  {12'b001100100111, 12'b100010100111};
			assign coef[381] =  {12'b001100100001, 12'b100010100100};
			assign coef[382] =  {12'b001100011011, 12'b100010100010};
			assign coef[383] =  {12'b001100010101, 12'b100010011111};
			assign coef[384] =  {12'b001100001111, 12'b100010011101};
			assign coef[385] =  {12'b001100001010, 12'b100010011010};
			assign coef[386] =  {12'b001100000100, 12'b100010011000};
			assign coef[387] =  {12'b001011111110, 12'b100010010110};
			assign coef[388] =  {12'b001011111000, 12'b100010010011};
			assign coef[389] =  {12'b001011110010, 12'b100010010001};
			assign coef[390] =  {12'b001011101100, 12'b100010001111};
			assign coef[391] =  {12'b001011100111, 12'b100010001100};
			assign coef[392] =  {12'b001011100001, 12'b100010001010};
			assign coef[393] =  {12'b001011011011, 12'b100010001000};
			assign coef[394] =  {12'b001011010101, 12'b100010000110};
			assign coef[395] =  {12'b001011001111, 12'b100010000011};
			assign coef[396] =  {12'b001011001001, 12'b100010000001};
			assign coef[397] =  {12'b001011000011, 12'b100001111111};
			assign coef[398] =  {12'b001010111101, 12'b100001111101};
			assign coef[399] =  {12'b001010111000, 12'b100001111011};
			assign coef[400] =  {12'b001010110010, 12'b100001111001};
			assign coef[401] =  {12'b001010101100, 12'b100001110111};
			assign coef[402] =  {12'b001010100110, 12'b100001110100};
			assign coef[403] =  {12'b001010100000, 12'b100001110010};
			assign coef[404] =  {12'b001010011010, 12'b100001110000};
			assign coef[405] =  {12'b001010010100, 12'b100001101110};
			assign coef[406] =  {12'b001010001110, 12'b100001101100};
			assign coef[407] =  {12'b001010001000, 12'b100001101010};
			assign coef[408] =  {12'b001010000010, 12'b100001101000};
			assign coef[409] =  {12'b001001111100, 12'b100001100110};
			assign coef[410] =  {12'b001001110110, 12'b100001100100};
			assign coef[411] =  {12'b001001110000, 12'b100001100010};
			assign coef[412] =  {12'b001001101010, 12'b100001100001};
			assign coef[413] =  {12'b001001100100, 12'b100001011111};
			assign coef[414] =  {12'b001001011110, 12'b100001011101};
			assign coef[415] =  {12'b001001011000, 12'b100001011011};
			assign coef[416] =  {12'b001001010010, 12'b100001011001};
			assign coef[417] =  {12'b001001001100, 12'b100001010111};
			assign coef[418] =  {12'b001001000110, 12'b100001010101};
			assign coef[419] =  {12'b001001000000, 12'b100001010100};
			assign coef[420] =  {12'b001000111010, 12'b100001010010};
			assign coef[421] =  {12'b001000110100, 12'b100001010000};
			assign coef[422] =  {12'b001000101110, 12'b100001001110};
			assign coef[423] =  {12'b001000101000, 12'b100001001101};
			assign coef[424] =  {12'b001000100010, 12'b100001001011};
			assign coef[425] =  {12'b001000011100, 12'b100001001001};
			assign coef[426] =  {12'b001000010110, 12'b100001001000};
			assign coef[427] =  {12'b001000010000, 12'b100001000110};
			assign coef[428] =  {12'b001000001010, 12'b100001000101};
			assign coef[429] =  {12'b001000000100, 12'b100001000011};
			assign coef[430] =  {12'b000111111110, 12'b100001000001};
			assign coef[431] =  {12'b000111111000, 12'b100001000000};
			assign coef[432] =  {12'b000111110001, 12'b100000111110};
			assign coef[433] =  {12'b000111101011, 12'b100000111101};
			assign coef[434] =  {12'b000111100101, 12'b100000111011};
			assign coef[435] =  {12'b000111011111, 12'b100000111010};
			assign coef[436] =  {12'b000111011001, 12'b100000111000};
			assign coef[437] =  {12'b000111010011, 12'b100000110111};
			assign coef[438] =  {12'b000111001101, 12'b100000110101};
			assign coef[439] =  {12'b000111000111, 12'b100000110100};
			assign coef[440] =  {12'b000111000001, 12'b100000110011};
			assign coef[441] =  {12'b000110111010, 12'b100000110001};
			assign coef[442] =  {12'b000110110100, 12'b100000110000};
			assign coef[443] =  {12'b000110101110, 12'b100000101111};
			assign coef[444] =  {12'b000110101000, 12'b100000101101};
			assign coef[445] =  {12'b000110100010, 12'b100000101100};
			assign coef[446] =  {12'b000110011100, 12'b100000101011};
			assign coef[447] =  {12'b000110010110, 12'b100000101010};
			assign coef[448] =  {12'b000110001111, 12'b100000101000};
			assign coef[449] =  {12'b000110001001, 12'b100000100111};
			assign coef[450] =  {12'b000110000011, 12'b100000100110};
			assign coef[451] =  {12'b000101111101, 12'b100000100101};
			assign coef[452] =  {12'b000101110111, 12'b100000100100};
			assign coef[453] =  {12'b000101110001, 12'b100000100010};
			assign coef[454] =  {12'b000101101010, 12'b100000100001};
			assign coef[455] =  {12'b000101100100, 12'b100000100000};
			assign coef[456] =  {12'b000101011110, 12'b100000011111};
			assign coef[457] =  {12'b000101011000, 12'b100000011110};
			assign coef[458] =  {12'b000101010010, 12'b100000011101};
			assign coef[459] =  {12'b000101001011, 12'b100000011100};
			assign coef[460] =  {12'b000101000101, 12'b100000011011};
			assign coef[461] =  {12'b000100111111, 12'b100000011010};
			assign coef[462] =  {12'b000100111001, 12'b100000011001};
			assign coef[463] =  {12'b000100110011, 12'b100000011000};
			assign coef[464] =  {12'b000100101100, 12'b100000010111};
			assign coef[465] =  {12'b000100100110, 12'b100000010110};
			assign coef[466] =  {12'b000100100000, 12'b100000010101};
			assign coef[467] =  {12'b000100011010, 12'b100000010100};
			assign coef[468] =  {12'b000100010100, 12'b100000010100};
			assign coef[469] =  {12'b000100001101, 12'b100000010011};
			assign coef[470] =  {12'b000100000111, 12'b100000010010};
			assign coef[471] =  {12'b000100000001, 12'b100000010001};
			assign coef[472] =  {12'b000011111011, 12'b100000010000};
			assign coef[473] =  {12'b000011110100, 12'b100000010000};
			assign coef[474] =  {12'b000011101110, 12'b100000001111};
			assign coef[475] =  {12'b000011101000, 12'b100000001110};
			assign coef[476] =  {12'b000011100010, 12'b100000001101};
			assign coef[477] =  {12'b000011011011, 12'b100000001101};
			assign coef[478] =  {12'b000011010101, 12'b100000001100};
			assign coef[479] =  {12'b000011001111, 12'b100000001011};
			assign coef[480] =  {12'b000011001001, 12'b100000001011};
			assign coef[481] =  {12'b000011000010, 12'b100000001010};
			assign coef[482] =  {12'b000010111100, 12'b100000001010};
			assign coef[483] =  {12'b000010110110, 12'b100000001001};
			assign coef[484] =  {12'b000010110000, 12'b100000001000};
			assign coef[485] =  {12'b000010101001, 12'b100000001000};
			assign coef[486] =  {12'b000010100011, 12'b100000000111};
			assign coef[487] =  {12'b000010011101, 12'b100000000111};
			assign coef[488] =  {12'b000010010111, 12'b100000000110};
			assign coef[489] =  {12'b000010010000, 12'b100000000110};
			assign coef[490] =  {12'b000010001010, 12'b100000000110};
			assign coef[491] =  {12'b000010000100, 12'b100000000101};
			assign coef[492] =  {12'b000001111110, 12'b100000000101};
			assign coef[493] =  {12'b000001110111, 12'b100000000100};
			assign coef[494] =  {12'b000001110001, 12'b100000000100};
			assign coef[495] =  {12'b000001101011, 12'b100000000100};
			assign coef[496] =  {12'b000001100100, 12'b100000000011};
			assign coef[497] =  {12'b000001011110, 12'b100000000011};
			assign coef[498] =  {12'b000001011000, 12'b100000000011};
			assign coef[499] =  {12'b000001010010, 12'b100000000011};
			assign coef[500] =  {12'b000001001011, 12'b100000000010};
			assign coef[501] =  {12'b000001000101, 12'b100000000010};
			assign coef[502] =  {12'b000000111111, 12'b100000000010};
			assign coef[503] =  {12'b000000111001, 12'b100000000010};
			assign coef[504] =  {12'b000000110010, 12'b100000000010};
			assign coef[505] =  {12'b000000101100, 12'b100000000001};
			assign coef[506] =  {12'b000000100110, 12'b100000000001};
			assign coef[507] =  {12'b000000011111, 12'b100000000001};
			assign coef[508] =  {12'b000000011001, 12'b100000000001};
			assign coef[509] =  {12'b000000010011, 12'b100000000001};
			assign coef[510] =  {12'b000000001101, 12'b100000000001};
			assign coef[511] =  {12'b000000000110, 12'b100000000001};
			assign coef[512] =  {12'b000000000000, 12'b100000000001};
			assign coef[513] =  {12'b111111111010, 12'b100000000001};
			assign coef[514] =  {12'b111111110011, 12'b100000000001};
			assign coef[515] =  {12'b111111101101, 12'b100000000001};
			assign coef[516] =  {12'b111111100111, 12'b100000000001};
			assign coef[517] =  {12'b111111100001, 12'b100000000001};
			assign coef[518] =  {12'b111111011010, 12'b100000000001};
			assign coef[519] =  {12'b111111010100, 12'b100000000001};
			assign coef[520] =  {12'b111111001110, 12'b100000000010};
			assign coef[521] =  {12'b111111000111, 12'b100000000010};
			assign coef[522] =  {12'b111111000001, 12'b100000000010};
			assign coef[523] =  {12'b111110111011, 12'b100000000010};
			assign coef[524] =  {12'b111110110101, 12'b100000000010};
			assign coef[525] =  {12'b111110101110, 12'b100000000011};
			assign coef[526] =  {12'b111110101000, 12'b100000000011};
			assign coef[527] =  {12'b111110100010, 12'b100000000011};
			assign coef[528] =  {12'b111110011100, 12'b100000000011};
			assign coef[529] =  {12'b111110010101, 12'b100000000100};
			assign coef[530] =  {12'b111110001111, 12'b100000000100};
			assign coef[531] =  {12'b111110001001, 12'b100000000100};
			assign coef[532] =  {12'b111110000010, 12'b100000000101};
			assign coef[533] =  {12'b111101111100, 12'b100000000101};
			assign coef[534] =  {12'b111101110110, 12'b100000000110};
			assign coef[535] =  {12'b111101110000, 12'b100000000110};
			assign coef[536] =  {12'b111101101001, 12'b100000000110};
			assign coef[537] =  {12'b111101100011, 12'b100000000111};
			assign coef[538] =  {12'b111101011101, 12'b100000000111};
			assign coef[539] =  {12'b111101010111, 12'b100000001000};
			assign coef[540] =  {12'b111101010000, 12'b100000001000};
			assign coef[541] =  {12'b111101001010, 12'b100000001001};
			assign coef[542] =  {12'b111101000100, 12'b100000001010};
			assign coef[543] =  {12'b111100111110, 12'b100000001010};
			assign coef[544] =  {12'b111100110111, 12'b100000001011};
			assign coef[545] =  {12'b111100110001, 12'b100000001011};
			assign coef[546] =  {12'b111100101011, 12'b100000001100};
			assign coef[547] =  {12'b111100100101, 12'b100000001101};
			assign coef[548] =  {12'b111100011110, 12'b100000001101};
			assign coef[549] =  {12'b111100011000, 12'b100000001110};
			assign coef[550] =  {12'b111100010010, 12'b100000001111};
			assign coef[551] =  {12'b111100001100, 12'b100000010000};
			assign coef[552] =  {12'b111100000101, 12'b100000010000};
			assign coef[553] =  {12'b111011111111, 12'b100000010001};
			assign coef[554] =  {12'b111011111001, 12'b100000010010};
			assign coef[555] =  {12'b111011110011, 12'b100000010011};
			assign coef[556] =  {12'b111011101100, 12'b100000010100};
			assign coef[557] =  {12'b111011100110, 12'b100000010100};
			assign coef[558] =  {12'b111011100000, 12'b100000010101};
			assign coef[559] =  {12'b111011011010, 12'b100000010110};
			assign coef[560] =  {12'b111011010100, 12'b100000010111};
			assign coef[561] =  {12'b111011001101, 12'b100000011000};
			assign coef[562] =  {12'b111011000111, 12'b100000011001};
			assign coef[563] =  {12'b111011000001, 12'b100000011010};
			assign coef[564] =  {12'b111010111011, 12'b100000011011};
			assign coef[565] =  {12'b111010110101, 12'b100000011100};
			assign coef[566] =  {12'b111010101110, 12'b100000011101};
			assign coef[567] =  {12'b111010101000, 12'b100000011110};
			assign coef[568] =  {12'b111010100010, 12'b100000011111};
			assign coef[569] =  {12'b111010011100, 12'b100000100000};
			assign coef[570] =  {12'b111010010110, 12'b100000100001};
			assign coef[571] =  {12'b111010001111, 12'b100000100010};
			assign coef[572] =  {12'b111010001001, 12'b100000100100};
			assign coef[573] =  {12'b111010000011, 12'b100000100101};
			assign coef[574] =  {12'b111001111101, 12'b100000100110};
			assign coef[575] =  {12'b111001110111, 12'b100000100111};
			assign coef[576] =  {12'b111001110001, 12'b100000101000};
			assign coef[577] =  {12'b111001101010, 12'b100000101010};
			assign coef[578] =  {12'b111001100100, 12'b100000101011};
			assign coef[579] =  {12'b111001011110, 12'b100000101100};
			assign coef[580] =  {12'b111001011000, 12'b100000101101};
			assign coef[581] =  {12'b111001010010, 12'b100000101111};
			assign coef[582] =  {12'b111001001100, 12'b100000110000};
			assign coef[583] =  {12'b111001000110, 12'b100000110001};
			assign coef[584] =  {12'b111000111111, 12'b100000110011};
			assign coef[585] =  {12'b111000111001, 12'b100000110100};
			assign coef[586] =  {12'b111000110011, 12'b100000110101};
			assign coef[587] =  {12'b111000101101, 12'b100000110111};
			assign coef[588] =  {12'b111000100111, 12'b100000111000};
			assign coef[589] =  {12'b111000100001, 12'b100000111010};
			assign coef[590] =  {12'b111000011011, 12'b100000111011};
			assign coef[591] =  {12'b111000010101, 12'b100000111101};
			assign coef[592] =  {12'b111000001111, 12'b100000111110};
			assign coef[593] =  {12'b111000001000, 12'b100001000000};
			assign coef[594] =  {12'b111000000010, 12'b100001000001};
			assign coef[595] =  {12'b110111111100, 12'b100001000011};
			assign coef[596] =  {12'b110111110110, 12'b100001000101};
			assign coef[597] =  {12'b110111110000, 12'b100001000110};
			assign coef[598] =  {12'b110111101010, 12'b100001001000};
			assign coef[599] =  {12'b110111100100, 12'b100001001001};
			assign coef[600] =  {12'b110111011110, 12'b100001001011};
			assign coef[601] =  {12'b110111011000, 12'b100001001101};
			assign coef[602] =  {12'b110111010010, 12'b100001001110};
			assign coef[603] =  {12'b110111001100, 12'b100001010000};
			assign coef[604] =  {12'b110111000110, 12'b100001010010};
			assign coef[605] =  {12'b110111000000, 12'b100001010100};
			assign coef[606] =  {12'b110110111010, 12'b100001010101};
			assign coef[607] =  {12'b110110110100, 12'b100001010111};
			assign coef[608] =  {12'b110110101110, 12'b100001011001};
			assign coef[609] =  {12'b110110101000, 12'b100001011011};
			assign coef[610] =  {12'b110110100010, 12'b100001011101};
			assign coef[611] =  {12'b110110011100, 12'b100001011111};
			assign coef[612] =  {12'b110110010110, 12'b100001100001};
			assign coef[613] =  {12'b110110010000, 12'b100001100010};
			assign coef[614] =  {12'b110110001010, 12'b100001100100};
			assign coef[615] =  {12'b110110000100, 12'b100001100110};
			assign coef[616] =  {12'b110101111110, 12'b100001101000};
			assign coef[617] =  {12'b110101111000, 12'b100001101010};
			assign coef[618] =  {12'b110101110010, 12'b100001101100};
			assign coef[619] =  {12'b110101101100, 12'b100001101110};
			assign coef[620] =  {12'b110101100110, 12'b100001110000};
			assign coef[621] =  {12'b110101100000, 12'b100001110010};
			assign coef[622] =  {12'b110101011010, 12'b100001110100};
			assign coef[623] =  {12'b110101010100, 12'b100001110111};
			assign coef[624] =  {12'b110101001110, 12'b100001111001};
			assign coef[625] =  {12'b110101001000, 12'b100001111011};
			assign coef[626] =  {12'b110101000011, 12'b100001111101};
			assign coef[627] =  {12'b110100111101, 12'b100001111111};
			assign coef[628] =  {12'b110100110111, 12'b100010000001};
			assign coef[629] =  {12'b110100110001, 12'b100010000011};
			assign coef[630] =  {12'b110100101011, 12'b100010000110};
			assign coef[631] =  {12'b110100100101, 12'b100010001000};
			assign coef[632] =  {12'b110100011111, 12'b100010001010};
			assign coef[633] =  {12'b110100011001, 12'b100010001100};
			assign coef[634] =  {12'b110100010100, 12'b100010001111};
			assign coef[635] =  {12'b110100001110, 12'b100010010001};
			assign coef[636] =  {12'b110100001000, 12'b100010010011};
			assign coef[637] =  {12'b110100000010, 12'b100010010110};
			assign coef[638] =  {12'b110011111100, 12'b100010011000};
			assign coef[639] =  {12'b110011110110, 12'b100010011010};
			assign coef[640] =  {12'b110011110001, 12'b100010011101};
			assign coef[641] =  {12'b110011101011, 12'b100010011111};
			assign coef[642] =  {12'b110011100101, 12'b100010100010};
			assign coef[643] =  {12'b110011011111, 12'b100010100100};
			assign coef[644] =  {12'b110011011001, 12'b100010100111};
			assign coef[645] =  {12'b110011010100, 12'b100010101001};
			assign coef[646] =  {12'b110011001110, 12'b100010101100};
			assign coef[647] =  {12'b110011001000, 12'b100010101110};
			assign coef[648] =  {12'b110011000010, 12'b100010110001};
			assign coef[649] =  {12'b110010111101, 12'b100010110011};
			assign coef[650] =  {12'b110010110111, 12'b100010110110};
			assign coef[651] =  {12'b110010110001, 12'b100010111000};
			assign coef[652] =  {12'b110010101100, 12'b100010111011};
			assign coef[653] =  {12'b110010100110, 12'b100010111110};
			assign coef[654] =  {12'b110010100000, 12'b100011000000};
			assign coef[655] =  {12'b110010011010, 12'b100011000011};
			assign coef[656] =  {12'b110010010101, 12'b100011000101};
			assign coef[657] =  {12'b110010001111, 12'b100011001000};
			assign coef[658] =  {12'b110010001001, 12'b100011001011};
			assign coef[659] =  {12'b110010000100, 12'b100011001110};
			assign coef[660] =  {12'b110001111110, 12'b100011010000};
			assign coef[661] =  {12'b110001111000, 12'b100011010011};
			assign coef[662] =  {12'b110001110011, 12'b100011010110};
			assign coef[663] =  {12'b110001101101, 12'b100011011001};
			assign coef[664] =  {12'b110001101000, 12'b100011011100};
			assign coef[665] =  {12'b110001100010, 12'b100011011110};
			assign coef[666] =  {12'b110001011100, 12'b100011100001};
			assign coef[667] =  {12'b110001010111, 12'b100011100100};
			assign coef[668] =  {12'b110001010001, 12'b100011100111};
			assign coef[669] =  {12'b110001001100, 12'b100011101010};
			assign coef[670] =  {12'b110001000110, 12'b100011101101};
			assign coef[671] =  {12'b110001000001, 12'b100011110000};
			assign coef[672] =  {12'b110000111011, 12'b100011110011};
			assign coef[673] =  {12'b110000110101, 12'b100011110110};
			assign coef[674] =  {12'b110000110000, 12'b100011111001};
			assign coef[675] =  {12'b110000101010, 12'b100011111100};
			assign coef[676] =  {12'b110000100101, 12'b100011111111};
			assign coef[677] =  {12'b110000011111, 12'b100100000010};
			assign coef[678] =  {12'b110000011010, 12'b100100000101};
			assign coef[679] =  {12'b110000010100, 12'b100100001000};
			assign coef[680] =  {12'b110000001111, 12'b100100001011};
			assign coef[681] =  {12'b110000001010, 12'b100100001110};
			assign coef[682] =  {12'b110000000100, 12'b100100010001};
			assign coef[683] =  {12'b101111111111, 12'b100100010100};
			assign coef[684] =  {12'b101111111001, 12'b100100010111};
			assign coef[685] =  {12'b101111110100, 12'b100100011011};
			assign coef[686] =  {12'b101111101110, 12'b100100011110};
			assign coef[687] =  {12'b101111101001, 12'b100100100001};
			assign coef[688] =  {12'b101111100100, 12'b100100100100};
			assign coef[689] =  {12'b101111011110, 12'b100100100111};
			assign coef[690] =  {12'b101111011001, 12'b100100101011};
			assign coef[691] =  {12'b101111010011, 12'b100100101110};
			assign coef[692] =  {12'b101111001110, 12'b100100110001};
			assign coef[693] =  {12'b101111001001, 12'b100100110101};
			assign coef[694] =  {12'b101111000011, 12'b100100111000};
			assign coef[695] =  {12'b101110111110, 12'b100100111011};
			assign coef[696] =  {12'b101110111001, 12'b100100111111};
			assign coef[697] =  {12'b101110110100, 12'b100101000010};
			assign coef[698] =  {12'b101110101110, 12'b100101000101};
			assign coef[699] =  {12'b101110101001, 12'b100101001001};
			assign coef[700] =  {12'b101110100100, 12'b100101001100};
			assign coef[701] =  {12'b101110011110, 12'b100101010000};
			assign coef[702] =  {12'b101110011001, 12'b100101010011};
			assign coef[703] =  {12'b101110010100, 12'b100101010110};
			assign coef[704] =  {12'b101110001111, 12'b100101011010};
			assign coef[705] =  {12'b101110001001, 12'b100101011101};
			assign coef[706] =  {12'b101110000100, 12'b100101100001};
			assign coef[707] =  {12'b101101111111, 12'b100101100100};
			assign coef[708] =  {12'b101101111010, 12'b100101101000};
			assign coef[709] =  {12'b101101110101, 12'b100101101100};
			assign coef[710] =  {12'b101101110000, 12'b100101101111};
			assign coef[711] =  {12'b101101101010, 12'b100101110011};
			assign coef[712] =  {12'b101101100101, 12'b100101110110};
			assign coef[713] =  {12'b101101100000, 12'b100101111010};
			assign coef[714] =  {12'b101101011011, 12'b100101111110};
			assign coef[715] =  {12'b101101010110, 12'b100110000001};
			assign coef[716] =  {12'b101101010001, 12'b100110000101};
			assign coef[717] =  {12'b101101001100, 12'b100110001001};
			assign coef[718] =  {12'b101101000111, 12'b100110001100};
			assign coef[719] =  {12'b101101000010, 12'b100110010000};
			assign coef[720] =  {12'b101100111101, 12'b100110010100};
			assign coef[721] =  {12'b101100111000, 12'b100110011000};
			assign coef[722] =  {12'b101100110010, 12'b100110011011};
			assign coef[723] =  {12'b101100101101, 12'b100110011111};
			assign coef[724] =  {12'b101100101000, 12'b100110100011};
			assign coef[725] =  {12'b101100100011, 12'b100110100111};
			assign coef[726] =  {12'b101100011110, 12'b100110101011};
			assign coef[727] =  {12'b101100011010, 12'b100110101110};
			assign coef[728] =  {12'b101100010101, 12'b100110110010};
			assign coef[729] =  {12'b101100010000, 12'b100110110110};
			assign coef[730] =  {12'b101100001011, 12'b100110111010};
			assign coef[731] =  {12'b101100000110, 12'b100110111110};
			assign coef[732] =  {12'b101100000001, 12'b100111000010};
			assign coef[733] =  {12'b101011111100, 12'b100111000110};
			assign coef[734] =  {12'b101011110111, 12'b100111001010};
			assign coef[735] =  {12'b101011110010, 12'b100111001110};
			assign coef[736] =  {12'b101011101101, 12'b100111010010};
			assign coef[737] =  {12'b101011101000, 12'b100111010110};
			assign coef[738] =  {12'b101011100100, 12'b100111011010};
			assign coef[739] =  {12'b101011011111, 12'b100111011110};
			assign coef[740] =  {12'b101011011010, 12'b100111100010};
			assign coef[741] =  {12'b101011010101, 12'b100111100110};
			assign coef[742] =  {12'b101011010000, 12'b100111101010};
			assign coef[743] =  {12'b101011001100, 12'b100111101110};
			assign coef[744] =  {12'b101011000111, 12'b100111110010};
			assign coef[745] =  {12'b101011000010, 12'b100111110110};
			assign coef[746] =  {12'b101010111101, 12'b100111111010};
			assign coef[747] =  {12'b101010111001, 12'b100111111110};
			assign coef[748] =  {12'b101010110100, 12'b101000000010};
			assign coef[749] =  {12'b101010101111, 12'b101000000111};
			assign coef[750] =  {12'b101010101011, 12'b101000001011};
			assign coef[751] =  {12'b101010100110, 12'b101000001111};
			assign coef[752] =  {12'b101010100001, 12'b101000010011};
			assign coef[753] =  {12'b101010011101, 12'b101000010111};
			assign coef[754] =  {12'b101010011000, 12'b101000011100};
			assign coef[755] =  {12'b101010010011, 12'b101000100000};
			assign coef[756] =  {12'b101010001111, 12'b101000100100};
			assign coef[757] =  {12'b101010001010, 12'b101000101000};
			assign coef[758] =  {12'b101010000110, 12'b101000101101};
			assign coef[759] =  {12'b101010000001, 12'b101000110001};
			assign coef[760] =  {12'b101001111100, 12'b101000110101};
			assign coef[761] =  {12'b101001111000, 12'b101000111010};
			assign coef[762] =  {12'b101001110011, 12'b101000111110};
			assign coef[763] =  {12'b101001101111, 12'b101001000010};
			assign coef[764] =  {12'b101001101010, 12'b101001000111};
			assign coef[765] =  {12'b101001100110, 12'b101001001011};
			assign coef[766] =  {12'b101001100001, 12'b101001010000};
			assign coef[767] =  {12'b101001011101, 12'b101001010100};
			assign coef[768] =  {12'b101001011001, 12'b101001011001};
			assign coef[769] =  {12'b101001010100, 12'b101001011101};
			assign coef[770] =  {12'b101001010000, 12'b101001100001};
			assign coef[771] =  {12'b101001001011, 12'b101001100110};
			assign coef[772] =  {12'b101001000111, 12'b101001101010};
			assign coef[773] =  {12'b101001000010, 12'b101001101111};
			assign coef[774] =  {12'b101000111110, 12'b101001110011};
			assign coef[775] =  {12'b101000111010, 12'b101001111000};
			assign coef[776] =  {12'b101000110101, 12'b101001111100};
			assign coef[777] =  {12'b101000110001, 12'b101010000001};
			assign coef[778] =  {12'b101000101101, 12'b101010000110};
			assign coef[779] =  {12'b101000101000, 12'b101010001010};
			assign coef[780] =  {12'b101000100100, 12'b101010001111};
			assign coef[781] =  {12'b101000100000, 12'b101010010011};
			assign coef[782] =  {12'b101000011100, 12'b101010011000};
			assign coef[783] =  {12'b101000010111, 12'b101010011101};
			assign coef[784] =  {12'b101000010011, 12'b101010100001};
			assign coef[785] =  {12'b101000001111, 12'b101010100110};
			assign coef[786] =  {12'b101000001011, 12'b101010101011};
			assign coef[787] =  {12'b101000000111, 12'b101010101111};
			assign coef[788] =  {12'b101000000010, 12'b101010110100};
			assign coef[789] =  {12'b100111111110, 12'b101010111001};
			assign coef[790] =  {12'b100111111010, 12'b101010111101};
			assign coef[791] =  {12'b100111110110, 12'b101011000010};
			assign coef[792] =  {12'b100111110010, 12'b101011000111};
			assign coef[793] =  {12'b100111101110, 12'b101011001100};
			assign coef[794] =  {12'b100111101010, 12'b101011010000};
			assign coef[795] =  {12'b100111100110, 12'b101011010101};
			assign coef[796] =  {12'b100111100010, 12'b101011011010};
			assign coef[797] =  {12'b100111011110, 12'b101011011111};
			assign coef[798] =  {12'b100111011010, 12'b101011100100};
			assign coef[799] =  {12'b100111010110, 12'b101011101000};
			assign coef[800] =  {12'b100111010010, 12'b101011101101};
			assign coef[801] =  {12'b100111001110, 12'b101011110010};
			assign coef[802] =  {12'b100111001010, 12'b101011110111};
			assign coef[803] =  {12'b100111000110, 12'b101011111100};
			assign coef[804] =  {12'b100111000010, 12'b101100000001};
			assign coef[805] =  {12'b100110111110, 12'b101100000110};
			assign coef[806] =  {12'b100110111010, 12'b101100001011};
			assign coef[807] =  {12'b100110110110, 12'b101100010000};
			assign coef[808] =  {12'b100110110010, 12'b101100010101};
			assign coef[809] =  {12'b100110101110, 12'b101100011010};
			assign coef[810] =  {12'b100110101011, 12'b101100011110};
			assign coef[811] =  {12'b100110100111, 12'b101100100011};
			assign coef[812] =  {12'b100110100011, 12'b101100101000};
			assign coef[813] =  {12'b100110011111, 12'b101100101101};
			assign coef[814] =  {12'b100110011011, 12'b101100110010};
			assign coef[815] =  {12'b100110011000, 12'b101100111000};
			assign coef[816] =  {12'b100110010100, 12'b101100111101};
			assign coef[817] =  {12'b100110010000, 12'b101101000010};
			assign coef[818] =  {12'b100110001100, 12'b101101000111};
			assign coef[819] =  {12'b100110001001, 12'b101101001100};
			assign coef[820] =  {12'b100110000101, 12'b101101010001};
			assign coef[821] =  {12'b100110000001, 12'b101101010110};
			assign coef[822] =  {12'b100101111110, 12'b101101011011};
			assign coef[823] =  {12'b100101111010, 12'b101101100000};
			assign coef[824] =  {12'b100101110110, 12'b101101100101};
			assign coef[825] =  {12'b100101110011, 12'b101101101010};
			assign coef[826] =  {12'b100101101111, 12'b101101110000};
			assign coef[827] =  {12'b100101101100, 12'b101101110101};
			assign coef[828] =  {12'b100101101000, 12'b101101111010};
			assign coef[829] =  {12'b100101100100, 12'b101101111111};
			assign coef[830] =  {12'b100101100001, 12'b101110000100};
			assign coef[831] =  {12'b100101011101, 12'b101110001001};
			assign coef[832] =  {12'b100101011010, 12'b101110001111};
			assign coef[833] =  {12'b100101010110, 12'b101110010100};
			assign coef[834] =  {12'b100101010011, 12'b101110011001};
			assign coef[835] =  {12'b100101010000, 12'b101110011110};
			assign coef[836] =  {12'b100101001100, 12'b101110100100};
			assign coef[837] =  {12'b100101001001, 12'b101110101001};
			assign coef[838] =  {12'b100101000101, 12'b101110101110};
			assign coef[839] =  {12'b100101000010, 12'b101110110100};
			assign coef[840] =  {12'b100100111111, 12'b101110111001};
			assign coef[841] =  {12'b100100111011, 12'b101110111110};
			assign coef[842] =  {12'b100100111000, 12'b101111000011};
			assign coef[843] =  {12'b100100110101, 12'b101111001001};
			assign coef[844] =  {12'b100100110001, 12'b101111001110};
			assign coef[845] =  {12'b100100101110, 12'b101111010011};
			assign coef[846] =  {12'b100100101011, 12'b101111011001};
			assign coef[847] =  {12'b100100100111, 12'b101111011110};
			assign coef[848] =  {12'b100100100100, 12'b101111100100};
			assign coef[849] =  {12'b100100100001, 12'b101111101001};
			assign coef[850] =  {12'b100100011110, 12'b101111101110};
			assign coef[851] =  {12'b100100011011, 12'b101111110100};
			assign coef[852] =  {12'b100100010111, 12'b101111111001};
			assign coef[853] =  {12'b100100010100, 12'b101111111111};
			assign coef[854] =  {12'b100100010001, 12'b110000000100};
			assign coef[855] =  {12'b100100001110, 12'b110000001010};
			assign coef[856] =  {12'b100100001011, 12'b110000001111};
			assign coef[857] =  {12'b100100001000, 12'b110000010100};
			assign coef[858] =  {12'b100100000101, 12'b110000011010};
			assign coef[859] =  {12'b100100000010, 12'b110000011111};
			assign coef[860] =  {12'b100011111111, 12'b110000100101};
			assign coef[861] =  {12'b100011111100, 12'b110000101010};
			assign coef[862] =  {12'b100011111001, 12'b110000110000};
			assign coef[863] =  {12'b100011110110, 12'b110000110101};
			assign coef[864] =  {12'b100011110011, 12'b110000111011};
			assign coef[865] =  {12'b100011110000, 12'b110001000001};
			assign coef[866] =  {12'b100011101101, 12'b110001000110};
			assign coef[867] =  {12'b100011101010, 12'b110001001100};
			assign coef[868] =  {12'b100011100111, 12'b110001010001};
			assign coef[869] =  {12'b100011100100, 12'b110001010111};
			assign coef[870] =  {12'b100011100001, 12'b110001011100};
			assign coef[871] =  {12'b100011011110, 12'b110001100010};
			assign coef[872] =  {12'b100011011100, 12'b110001101000};
			assign coef[873] =  {12'b100011011001, 12'b110001101101};
			assign coef[874] =  {12'b100011010110, 12'b110001110011};
			assign coef[875] =  {12'b100011010011, 12'b110001111000};
			assign coef[876] =  {12'b100011010000, 12'b110001111110};
			assign coef[877] =  {12'b100011001110, 12'b110010000100};
			assign coef[878] =  {12'b100011001011, 12'b110010001001};
			assign coef[879] =  {12'b100011001000, 12'b110010001111};
			assign coef[880] =  {12'b100011000101, 12'b110010010101};
			assign coef[881] =  {12'b100011000011, 12'b110010011010};
			assign coef[882] =  {12'b100011000000, 12'b110010100000};
			assign coef[883] =  {12'b100010111110, 12'b110010100110};
			assign coef[884] =  {12'b100010111011, 12'b110010101100};
			assign coef[885] =  {12'b100010111000, 12'b110010110001};
			assign coef[886] =  {12'b100010110110, 12'b110010110111};
			assign coef[887] =  {12'b100010110011, 12'b110010111101};
			assign coef[888] =  {12'b100010110001, 12'b110011000010};
			assign coef[889] =  {12'b100010101110, 12'b110011001000};
			assign coef[890] =  {12'b100010101100, 12'b110011001110};
			assign coef[891] =  {12'b100010101001, 12'b110011010100};
			assign coef[892] =  {12'b100010100111, 12'b110011011001};
			assign coef[893] =  {12'b100010100100, 12'b110011011111};
			assign coef[894] =  {12'b100010100010, 12'b110011100101};
			assign coef[895] =  {12'b100010011111, 12'b110011101011};
			assign coef[896] =  {12'b100010011101, 12'b110011110001};
			assign coef[897] =  {12'b100010011010, 12'b110011110110};
			assign coef[898] =  {12'b100010011000, 12'b110011111100};
			assign coef[899] =  {12'b100010010110, 12'b110100000010};
			assign coef[900] =  {12'b100010010011, 12'b110100001000};
			assign coef[901] =  {12'b100010010001, 12'b110100001110};
			assign coef[902] =  {12'b100010001111, 12'b110100010100};
			assign coef[903] =  {12'b100010001100, 12'b110100011001};
			assign coef[904] =  {12'b100010001010, 12'b110100011111};
			assign coef[905] =  {12'b100010001000, 12'b110100100101};
			assign coef[906] =  {12'b100010000110, 12'b110100101011};
			assign coef[907] =  {12'b100010000011, 12'b110100110001};
			assign coef[908] =  {12'b100010000001, 12'b110100110111};
			assign coef[909] =  {12'b100001111111, 12'b110100111101};
			assign coef[910] =  {12'b100001111101, 12'b110101000011};
			assign coef[911] =  {12'b100001111011, 12'b110101001000};
			assign coef[912] =  {12'b100001111001, 12'b110101001110};
			assign coef[913] =  {12'b100001110111, 12'b110101010100};
			assign coef[914] =  {12'b100001110100, 12'b110101011010};
			assign coef[915] =  {12'b100001110010, 12'b110101100000};
			assign coef[916] =  {12'b100001110000, 12'b110101100110};
			assign coef[917] =  {12'b100001101110, 12'b110101101100};
			assign coef[918] =  {12'b100001101100, 12'b110101110010};
			assign coef[919] =  {12'b100001101010, 12'b110101111000};
			assign coef[920] =  {12'b100001101000, 12'b110101111110};
			assign coef[921] =  {12'b100001100110, 12'b110110000100};
			assign coef[922] =  {12'b100001100100, 12'b110110001010};
			assign coef[923] =  {12'b100001100010, 12'b110110010000};
			assign coef[924] =  {12'b100001100001, 12'b110110010110};
			assign coef[925] =  {12'b100001011111, 12'b110110011100};
			assign coef[926] =  {12'b100001011101, 12'b110110100010};
			assign coef[927] =  {12'b100001011011, 12'b110110101000};
			assign coef[928] =  {12'b100001011001, 12'b110110101110};
			assign coef[929] =  {12'b100001010111, 12'b110110110100};
			assign coef[930] =  {12'b100001010101, 12'b110110111010};
			assign coef[931] =  {12'b100001010100, 12'b110111000000};
			assign coef[932] =  {12'b100001010010, 12'b110111000110};
			assign coef[933] =  {12'b100001010000, 12'b110111001100};
			assign coef[934] =  {12'b100001001110, 12'b110111010010};
			assign coef[935] =  {12'b100001001101, 12'b110111011000};
			assign coef[936] =  {12'b100001001011, 12'b110111011110};
			assign coef[937] =  {12'b100001001001, 12'b110111100100};
			assign coef[938] =  {12'b100001001000, 12'b110111101010};
			assign coef[939] =  {12'b100001000110, 12'b110111110000};
			assign coef[940] =  {12'b100001000101, 12'b110111110110};
			assign coef[941] =  {12'b100001000011, 12'b110111111100};
			assign coef[942] =  {12'b100001000001, 12'b111000000010};
			assign coef[943] =  {12'b100001000000, 12'b111000001000};
			assign coef[944] =  {12'b100000111110, 12'b111000001111};
			assign coef[945] =  {12'b100000111101, 12'b111000010101};
			assign coef[946] =  {12'b100000111011, 12'b111000011011};
			assign coef[947] =  {12'b100000111010, 12'b111000100001};
			assign coef[948] =  {12'b100000111000, 12'b111000100111};
			assign coef[949] =  {12'b100000110111, 12'b111000101101};
			assign coef[950] =  {12'b100000110101, 12'b111000110011};
			assign coef[951] =  {12'b100000110100, 12'b111000111001};
			assign coef[952] =  {12'b100000110011, 12'b111000111111};
			assign coef[953] =  {12'b100000110001, 12'b111001000110};
			assign coef[954] =  {12'b100000110000, 12'b111001001100};
			assign coef[955] =  {12'b100000101111, 12'b111001010010};
			assign coef[956] =  {12'b100000101101, 12'b111001011000};
			assign coef[957] =  {12'b100000101100, 12'b111001011110};
			assign coef[958] =  {12'b100000101011, 12'b111001100100};
			assign coef[959] =  {12'b100000101010, 12'b111001101010};
			assign coef[960] =  {12'b100000101000, 12'b111001110001};
			assign coef[961] =  {12'b100000100111, 12'b111001110111};
			assign coef[962] =  {12'b100000100110, 12'b111001111101};
			assign coef[963] =  {12'b100000100101, 12'b111010000011};
			assign coef[964] =  {12'b100000100100, 12'b111010001001};
			assign coef[965] =  {12'b100000100010, 12'b111010001111};
			assign coef[966] =  {12'b100000100001, 12'b111010010110};
			assign coef[967] =  {12'b100000100000, 12'b111010011100};
			assign coef[968] =  {12'b100000011111, 12'b111010100010};
			assign coef[969] =  {12'b100000011110, 12'b111010101000};
			assign coef[970] =  {12'b100000011101, 12'b111010101110};
			assign coef[971] =  {12'b100000011100, 12'b111010110101};
			assign coef[972] =  {12'b100000011011, 12'b111010111011};
			assign coef[973] =  {12'b100000011010, 12'b111011000001};
			assign coef[974] =  {12'b100000011001, 12'b111011000111};
			assign coef[975] =  {12'b100000011000, 12'b111011001101};
			assign coef[976] =  {12'b100000010111, 12'b111011010100};
			assign coef[977] =  {12'b100000010110, 12'b111011011010};
			assign coef[978] =  {12'b100000010101, 12'b111011100000};
			assign coef[979] =  {12'b100000010100, 12'b111011100110};
			assign coef[980] =  {12'b100000010100, 12'b111011101100};
			assign coef[981] =  {12'b100000010011, 12'b111011110011};
			assign coef[982] =  {12'b100000010010, 12'b111011111001};
			assign coef[983] =  {12'b100000010001, 12'b111011111111};
			assign coef[984] =  {12'b100000010000, 12'b111100000101};
			assign coef[985] =  {12'b100000010000, 12'b111100001100};
			assign coef[986] =  {12'b100000001111, 12'b111100010010};
			assign coef[987] =  {12'b100000001110, 12'b111100011000};
			assign coef[988] =  {12'b100000001101, 12'b111100011110};
			assign coef[989] =  {12'b100000001101, 12'b111100100101};
			assign coef[990] =  {12'b100000001100, 12'b111100101011};
			assign coef[991] =  {12'b100000001011, 12'b111100110001};
			assign coef[992] =  {12'b100000001011, 12'b111100110111};
			assign coef[993] =  {12'b100000001010, 12'b111100111110};
			assign coef[994] =  {12'b100000001010, 12'b111101000100};
			assign coef[995] =  {12'b100000001001, 12'b111101001010};
			assign coef[996] =  {12'b100000001000, 12'b111101010000};
			assign coef[997] =  {12'b100000001000, 12'b111101010111};
			assign coef[998] =  {12'b100000000111, 12'b111101011101};
			assign coef[999] =  {12'b100000000111, 12'b111101100011};
			assign coef[1000] = {12'b100000000110, 12'b111101101001};
			assign coef[1001] = {12'b100000000110, 12'b111101110000};
			assign coef[1002] = {12'b100000000110, 12'b111101110110};
			assign coef[1003] = {12'b100000000101, 12'b111101111100};
			assign coef[1004] = {12'b100000000101, 12'b111110000010};
			assign coef[1005] = {12'b100000000100, 12'b111110001001};
			assign coef[1006] = {12'b100000000100, 12'b111110001111};
			assign coef[1007] = {12'b100000000100, 12'b111110010101};
			assign coef[1008] = {12'b100000000011, 12'b111110011100};
			assign coef[1009] = {12'b100000000011, 12'b111110100010};
			assign coef[1010] = {12'b100000000011, 12'b111110101000};
			assign coef[1011] = {12'b100000000011, 12'b111110101110};
			assign coef[1012] = {12'b100000000010, 12'b111110110101};
			assign coef[1013] = {12'b100000000010, 12'b111110111011};
			assign coef[1014] = {12'b100000000010, 12'b111111000001};
			assign coef[1015] = {12'b100000000010, 12'b111111000111};
			assign coef[1016] = {12'b100000000010, 12'b111111001110};
			assign coef[1017] = {12'b100000000001, 12'b111111010100};
			assign coef[1018] = {12'b100000000001, 12'b111111011010};
			assign coef[1019] = {12'b100000000001, 12'b111111100001};
			assign coef[1020] = {12'b100000000001, 12'b111111100111};
			assign coef[1021] = {12'b100000000001, 12'b111111101101};
			assign coef[1022] = {12'b100000000001, 12'b111111110011};
			assign coef[1023] = {12'b100000000001, 12'b111111111010};

		//--- fifo stage
			localparam depth=`LOG2(size);
			fifo #(.depth(depth)) inst_fifo(.clk(clk), .rst(rst), .stall_in(stall), .stall_out(stall_out));

			assign comb_stall = stall_out & stall;

		//--- input stage
			always @(posedge clk or posedge rst) begin
				if (rst) begin
					a0_wr[0]       <= 0;                           
					a0_wr[1]       <= 0;                           
					a0_wr[2]       <= 0;                           
					a0_wr[3]       <= 0;                           
					a0_wr[4]       <= 0;                           
					a0_wr[5]       <= 0;                           
					a0_wr[6]       <= 0;                           
					a0_wr[7]       <= 0;                           
					a0_wr[8]       <= 0;                           
					a0_wr[9]       <= 0;                           
					a0_wr[10]      <= 0;                           
					a0_wr[11]      <= 0;                           
					a0_wr[12]      <= 0;                           
					a0_wr[13]      <= 0;                           
					a0_wr[14]      <= 0;                           
					a0_wr[15]      <= 0;                           
					a0_wr[16]      <= 0;                           
					a0_wr[17]      <= 0;                           
					a0_wr[18]      <= 0;                           
					a0_wr[19]      <= 0;                           
					a0_wr[20]      <= 0;                           
					a0_wr[21]      <= 0;                           
					a0_wr[22]      <= 0;                           
					a0_wr[23]      <= 0;                           
					a0_wr[24]      <= 0;                           
					a0_wr[25]      <= 0;                           
					a0_wr[26]      <= 0;                           
					a0_wr[27]      <= 0;                           
					a0_wr[28]      <= 0;                           
					a0_wr[29]      <= 0;                           
					a0_wr[30]      <= 0;                           
					a0_wr[31]      <= 0;                           
					a0_wr[32]      <= 0;                           
					a0_wr[33]      <= 0;                           
					a0_wr[34]      <= 0;                           
					a0_wr[35]      <= 0;                           
					a0_wr[36]      <= 0;                           
					a0_wr[37]      <= 0;                           
					a0_wr[38]      <= 0;                           
					a0_wr[39]      <= 0;                           
					a0_wr[40]      <= 0;                           
					a0_wr[41]      <= 0;                           
					a0_wr[42]      <= 0;                           
					a0_wr[43]      <= 0;                           
					a0_wr[44]      <= 0;                           
					a0_wr[45]      <= 0;                           
					a0_wr[46]      <= 0;                           
					a0_wr[47]      <= 0;                           
					a0_wr[48]      <= 0;                           
					a0_wr[49]      <= 0;                           
					a0_wr[50]      <= 0;                           
					a0_wr[51]      <= 0;                           
					a0_wr[52]      <= 0;                           
					a0_wr[53]      <= 0;                           
					a0_wr[54]      <= 0;                           
					a0_wr[55]      <= 0;                           
					a0_wr[56]      <= 0;                           
					a0_wr[57]      <= 0;                           
					a0_wr[58]      <= 0;                           
					a0_wr[59]      <= 0;                           
					a0_wr[60]      <= 0;                           
					a0_wr[61]      <= 0;                           
					a0_wr[62]      <= 0;                           
					a0_wr[63]      <= 0;                           
					a0_wr[64]      <= 0;                           
					a0_wr[65]      <= 0;                           
					a0_wr[66]      <= 0;                           
					a0_wr[67]      <= 0;                           
					a0_wr[68]      <= 0;                           
					a0_wr[69]      <= 0;                           
					a0_wr[70]      <= 0;                           
					a0_wr[71]      <= 0;                           
					a0_wr[72]      <= 0;                           
					a0_wr[73]      <= 0;                           
					a0_wr[74]      <= 0;                           
					a0_wr[75]      <= 0;                           
					a0_wr[76]      <= 0;                           
					a0_wr[77]      <= 0;                           
					a0_wr[78]      <= 0;                           
					a0_wr[79]      <= 0;                           
					a0_wr[80]      <= 0;                           
					a0_wr[81]      <= 0;                           
					a0_wr[82]      <= 0;                           
					a0_wr[83]      <= 0;                           
					a0_wr[84]      <= 0;                           
					a0_wr[85]      <= 0;                           
					a0_wr[86]      <= 0;                           
					a0_wr[87]      <= 0;                           
					a0_wr[88]      <= 0;                           
					a0_wr[89]      <= 0;                           
					a0_wr[90]      <= 0;                           
					a0_wr[91]      <= 0;                           
					a0_wr[92]      <= 0;                           
					a0_wr[93]      <= 0;                           
					a0_wr[94]      <= 0;                           
					a0_wr[95]      <= 0;                           
					a0_wr[96]      <= 0;                           
					a0_wr[97]      <= 0;                           
					a0_wr[98]      <= 0;                           
					a0_wr[99]      <= 0;                           
					a0_wr[100]     <= 0;                           
					a0_wr[101]     <= 0;                           
					a0_wr[102]     <= 0;                           
					a0_wr[103]     <= 0;                           
					a0_wr[104]     <= 0;                           
					a0_wr[105]     <= 0;                           
					a0_wr[106]     <= 0;                           
					a0_wr[107]     <= 0;                           
					a0_wr[108]     <= 0;                           
					a0_wr[109]     <= 0;                           
					a0_wr[110]     <= 0;                           
					a0_wr[111]     <= 0;                           
					a0_wr[112]     <= 0;                           
					a0_wr[113]     <= 0;                           
					a0_wr[114]     <= 0;                           
					a0_wr[115]     <= 0;                           
					a0_wr[116]     <= 0;                           
					a0_wr[117]     <= 0;                           
					a0_wr[118]     <= 0;                           
					a0_wr[119]     <= 0;                           
					a0_wr[120]     <= 0;                           
					a0_wr[121]     <= 0;                           
					a0_wr[122]     <= 0;                           
					a0_wr[123]     <= 0;                           
					a0_wr[124]     <= 0;                           
					a0_wr[125]     <= 0;                           
					a0_wr[126]     <= 0;                           
					a0_wr[127]     <= 0;                           
					a0_wr[128]     <= 0;                           
					a0_wr[129]     <= 0;                           
					a0_wr[130]     <= 0;                           
					a0_wr[131]     <= 0;                           
					a0_wr[132]     <= 0;                           
					a0_wr[133]     <= 0;                           
					a0_wr[134]     <= 0;                           
					a0_wr[135]     <= 0;                           
					a0_wr[136]     <= 0;                           
					a0_wr[137]     <= 0;                           
					a0_wr[138]     <= 0;                           
					a0_wr[139]     <= 0;                           
					a0_wr[140]     <= 0;                           
					a0_wr[141]     <= 0;                           
					a0_wr[142]     <= 0;                           
					a0_wr[143]     <= 0;                           
					a0_wr[144]     <= 0;                           
					a0_wr[145]     <= 0;                           
					a0_wr[146]     <= 0;                           
					a0_wr[147]     <= 0;                           
					a0_wr[148]     <= 0;                           
					a0_wr[149]     <= 0;                           
					a0_wr[150]     <= 0;                           
					a0_wr[151]     <= 0;                           
					a0_wr[152]     <= 0;                           
					a0_wr[153]     <= 0;                           
					a0_wr[154]     <= 0;                           
					a0_wr[155]     <= 0;                           
					a0_wr[156]     <= 0;                           
					a0_wr[157]     <= 0;                           
					a0_wr[158]     <= 0;                           
					a0_wr[159]     <= 0;                           
					a0_wr[160]     <= 0;                           
					a0_wr[161]     <= 0;                           
					a0_wr[162]     <= 0;                           
					a0_wr[163]     <= 0;                           
					a0_wr[164]     <= 0;                           
					a0_wr[165]     <= 0;                           
					a0_wr[166]     <= 0;                           
					a0_wr[167]     <= 0;                           
					a0_wr[168]     <= 0;                           
					a0_wr[169]     <= 0;                           
					a0_wr[170]     <= 0;                           
					a0_wr[171]     <= 0;                           
					a0_wr[172]     <= 0;                           
					a0_wr[173]     <= 0;                           
					a0_wr[174]     <= 0;                           
					a0_wr[175]     <= 0;                           
					a0_wr[176]     <= 0;                           
					a0_wr[177]     <= 0;                           
					a0_wr[178]     <= 0;                           
					a0_wr[179]     <= 0;                           
					a0_wr[180]     <= 0;                           
					a0_wr[181]     <= 0;                           
					a0_wr[182]     <= 0;                           
					a0_wr[183]     <= 0;                           
					a0_wr[184]     <= 0;                           
					a0_wr[185]     <= 0;                           
					a0_wr[186]     <= 0;                           
					a0_wr[187]     <= 0;                           
					a0_wr[188]     <= 0;                           
					a0_wr[189]     <= 0;                           
					a0_wr[190]     <= 0;                           
					a0_wr[191]     <= 0;                           
					a0_wr[192]     <= 0;                           
					a0_wr[193]     <= 0;                           
					a0_wr[194]     <= 0;                           
					a0_wr[195]     <= 0;                           
					a0_wr[196]     <= 0;                           
					a0_wr[197]     <= 0;                           
					a0_wr[198]     <= 0;                           
					a0_wr[199]     <= 0;                           
					a0_wr[200]     <= 0;                           
					a0_wr[201]     <= 0;                           
					a0_wr[202]     <= 0;                           
					a0_wr[203]     <= 0;                           
					a0_wr[204]     <= 0;                           
					a0_wr[205]     <= 0;                           
					a0_wr[206]     <= 0;                           
					a0_wr[207]     <= 0;                           
					a0_wr[208]     <= 0;                           
					a0_wr[209]     <= 0;                           
					a0_wr[210]     <= 0;                           
					a0_wr[211]     <= 0;                           
					a0_wr[212]     <= 0;                           
					a0_wr[213]     <= 0;                           
					a0_wr[214]     <= 0;                           
					a0_wr[215]     <= 0;                           
					a0_wr[216]     <= 0;                           
					a0_wr[217]     <= 0;                           
					a0_wr[218]     <= 0;                           
					a0_wr[219]     <= 0;                           
					a0_wr[220]     <= 0;                           
					a0_wr[221]     <= 0;                           
					a0_wr[222]     <= 0;                           
					a0_wr[223]     <= 0;                           
					a0_wr[224]     <= 0;                           
					a0_wr[225]     <= 0;                           
					a0_wr[226]     <= 0;                           
					a0_wr[227]     <= 0;                           
					a0_wr[228]     <= 0;                           
					a0_wr[229]     <= 0;                           
					a0_wr[230]     <= 0;                           
					a0_wr[231]     <= 0;                           
					a0_wr[232]     <= 0;                           
					a0_wr[233]     <= 0;                           
					a0_wr[234]     <= 0;                           
					a0_wr[235]     <= 0;                           
					a0_wr[236]     <= 0;                           
					a0_wr[237]     <= 0;                           
					a0_wr[238]     <= 0;                           
					a0_wr[239]     <= 0;                           
					a0_wr[240]     <= 0;                           
					a0_wr[241]     <= 0;                           
					a0_wr[242]     <= 0;                           
					a0_wr[243]     <= 0;                           
					a0_wr[244]     <= 0;                           
					a0_wr[245]     <= 0;                           
					a0_wr[246]     <= 0;                           
					a0_wr[247]     <= 0;                           
					a0_wr[248]     <= 0;                           
					a0_wr[249]     <= 0;                           
					a0_wr[250]     <= 0;                           
					a0_wr[251]     <= 0;                           
					a0_wr[252]     <= 0;                           
					a0_wr[253]     <= 0;                           
					a0_wr[254]     <= 0;                           
					a0_wr[255]     <= 0;                           
					a0_wr[256]     <= 0;                           
					a0_wr[257]     <= 0;                           
					a0_wr[258]     <= 0;                           
					a0_wr[259]     <= 0;                           
					a0_wr[260]     <= 0;                           
					a0_wr[261]     <= 0;                           
					a0_wr[262]     <= 0;                           
					a0_wr[263]     <= 0;                           
					a0_wr[264]     <= 0;                           
					a0_wr[265]     <= 0;                           
					a0_wr[266]     <= 0;                           
					a0_wr[267]     <= 0;                           
					a0_wr[268]     <= 0;                           
					a0_wr[269]     <= 0;                           
					a0_wr[270]     <= 0;                           
					a0_wr[271]     <= 0;                           
					a0_wr[272]     <= 0;                           
					a0_wr[273]     <= 0;                           
					a0_wr[274]     <= 0;                           
					a0_wr[275]     <= 0;                           
					a0_wr[276]     <= 0;                           
					a0_wr[277]     <= 0;                           
					a0_wr[278]     <= 0;                           
					a0_wr[279]     <= 0;                           
					a0_wr[280]     <= 0;                           
					a0_wr[281]     <= 0;                           
					a0_wr[282]     <= 0;                           
					a0_wr[283]     <= 0;                           
					a0_wr[284]     <= 0;                           
					a0_wr[285]     <= 0;                           
					a0_wr[286]     <= 0;                           
					a0_wr[287]     <= 0;                           
					a0_wr[288]     <= 0;                           
					a0_wr[289]     <= 0;                           
					a0_wr[290]     <= 0;                           
					a0_wr[291]     <= 0;                           
					a0_wr[292]     <= 0;                           
					a0_wr[293]     <= 0;                           
					a0_wr[294]     <= 0;                           
					a0_wr[295]     <= 0;                           
					a0_wr[296]     <= 0;                           
					a0_wr[297]     <= 0;                           
					a0_wr[298]     <= 0;                           
					a0_wr[299]     <= 0;                           
					a0_wr[300]     <= 0;                           
					a0_wr[301]     <= 0;                           
					a0_wr[302]     <= 0;                           
					a0_wr[303]     <= 0;                           
					a0_wr[304]     <= 0;                           
					a0_wr[305]     <= 0;                           
					a0_wr[306]     <= 0;                           
					a0_wr[307]     <= 0;                           
					a0_wr[308]     <= 0;                           
					a0_wr[309]     <= 0;                           
					a0_wr[310]     <= 0;                           
					a0_wr[311]     <= 0;                           
					a0_wr[312]     <= 0;                           
					a0_wr[313]     <= 0;                           
					a0_wr[314]     <= 0;                           
					a0_wr[315]     <= 0;                           
					a0_wr[316]     <= 0;                           
					a0_wr[317]     <= 0;                           
					a0_wr[318]     <= 0;                           
					a0_wr[319]     <= 0;                           
					a0_wr[320]     <= 0;                           
					a0_wr[321]     <= 0;                           
					a0_wr[322]     <= 0;                           
					a0_wr[323]     <= 0;                           
					a0_wr[324]     <= 0;                           
					a0_wr[325]     <= 0;                           
					a0_wr[326]     <= 0;                           
					a0_wr[327]     <= 0;                           
					a0_wr[328]     <= 0;                           
					a0_wr[329]     <= 0;                           
					a0_wr[330]     <= 0;                           
					a0_wr[331]     <= 0;                           
					a0_wr[332]     <= 0;                           
					a0_wr[333]     <= 0;                           
					a0_wr[334]     <= 0;                           
					a0_wr[335]     <= 0;                           
					a0_wr[336]     <= 0;                           
					a0_wr[337]     <= 0;                           
					a0_wr[338]     <= 0;                           
					a0_wr[339]     <= 0;                           
					a0_wr[340]     <= 0;                           
					a0_wr[341]     <= 0;                           
					a0_wr[342]     <= 0;                           
					a0_wr[343]     <= 0;                           
					a0_wr[344]     <= 0;                           
					a0_wr[345]     <= 0;                           
					a0_wr[346]     <= 0;                           
					a0_wr[347]     <= 0;                           
					a0_wr[348]     <= 0;                           
					a0_wr[349]     <= 0;                           
					a0_wr[350]     <= 0;                           
					a0_wr[351]     <= 0;                           
					a0_wr[352]     <= 0;                           
					a0_wr[353]     <= 0;                           
					a0_wr[354]     <= 0;                           
					a0_wr[355]     <= 0;                           
					a0_wr[356]     <= 0;                           
					a0_wr[357]     <= 0;                           
					a0_wr[358]     <= 0;                           
					a0_wr[359]     <= 0;                           
					a0_wr[360]     <= 0;                           
					a0_wr[361]     <= 0;                           
					a0_wr[362]     <= 0;                           
					a0_wr[363]     <= 0;                           
					a0_wr[364]     <= 0;                           
					a0_wr[365]     <= 0;                           
					a0_wr[366]     <= 0;                           
					a0_wr[367]     <= 0;                           
					a0_wr[368]     <= 0;                           
					a0_wr[369]     <= 0;                           
					a0_wr[370]     <= 0;                           
					a0_wr[371]     <= 0;                           
					a0_wr[372]     <= 0;                           
					a0_wr[373]     <= 0;                           
					a0_wr[374]     <= 0;                           
					a0_wr[375]     <= 0;                           
					a0_wr[376]     <= 0;                           
					a0_wr[377]     <= 0;                           
					a0_wr[378]     <= 0;                           
					a0_wr[379]     <= 0;                           
					a0_wr[380]     <= 0;                           
					a0_wr[381]     <= 0;                           
					a0_wr[382]     <= 0;                           
					a0_wr[383]     <= 0;                           
					a0_wr[384]     <= 0;                           
					a0_wr[385]     <= 0;                           
					a0_wr[386]     <= 0;                           
					a0_wr[387]     <= 0;                           
					a0_wr[388]     <= 0;                           
					a0_wr[389]     <= 0;                           
					a0_wr[390]     <= 0;                           
					a0_wr[391]     <= 0;                           
					a0_wr[392]     <= 0;                           
					a0_wr[393]     <= 0;                           
					a0_wr[394]     <= 0;                           
					a0_wr[395]     <= 0;                           
					a0_wr[396]     <= 0;                           
					a0_wr[397]     <= 0;                           
					a0_wr[398]     <= 0;                           
					a0_wr[399]     <= 0;                           
					a0_wr[400]     <= 0;                           
					a0_wr[401]     <= 0;                           
					a0_wr[402]     <= 0;                           
					a0_wr[403]     <= 0;                           
					a0_wr[404]     <= 0;                           
					a0_wr[405]     <= 0;                           
					a0_wr[406]     <= 0;                           
					a0_wr[407]     <= 0;                           
					a0_wr[408]     <= 0;                           
					a0_wr[409]     <= 0;                           
					a0_wr[410]     <= 0;                           
					a0_wr[411]     <= 0;                           
					a0_wr[412]     <= 0;                           
					a0_wr[413]     <= 0;                           
					a0_wr[414]     <= 0;                           
					a0_wr[415]     <= 0;                           
					a0_wr[416]     <= 0;                           
					a0_wr[417]     <= 0;                           
					a0_wr[418]     <= 0;                           
					a0_wr[419]     <= 0;                           
					a0_wr[420]     <= 0;                           
					a0_wr[421]     <= 0;                           
					a0_wr[422]     <= 0;                           
					a0_wr[423]     <= 0;                           
					a0_wr[424]     <= 0;                           
					a0_wr[425]     <= 0;                           
					a0_wr[426]     <= 0;                           
					a0_wr[427]     <= 0;                           
					a0_wr[428]     <= 0;                           
					a0_wr[429]     <= 0;                           
					a0_wr[430]     <= 0;                           
					a0_wr[431]     <= 0;                           
					a0_wr[432]     <= 0;                           
					a0_wr[433]     <= 0;                           
					a0_wr[434]     <= 0;                           
					a0_wr[435]     <= 0;                           
					a0_wr[436]     <= 0;                           
					a0_wr[437]     <= 0;                           
					a0_wr[438]     <= 0;                           
					a0_wr[439]     <= 0;                           
					a0_wr[440]     <= 0;                           
					a0_wr[441]     <= 0;                           
					a0_wr[442]     <= 0;                           
					a0_wr[443]     <= 0;                           
					a0_wr[444]     <= 0;                           
					a0_wr[445]     <= 0;                           
					a0_wr[446]     <= 0;                           
					a0_wr[447]     <= 0;                           
					a0_wr[448]     <= 0;                           
					a0_wr[449]     <= 0;                           
					a0_wr[450]     <= 0;                           
					a0_wr[451]     <= 0;                           
					a0_wr[452]     <= 0;                           
					a0_wr[453]     <= 0;                           
					a0_wr[454]     <= 0;                           
					a0_wr[455]     <= 0;                           
					a0_wr[456]     <= 0;                           
					a0_wr[457]     <= 0;                           
					a0_wr[458]     <= 0;                           
					a0_wr[459]     <= 0;                           
					a0_wr[460]     <= 0;                           
					a0_wr[461]     <= 0;                           
					a0_wr[462]     <= 0;                           
					a0_wr[463]     <= 0;                           
					a0_wr[464]     <= 0;                           
					a0_wr[465]     <= 0;                           
					a0_wr[466]     <= 0;                           
					a0_wr[467]     <= 0;                           
					a0_wr[468]     <= 0;                           
					a0_wr[469]     <= 0;                           
					a0_wr[470]     <= 0;                           
					a0_wr[471]     <= 0;                           
					a0_wr[472]     <= 0;                           
					a0_wr[473]     <= 0;                           
					a0_wr[474]     <= 0;                           
					a0_wr[475]     <= 0;                           
					a0_wr[476]     <= 0;                           
					a0_wr[477]     <= 0;                           
					a0_wr[478]     <= 0;                           
					a0_wr[479]     <= 0;                           
					a0_wr[480]     <= 0;                           
					a0_wr[481]     <= 0;                           
					a0_wr[482]     <= 0;                           
					a0_wr[483]     <= 0;                           
					a0_wr[484]     <= 0;                           
					a0_wr[485]     <= 0;                           
					a0_wr[486]     <= 0;                           
					a0_wr[487]     <= 0;                           
					a0_wr[488]     <= 0;                           
					a0_wr[489]     <= 0;                           
					a0_wr[490]     <= 0;                           
					a0_wr[491]     <= 0;                           
					a0_wr[492]     <= 0;                           
					a0_wr[493]     <= 0;                           
					a0_wr[494]     <= 0;                           
					a0_wr[495]     <= 0;                           
					a0_wr[496]     <= 0;                           
					a0_wr[497]     <= 0;                           
					a0_wr[498]     <= 0;                           
					a0_wr[499]     <= 0;                           
					a0_wr[500]     <= 0;                           
					a0_wr[501]     <= 0;                           
					a0_wr[502]     <= 0;                           
					a0_wr[503]     <= 0;                           
					a0_wr[504]     <= 0;                           
					a0_wr[505]     <= 0;                           
					a0_wr[506]     <= 0;                           
					a0_wr[507]     <= 0;                           
					a0_wr[508]     <= 0;                           
					a0_wr[509]     <= 0;                           
					a0_wr[510]     <= 0;                           
					a0_wr[511]     <= 0;                           
					a0_wr[512]     <= 0;                           
					a0_wr[513]     <= 0;                           
					a0_wr[514]     <= 0;                           
					a0_wr[515]     <= 0;                           
					a0_wr[516]     <= 0;                           
					a0_wr[517]     <= 0;                           
					a0_wr[518]     <= 0;                           
					a0_wr[519]     <= 0;                           
					a0_wr[520]     <= 0;                           
					a0_wr[521]     <= 0;                           
					a0_wr[522]     <= 0;                           
					a0_wr[523]     <= 0;                           
					a0_wr[524]     <= 0;                           
					a0_wr[525]     <= 0;                           
					a0_wr[526]     <= 0;                           
					a0_wr[527]     <= 0;                           
					a0_wr[528]     <= 0;                           
					a0_wr[529]     <= 0;                           
					a0_wr[530]     <= 0;                           
					a0_wr[531]     <= 0;                           
					a0_wr[532]     <= 0;                           
					a0_wr[533]     <= 0;                           
					a0_wr[534]     <= 0;                           
					a0_wr[535]     <= 0;                           
					a0_wr[536]     <= 0;                           
					a0_wr[537]     <= 0;                           
					a0_wr[538]     <= 0;                           
					a0_wr[539]     <= 0;                           
					a0_wr[540]     <= 0;                           
					a0_wr[541]     <= 0;                           
					a0_wr[542]     <= 0;                           
					a0_wr[543]     <= 0;                           
					a0_wr[544]     <= 0;                           
					a0_wr[545]     <= 0;                           
					a0_wr[546]     <= 0;                           
					a0_wr[547]     <= 0;                           
					a0_wr[548]     <= 0;                           
					a0_wr[549]     <= 0;                           
					a0_wr[550]     <= 0;                           
					a0_wr[551]     <= 0;                           
					a0_wr[552]     <= 0;                           
					a0_wr[553]     <= 0;                           
					a0_wr[554]     <= 0;                           
					a0_wr[555]     <= 0;                           
					a0_wr[556]     <= 0;                           
					a0_wr[557]     <= 0;                           
					a0_wr[558]     <= 0;                           
					a0_wr[559]     <= 0;                           
					a0_wr[560]     <= 0;                           
					a0_wr[561]     <= 0;                           
					a0_wr[562]     <= 0;                           
					a0_wr[563]     <= 0;                           
					a0_wr[564]     <= 0;                           
					a0_wr[565]     <= 0;                           
					a0_wr[566]     <= 0;                           
					a0_wr[567]     <= 0;                           
					a0_wr[568]     <= 0;                           
					a0_wr[569]     <= 0;                           
					a0_wr[570]     <= 0;                           
					a0_wr[571]     <= 0;                           
					a0_wr[572]     <= 0;                           
					a0_wr[573]     <= 0;                           
					a0_wr[574]     <= 0;                           
					a0_wr[575]     <= 0;                           
					a0_wr[576]     <= 0;                           
					a0_wr[577]     <= 0;                           
					a0_wr[578]     <= 0;                           
					a0_wr[579]     <= 0;                           
					a0_wr[580]     <= 0;                           
					a0_wr[581]     <= 0;                           
					a0_wr[582]     <= 0;                           
					a0_wr[583]     <= 0;                           
					a0_wr[584]     <= 0;                           
					a0_wr[585]     <= 0;                           
					a0_wr[586]     <= 0;                           
					a0_wr[587]     <= 0;                           
					a0_wr[588]     <= 0;                           
					a0_wr[589]     <= 0;                           
					a0_wr[590]     <= 0;                           
					a0_wr[591]     <= 0;                           
					a0_wr[592]     <= 0;                           
					a0_wr[593]     <= 0;                           
					a0_wr[594]     <= 0;                           
					a0_wr[595]     <= 0;                           
					a0_wr[596]     <= 0;                           
					a0_wr[597]     <= 0;                           
					a0_wr[598]     <= 0;                           
					a0_wr[599]     <= 0;                           
					a0_wr[600]     <= 0;                           
					a0_wr[601]     <= 0;                           
					a0_wr[602]     <= 0;                           
					a0_wr[603]     <= 0;                           
					a0_wr[604]     <= 0;                           
					a0_wr[605]     <= 0;                           
					a0_wr[606]     <= 0;                           
					a0_wr[607]     <= 0;                           
					a0_wr[608]     <= 0;                           
					a0_wr[609]     <= 0;                           
					a0_wr[610]     <= 0;                           
					a0_wr[611]     <= 0;                           
					a0_wr[612]     <= 0;                           
					a0_wr[613]     <= 0;                           
					a0_wr[614]     <= 0;                           
					a0_wr[615]     <= 0;                           
					a0_wr[616]     <= 0;                           
					a0_wr[617]     <= 0;                           
					a0_wr[618]     <= 0;                           
					a0_wr[619]     <= 0;                           
					a0_wr[620]     <= 0;                           
					a0_wr[621]     <= 0;                           
					a0_wr[622]     <= 0;                           
					a0_wr[623]     <= 0;                           
					a0_wr[624]     <= 0;                           
					a0_wr[625]     <= 0;                           
					a0_wr[626]     <= 0;                           
					a0_wr[627]     <= 0;                           
					a0_wr[628]     <= 0;                           
					a0_wr[629]     <= 0;                           
					a0_wr[630]     <= 0;                           
					a0_wr[631]     <= 0;                           
					a0_wr[632]     <= 0;                           
					a0_wr[633]     <= 0;                           
					a0_wr[634]     <= 0;                           
					a0_wr[635]     <= 0;                           
					a0_wr[636]     <= 0;                           
					a0_wr[637]     <= 0;                           
					a0_wr[638]     <= 0;                           
					a0_wr[639]     <= 0;                           
					a0_wr[640]     <= 0;                           
					a0_wr[641]     <= 0;                           
					a0_wr[642]     <= 0;                           
					a0_wr[643]     <= 0;                           
					a0_wr[644]     <= 0;                           
					a0_wr[645]     <= 0;                           
					a0_wr[646]     <= 0;                           
					a0_wr[647]     <= 0;                           
					a0_wr[648]     <= 0;                           
					a0_wr[649]     <= 0;                           
					a0_wr[650]     <= 0;                           
					a0_wr[651]     <= 0;                           
					a0_wr[652]     <= 0;                           
					a0_wr[653]     <= 0;                           
					a0_wr[654]     <= 0;                           
					a0_wr[655]     <= 0;                           
					a0_wr[656]     <= 0;                           
					a0_wr[657]     <= 0;                           
					a0_wr[658]     <= 0;                           
					a0_wr[659]     <= 0;                           
					a0_wr[660]     <= 0;                           
					a0_wr[661]     <= 0;                           
					a0_wr[662]     <= 0;                           
					a0_wr[663]     <= 0;                           
					a0_wr[664]     <= 0;                           
					a0_wr[665]     <= 0;                           
					a0_wr[666]     <= 0;                           
					a0_wr[667]     <= 0;                           
					a0_wr[668]     <= 0;                           
					a0_wr[669]     <= 0;                           
					a0_wr[670]     <= 0;                           
					a0_wr[671]     <= 0;                           
					a0_wr[672]     <= 0;                           
					a0_wr[673]     <= 0;                           
					a0_wr[674]     <= 0;                           
					a0_wr[675]     <= 0;                           
					a0_wr[676]     <= 0;                           
					a0_wr[677]     <= 0;                           
					a0_wr[678]     <= 0;                           
					a0_wr[679]     <= 0;                           
					a0_wr[680]     <= 0;                           
					a0_wr[681]     <= 0;                           
					a0_wr[682]     <= 0;                           
					a0_wr[683]     <= 0;                           
					a0_wr[684]     <= 0;                           
					a0_wr[685]     <= 0;                           
					a0_wr[686]     <= 0;                           
					a0_wr[687]     <= 0;                           
					a0_wr[688]     <= 0;                           
					a0_wr[689]     <= 0;                           
					a0_wr[690]     <= 0;                           
					a0_wr[691]     <= 0;                           
					a0_wr[692]     <= 0;                           
					a0_wr[693]     <= 0;                           
					a0_wr[694]     <= 0;                           
					a0_wr[695]     <= 0;                           
					a0_wr[696]     <= 0;                           
					a0_wr[697]     <= 0;                           
					a0_wr[698]     <= 0;                           
					a0_wr[699]     <= 0;                           
					a0_wr[700]     <= 0;                           
					a0_wr[701]     <= 0;                           
					a0_wr[702]     <= 0;                           
					a0_wr[703]     <= 0;                           
					a0_wr[704]     <= 0;                           
					a0_wr[705]     <= 0;                           
					a0_wr[706]     <= 0;                           
					a0_wr[707]     <= 0;                           
					a0_wr[708]     <= 0;                           
					a0_wr[709]     <= 0;                           
					a0_wr[710]     <= 0;                           
					a0_wr[711]     <= 0;                           
					a0_wr[712]     <= 0;                           
					a0_wr[713]     <= 0;                           
					a0_wr[714]     <= 0;                           
					a0_wr[715]     <= 0;                           
					a0_wr[716]     <= 0;                           
					a0_wr[717]     <= 0;                           
					a0_wr[718]     <= 0;                           
					a0_wr[719]     <= 0;                           
					a0_wr[720]     <= 0;                           
					a0_wr[721]     <= 0;                           
					a0_wr[722]     <= 0;                           
					a0_wr[723]     <= 0;                           
					a0_wr[724]     <= 0;                           
					a0_wr[725]     <= 0;                           
					a0_wr[726]     <= 0;                           
					a0_wr[727]     <= 0;                           
					a0_wr[728]     <= 0;                           
					a0_wr[729]     <= 0;                           
					a0_wr[730]     <= 0;                           
					a0_wr[731]     <= 0;                           
					a0_wr[732]     <= 0;                           
					a0_wr[733]     <= 0;                           
					a0_wr[734]     <= 0;                           
					a0_wr[735]     <= 0;                           
					a0_wr[736]     <= 0;                           
					a0_wr[737]     <= 0;                           
					a0_wr[738]     <= 0;                           
					a0_wr[739]     <= 0;                           
					a0_wr[740]     <= 0;                           
					a0_wr[741]     <= 0;                           
					a0_wr[742]     <= 0;                           
					a0_wr[743]     <= 0;                           
					a0_wr[744]     <= 0;                           
					a0_wr[745]     <= 0;                           
					a0_wr[746]     <= 0;                           
					a0_wr[747]     <= 0;                           
					a0_wr[748]     <= 0;                           
					a0_wr[749]     <= 0;                           
					a0_wr[750]     <= 0;                           
					a0_wr[751]     <= 0;                           
					a0_wr[752]     <= 0;                           
					a0_wr[753]     <= 0;                           
					a0_wr[754]     <= 0;                           
					a0_wr[755]     <= 0;                           
					a0_wr[756]     <= 0;                           
					a0_wr[757]     <= 0;                           
					a0_wr[758]     <= 0;                           
					a0_wr[759]     <= 0;                           
					a0_wr[760]     <= 0;                           
					a0_wr[761]     <= 0;                           
					a0_wr[762]     <= 0;                           
					a0_wr[763]     <= 0;                           
					a0_wr[764]     <= 0;                           
					a0_wr[765]     <= 0;                           
					a0_wr[766]     <= 0;                           
					a0_wr[767]     <= 0;                           
					a0_wr[768]     <= 0;                           
					a0_wr[769]     <= 0;                           
					a0_wr[770]     <= 0;                           
					a0_wr[771]     <= 0;                           
					a0_wr[772]     <= 0;                           
					a0_wr[773]     <= 0;                           
					a0_wr[774]     <= 0;                           
					a0_wr[775]     <= 0;                           
					a0_wr[776]     <= 0;                           
					a0_wr[777]     <= 0;                           
					a0_wr[778]     <= 0;                           
					a0_wr[779]     <= 0;                           
					a0_wr[780]     <= 0;                           
					a0_wr[781]     <= 0;                           
					a0_wr[782]     <= 0;                           
					a0_wr[783]     <= 0;                           
					a0_wr[784]     <= 0;                           
					a0_wr[785]     <= 0;                           
					a0_wr[786]     <= 0;                           
					a0_wr[787]     <= 0;                           
					a0_wr[788]     <= 0;                           
					a0_wr[789]     <= 0;                           
					a0_wr[790]     <= 0;                           
					a0_wr[791]     <= 0;                           
					a0_wr[792]     <= 0;                           
					a0_wr[793]     <= 0;                           
					a0_wr[794]     <= 0;                           
					a0_wr[795]     <= 0;                           
					a0_wr[796]     <= 0;                           
					a0_wr[797]     <= 0;                           
					a0_wr[798]     <= 0;                           
					a0_wr[799]     <= 0;                           
					a0_wr[800]     <= 0;                           
					a0_wr[801]     <= 0;                           
					a0_wr[802]     <= 0;                           
					a0_wr[803]     <= 0;                           
					a0_wr[804]     <= 0;                           
					a0_wr[805]     <= 0;                           
					a0_wr[806]     <= 0;                           
					a0_wr[807]     <= 0;                           
					a0_wr[808]     <= 0;                           
					a0_wr[809]     <= 0;                           
					a0_wr[810]     <= 0;                           
					a0_wr[811]     <= 0;                           
					a0_wr[812]     <= 0;                           
					a0_wr[813]     <= 0;                           
					a0_wr[814]     <= 0;                           
					a0_wr[815]     <= 0;                           
					a0_wr[816]     <= 0;                           
					a0_wr[817]     <= 0;                           
					a0_wr[818]     <= 0;                           
					a0_wr[819]     <= 0;                           
					a0_wr[820]     <= 0;                           
					a0_wr[821]     <= 0;                           
					a0_wr[822]     <= 0;                           
					a0_wr[823]     <= 0;                           
					a0_wr[824]     <= 0;                           
					a0_wr[825]     <= 0;                           
					a0_wr[826]     <= 0;                           
					a0_wr[827]     <= 0;                           
					a0_wr[828]     <= 0;                           
					a0_wr[829]     <= 0;                           
					a0_wr[830]     <= 0;                           
					a0_wr[831]     <= 0;                           
					a0_wr[832]     <= 0;                           
					a0_wr[833]     <= 0;                           
					a0_wr[834]     <= 0;                           
					a0_wr[835]     <= 0;                           
					a0_wr[836]     <= 0;                           
					a0_wr[837]     <= 0;                           
					a0_wr[838]     <= 0;                           
					a0_wr[839]     <= 0;                           
					a0_wr[840]     <= 0;                           
					a0_wr[841]     <= 0;                           
					a0_wr[842]     <= 0;                           
					a0_wr[843]     <= 0;                           
					a0_wr[844]     <= 0;                           
					a0_wr[845]     <= 0;                           
					a0_wr[846]     <= 0;                           
					a0_wr[847]     <= 0;                           
					a0_wr[848]     <= 0;                           
					a0_wr[849]     <= 0;                           
					a0_wr[850]     <= 0;                           
					a0_wr[851]     <= 0;                           
					a0_wr[852]     <= 0;                           
					a0_wr[853]     <= 0;                           
					a0_wr[854]     <= 0;                           
					a0_wr[855]     <= 0;                           
					a0_wr[856]     <= 0;                           
					a0_wr[857]     <= 0;                           
					a0_wr[858]     <= 0;                           
					a0_wr[859]     <= 0;                           
					a0_wr[860]     <= 0;                           
					a0_wr[861]     <= 0;                           
					a0_wr[862]     <= 0;                           
					a0_wr[863]     <= 0;                           
					a0_wr[864]     <= 0;                           
					a0_wr[865]     <= 0;                           
					a0_wr[866]     <= 0;                           
					a0_wr[867]     <= 0;                           
					a0_wr[868]     <= 0;                           
					a0_wr[869]     <= 0;                           
					a0_wr[870]     <= 0;                           
					a0_wr[871]     <= 0;                           
					a0_wr[872]     <= 0;                           
					a0_wr[873]     <= 0;                           
					a0_wr[874]     <= 0;                           
					a0_wr[875]     <= 0;                           
					a0_wr[876]     <= 0;                           
					a0_wr[877]     <= 0;                           
					a0_wr[878]     <= 0;                           
					a0_wr[879]     <= 0;                           
					a0_wr[880]     <= 0;                           
					a0_wr[881]     <= 0;                           
					a0_wr[882]     <= 0;                           
					a0_wr[883]     <= 0;                           
					a0_wr[884]     <= 0;                           
					a0_wr[885]     <= 0;                           
					a0_wr[886]     <= 0;                           
					a0_wr[887]     <= 0;                           
					a0_wr[888]     <= 0;                           
					a0_wr[889]     <= 0;                           
					a0_wr[890]     <= 0;                           
					a0_wr[891]     <= 0;                           
					a0_wr[892]     <= 0;                           
					a0_wr[893]     <= 0;                           
					a0_wr[894]     <= 0;                           
					a0_wr[895]     <= 0;                           
					a0_wr[896]     <= 0;                           
					a0_wr[897]     <= 0;                           
					a0_wr[898]     <= 0;                           
					a0_wr[899]     <= 0;                           
					a0_wr[900]     <= 0;                           
					a0_wr[901]     <= 0;                           
					a0_wr[902]     <= 0;                           
					a0_wr[903]     <= 0;                           
					a0_wr[904]     <= 0;                           
					a0_wr[905]     <= 0;                           
					a0_wr[906]     <= 0;                           
					a0_wr[907]     <= 0;                           
					a0_wr[908]     <= 0;                           
					a0_wr[909]     <= 0;                           
					a0_wr[910]     <= 0;                           
					a0_wr[911]     <= 0;                           
					a0_wr[912]     <= 0;                           
					a0_wr[913]     <= 0;                           
					a0_wr[914]     <= 0;                           
					a0_wr[915]     <= 0;                           
					a0_wr[916]     <= 0;                           
					a0_wr[917]     <= 0;                           
					a0_wr[918]     <= 0;                           
					a0_wr[919]     <= 0;                           
					a0_wr[920]     <= 0;                           
					a0_wr[921]     <= 0;                           
					a0_wr[922]     <= 0;                           
					a0_wr[923]     <= 0;                           
					a0_wr[924]     <= 0;                           
					a0_wr[925]     <= 0;                           
					a0_wr[926]     <= 0;                           
					a0_wr[927]     <= 0;                           
					a0_wr[928]     <= 0;                           
					a0_wr[929]     <= 0;                           
					a0_wr[930]     <= 0;                           
					a0_wr[931]     <= 0;                           
					a0_wr[932]     <= 0;                           
					a0_wr[933]     <= 0;                           
					a0_wr[934]     <= 0;                           
					a0_wr[935]     <= 0;                           
					a0_wr[936]     <= 0;                           
					a0_wr[937]     <= 0;                           
					a0_wr[938]     <= 0;                           
					a0_wr[939]     <= 0;                           
					a0_wr[940]     <= 0;                           
					a0_wr[941]     <= 0;                           
					a0_wr[942]     <= 0;                           
					a0_wr[943]     <= 0;                           
					a0_wr[944]     <= 0;                           
					a0_wr[945]     <= 0;                           
					a0_wr[946]     <= 0;                           
					a0_wr[947]     <= 0;                           
					a0_wr[948]     <= 0;                           
					a0_wr[949]     <= 0;                           
					a0_wr[950]     <= 0;                           
					a0_wr[951]     <= 0;                           
					a0_wr[952]     <= 0;                           
					a0_wr[953]     <= 0;                           
					a0_wr[954]     <= 0;                           
					a0_wr[955]     <= 0;                           
					a0_wr[956]     <= 0;                           
					a0_wr[957]     <= 0;                           
					a0_wr[958]     <= 0;                           
					a0_wr[959]     <= 0;                           
					a0_wr[960]     <= 0;                           
					a0_wr[961]     <= 0;                           
					a0_wr[962]     <= 0;                           
					a0_wr[963]     <= 0;                           
					a0_wr[964]     <= 0;                           
					a0_wr[965]     <= 0;                           
					a0_wr[966]     <= 0;                           
					a0_wr[967]     <= 0;                           
					a0_wr[968]     <= 0;                           
					a0_wr[969]     <= 0;                           
					a0_wr[970]     <= 0;                           
					a0_wr[971]     <= 0;                           
					a0_wr[972]     <= 0;                           
					a0_wr[973]     <= 0;                           
					a0_wr[974]     <= 0;                           
					a0_wr[975]     <= 0;                           
					a0_wr[976]     <= 0;                           
					a0_wr[977]     <= 0;                           
					a0_wr[978]     <= 0;                           
					a0_wr[979]     <= 0;                           
					a0_wr[980]     <= 0;                           
					a0_wr[981]     <= 0;                           
					a0_wr[982]     <= 0;                           
					a0_wr[983]     <= 0;                           
					a0_wr[984]     <= 0;                           
					a0_wr[985]     <= 0;                           
					a0_wr[986]     <= 0;                           
					a0_wr[987]     <= 0;                           
					a0_wr[988]     <= 0;                           
					a0_wr[989]     <= 0;                           
					a0_wr[990]     <= 0;                           
					a0_wr[991]     <= 0;                           
					a0_wr[992]     <= 0;                           
					a0_wr[993]     <= 0;                           
					a0_wr[994]     <= 0;                           
					a0_wr[995]     <= 0;                           
					a0_wr[996]     <= 0;                           
					a0_wr[997]     <= 0;                           
					a0_wr[998]     <= 0;                           
					a0_wr[999]     <= 0;                           
					a0_wr[1000]    <= 0;                           
					a0_wr[1001]    <= 0;                           
					a0_wr[1002]    <= 0;                           
					a0_wr[1003]    <= 0;                           
					a0_wr[1004]    <= 0;                           
					a0_wr[1005]    <= 0;                           
					a0_wr[1006]    <= 0;                           
					a0_wr[1007]    <= 0;                           
					a0_wr[1008]    <= 0;                           
					a0_wr[1009]    <= 0;                           
					a0_wr[1010]    <= 0;                           
					a0_wr[1011]    <= 0;                           
					a0_wr[1012]    <= 0;                           
					a0_wr[1013]    <= 0;                           
					a0_wr[1014]    <= 0;                           
					a0_wr[1015]    <= 0;                           
					a0_wr[1016]    <= 0;                           
					a0_wr[1017]    <= 0;                           
					a0_wr[1018]    <= 0;                           
					a0_wr[1019]    <= 0;                           
					a0_wr[1020]    <= 0;                           
					a0_wr[1021]    <= 0;                           
					a0_wr[1022]    <= 0;                           
					a0_wr[1023]    <= 0;                           
					a0_wr[1024]    <= 0;                           
					a0_wr[1025]    <= 0;                           
					a0_wr[1026]    <= 0;                           
					a0_wr[1027]    <= 0;                           
					a0_wr[1028]    <= 0;                           
					a0_wr[1029]    <= 0;                           
					a0_wr[1030]    <= 0;                           
					a0_wr[1031]    <= 0;                           
					a0_wr[1032]    <= 0;                           
					a0_wr[1033]    <= 0;                           
					a0_wr[1034]    <= 0;                           
					a0_wr[1035]    <= 0;                           
					a0_wr[1036]    <= 0;                           
					a0_wr[1037]    <= 0;                           
					a0_wr[1038]    <= 0;                           
					a0_wr[1039]    <= 0;                           
					a0_wr[1040]    <= 0;                           
					a0_wr[1041]    <= 0;                           
					a0_wr[1042]    <= 0;                           
					a0_wr[1043]    <= 0;                           
					a0_wr[1044]    <= 0;                           
					a0_wr[1045]    <= 0;                           
					a0_wr[1046]    <= 0;                           
					a0_wr[1047]    <= 0;                           
					a0_wr[1048]    <= 0;                           
					a0_wr[1049]    <= 0;                           
					a0_wr[1050]    <= 0;                           
					a0_wr[1051]    <= 0;                           
					a0_wr[1052]    <= 0;                           
					a0_wr[1053]    <= 0;                           
					a0_wr[1054]    <= 0;                           
					a0_wr[1055]    <= 0;                           
					a0_wr[1056]    <= 0;                           
					a0_wr[1057]    <= 0;                           
					a0_wr[1058]    <= 0;                           
					a0_wr[1059]    <= 0;                           
					a0_wr[1060]    <= 0;                           
					a0_wr[1061]    <= 0;                           
					a0_wr[1062]    <= 0;                           
					a0_wr[1063]    <= 0;                           
					a0_wr[1064]    <= 0;                           
					a0_wr[1065]    <= 0;                           
					a0_wr[1066]    <= 0;                           
					a0_wr[1067]    <= 0;                           
					a0_wr[1068]    <= 0;                           
					a0_wr[1069]    <= 0;                           
					a0_wr[1070]    <= 0;                           
					a0_wr[1071]    <= 0;                           
					a0_wr[1072]    <= 0;                           
					a0_wr[1073]    <= 0;                           
					a0_wr[1074]    <= 0;                           
					a0_wr[1075]    <= 0;                           
					a0_wr[1076]    <= 0;                           
					a0_wr[1077]    <= 0;                           
					a0_wr[1078]    <= 0;                           
					a0_wr[1079]    <= 0;                           
					a0_wr[1080]    <= 0;                           
					a0_wr[1081]    <= 0;                           
					a0_wr[1082]    <= 0;                           
					a0_wr[1083]    <= 0;                           
					a0_wr[1084]    <= 0;                           
					a0_wr[1085]    <= 0;                           
					a0_wr[1086]    <= 0;                           
					a0_wr[1087]    <= 0;                           
					a0_wr[1088]    <= 0;                           
					a0_wr[1089]    <= 0;                           
					a0_wr[1090]    <= 0;                           
					a0_wr[1091]    <= 0;                           
					a0_wr[1092]    <= 0;                           
					a0_wr[1093]    <= 0;                           
					a0_wr[1094]    <= 0;                           
					a0_wr[1095]    <= 0;                           
					a0_wr[1096]    <= 0;                           
					a0_wr[1097]    <= 0;                           
					a0_wr[1098]    <= 0;                           
					a0_wr[1099]    <= 0;                           
					a0_wr[1100]    <= 0;                           
					a0_wr[1101]    <= 0;                           
					a0_wr[1102]    <= 0;                           
					a0_wr[1103]    <= 0;                           
					a0_wr[1104]    <= 0;                           
					a0_wr[1105]    <= 0;                           
					a0_wr[1106]    <= 0;                           
					a0_wr[1107]    <= 0;                           
					a0_wr[1108]    <= 0;                           
					a0_wr[1109]    <= 0;                           
					a0_wr[1110]    <= 0;                           
					a0_wr[1111]    <= 0;                           
					a0_wr[1112]    <= 0;                           
					a0_wr[1113]    <= 0;                           
					a0_wr[1114]    <= 0;                           
					a0_wr[1115]    <= 0;                           
					a0_wr[1116]    <= 0;                           
					a0_wr[1117]    <= 0;                           
					a0_wr[1118]    <= 0;                           
					a0_wr[1119]    <= 0;                           
					a0_wr[1120]    <= 0;                           
					a0_wr[1121]    <= 0;                           
					a0_wr[1122]    <= 0;                           
					a0_wr[1123]    <= 0;                           
					a0_wr[1124]    <= 0;                           
					a0_wr[1125]    <= 0;                           
					a0_wr[1126]    <= 0;                           
					a0_wr[1127]    <= 0;                           
					a0_wr[1128]    <= 0;                           
					a0_wr[1129]    <= 0;                           
					a0_wr[1130]    <= 0;                           
					a0_wr[1131]    <= 0;                           
					a0_wr[1132]    <= 0;                           
					a0_wr[1133]    <= 0;                           
					a0_wr[1134]    <= 0;                           
					a0_wr[1135]    <= 0;                           
					a0_wr[1136]    <= 0;                           
					a0_wr[1137]    <= 0;                           
					a0_wr[1138]    <= 0;                           
					a0_wr[1139]    <= 0;                           
					a0_wr[1140]    <= 0;                           
					a0_wr[1141]    <= 0;                           
					a0_wr[1142]    <= 0;                           
					a0_wr[1143]    <= 0;                           
					a0_wr[1144]    <= 0;                           
					a0_wr[1145]    <= 0;                           
					a0_wr[1146]    <= 0;                           
					a0_wr[1147]    <= 0;                           
					a0_wr[1148]    <= 0;                           
					a0_wr[1149]    <= 0;                           
					a0_wr[1150]    <= 0;                           
					a0_wr[1151]    <= 0;                           
					a0_wr[1152]    <= 0;                           
					a0_wr[1153]    <= 0;                           
					a0_wr[1154]    <= 0;                           
					a0_wr[1155]    <= 0;                           
					a0_wr[1156]    <= 0;                           
					a0_wr[1157]    <= 0;                           
					a0_wr[1158]    <= 0;                           
					a0_wr[1159]    <= 0;                           
					a0_wr[1160]    <= 0;                           
					a0_wr[1161]    <= 0;                           
					a0_wr[1162]    <= 0;                           
					a0_wr[1163]    <= 0;                           
					a0_wr[1164]    <= 0;                           
					a0_wr[1165]    <= 0;                           
					a0_wr[1166]    <= 0;                           
					a0_wr[1167]    <= 0;                           
					a0_wr[1168]    <= 0;                           
					a0_wr[1169]    <= 0;                           
					a0_wr[1170]    <= 0;                           
					a0_wr[1171]    <= 0;                           
					a0_wr[1172]    <= 0;                           
					a0_wr[1173]    <= 0;                           
					a0_wr[1174]    <= 0;                           
					a0_wr[1175]    <= 0;                           
					a0_wr[1176]    <= 0;                           
					a0_wr[1177]    <= 0;                           
					a0_wr[1178]    <= 0;                           
					a0_wr[1179]    <= 0;                           
					a0_wr[1180]    <= 0;                           
					a0_wr[1181]    <= 0;                           
					a0_wr[1182]    <= 0;                           
					a0_wr[1183]    <= 0;                           
					a0_wr[1184]    <= 0;                           
					a0_wr[1185]    <= 0;                           
					a0_wr[1186]    <= 0;                           
					a0_wr[1187]    <= 0;                           
					a0_wr[1188]    <= 0;                           
					a0_wr[1189]    <= 0;                           
					a0_wr[1190]    <= 0;                           
					a0_wr[1191]    <= 0;                           
					a0_wr[1192]    <= 0;                           
					a0_wr[1193]    <= 0;                           
					a0_wr[1194]    <= 0;                           
					a0_wr[1195]    <= 0;                           
					a0_wr[1196]    <= 0;                           
					a0_wr[1197]    <= 0;                           
					a0_wr[1198]    <= 0;                           
					a0_wr[1199]    <= 0;                           
					a0_wr[1200]    <= 0;                           
					a0_wr[1201]    <= 0;                           
					a0_wr[1202]    <= 0;                           
					a0_wr[1203]    <= 0;                           
					a0_wr[1204]    <= 0;                           
					a0_wr[1205]    <= 0;                           
					a0_wr[1206]    <= 0;                           
					a0_wr[1207]    <= 0;                           
					a0_wr[1208]    <= 0;                           
					a0_wr[1209]    <= 0;                           
					a0_wr[1210]    <= 0;                           
					a0_wr[1211]    <= 0;                           
					a0_wr[1212]    <= 0;                           
					a0_wr[1213]    <= 0;                           
					a0_wr[1214]    <= 0;                           
					a0_wr[1215]    <= 0;                           
					a0_wr[1216]    <= 0;                           
					a0_wr[1217]    <= 0;                           
					a0_wr[1218]    <= 0;                           
					a0_wr[1219]    <= 0;                           
					a0_wr[1220]    <= 0;                           
					a0_wr[1221]    <= 0;                           
					a0_wr[1222]    <= 0;                           
					a0_wr[1223]    <= 0;                           
					a0_wr[1224]    <= 0;                           
					a0_wr[1225]    <= 0;                           
					a0_wr[1226]    <= 0;                           
					a0_wr[1227]    <= 0;                           
					a0_wr[1228]    <= 0;                           
					a0_wr[1229]    <= 0;                           
					a0_wr[1230]    <= 0;                           
					a0_wr[1231]    <= 0;                           
					a0_wr[1232]    <= 0;                           
					a0_wr[1233]    <= 0;                           
					a0_wr[1234]    <= 0;                           
					a0_wr[1235]    <= 0;                           
					a0_wr[1236]    <= 0;                           
					a0_wr[1237]    <= 0;                           
					a0_wr[1238]    <= 0;                           
					a0_wr[1239]    <= 0;                           
					a0_wr[1240]    <= 0;                           
					a0_wr[1241]    <= 0;                           
					a0_wr[1242]    <= 0;                           
					a0_wr[1243]    <= 0;                           
					a0_wr[1244]    <= 0;                           
					a0_wr[1245]    <= 0;                           
					a0_wr[1246]    <= 0;                           
					a0_wr[1247]    <= 0;                           
					a0_wr[1248]    <= 0;                           
					a0_wr[1249]    <= 0;                           
					a0_wr[1250]    <= 0;                           
					a0_wr[1251]    <= 0;                           
					a0_wr[1252]    <= 0;                           
					a0_wr[1253]    <= 0;                           
					a0_wr[1254]    <= 0;                           
					a0_wr[1255]    <= 0;                           
					a0_wr[1256]    <= 0;                           
					a0_wr[1257]    <= 0;                           
					a0_wr[1258]    <= 0;                           
					a0_wr[1259]    <= 0;                           
					a0_wr[1260]    <= 0;                           
					a0_wr[1261]    <= 0;                           
					a0_wr[1262]    <= 0;                           
					a0_wr[1263]    <= 0;                           
					a0_wr[1264]    <= 0;                           
					a0_wr[1265]    <= 0;                           
					a0_wr[1266]    <= 0;                           
					a0_wr[1267]    <= 0;                           
					a0_wr[1268]    <= 0;                           
					a0_wr[1269]    <= 0;                           
					a0_wr[1270]    <= 0;                           
					a0_wr[1271]    <= 0;                           
					a0_wr[1272]    <= 0;                           
					a0_wr[1273]    <= 0;                           
					a0_wr[1274]    <= 0;                           
					a0_wr[1275]    <= 0;                           
					a0_wr[1276]    <= 0;                           
					a0_wr[1277]    <= 0;                           
					a0_wr[1278]    <= 0;                           
					a0_wr[1279]    <= 0;                           
					a0_wr[1280]    <= 0;                           
					a0_wr[1281]    <= 0;                           
					a0_wr[1282]    <= 0;                           
					a0_wr[1283]    <= 0;                           
					a0_wr[1284]    <= 0;                           
					a0_wr[1285]    <= 0;                           
					a0_wr[1286]    <= 0;                           
					a0_wr[1287]    <= 0;                           
					a0_wr[1288]    <= 0;                           
					a0_wr[1289]    <= 0;                           
					a0_wr[1290]    <= 0;                           
					a0_wr[1291]    <= 0;                           
					a0_wr[1292]    <= 0;                           
					a0_wr[1293]    <= 0;                           
					a0_wr[1294]    <= 0;                           
					a0_wr[1295]    <= 0;                           
					a0_wr[1296]    <= 0;                           
					a0_wr[1297]    <= 0;                           
					a0_wr[1298]    <= 0;                           
					a0_wr[1299]    <= 0;                           
					a0_wr[1300]    <= 0;                           
					a0_wr[1301]    <= 0;                           
					a0_wr[1302]    <= 0;                           
					a0_wr[1303]    <= 0;                           
					a0_wr[1304]    <= 0;                           
					a0_wr[1305]    <= 0;                           
					a0_wr[1306]    <= 0;                           
					a0_wr[1307]    <= 0;                           
					a0_wr[1308]    <= 0;                           
					a0_wr[1309]    <= 0;                           
					a0_wr[1310]    <= 0;                           
					a0_wr[1311]    <= 0;                           
					a0_wr[1312]    <= 0;                           
					a0_wr[1313]    <= 0;                           
					a0_wr[1314]    <= 0;                           
					a0_wr[1315]    <= 0;                           
					a0_wr[1316]    <= 0;                           
					a0_wr[1317]    <= 0;                           
					a0_wr[1318]    <= 0;                           
					a0_wr[1319]    <= 0;                           
					a0_wr[1320]    <= 0;                           
					a0_wr[1321]    <= 0;                           
					a0_wr[1322]    <= 0;                           
					a0_wr[1323]    <= 0;                           
					a0_wr[1324]    <= 0;                           
					a0_wr[1325]    <= 0;                           
					a0_wr[1326]    <= 0;                           
					a0_wr[1327]    <= 0;                           
					a0_wr[1328]    <= 0;                           
					a0_wr[1329]    <= 0;                           
					a0_wr[1330]    <= 0;                           
					a0_wr[1331]    <= 0;                           
					a0_wr[1332]    <= 0;                           
					a0_wr[1333]    <= 0;                           
					a0_wr[1334]    <= 0;                           
					a0_wr[1335]    <= 0;                           
					a0_wr[1336]    <= 0;                           
					a0_wr[1337]    <= 0;                           
					a0_wr[1338]    <= 0;                           
					a0_wr[1339]    <= 0;                           
					a0_wr[1340]    <= 0;                           
					a0_wr[1341]    <= 0;                           
					a0_wr[1342]    <= 0;                           
					a0_wr[1343]    <= 0;                           
					a0_wr[1344]    <= 0;                           
					a0_wr[1345]    <= 0;                           
					a0_wr[1346]    <= 0;                           
					a0_wr[1347]    <= 0;                           
					a0_wr[1348]    <= 0;                           
					a0_wr[1349]    <= 0;                           
					a0_wr[1350]    <= 0;                           
					a0_wr[1351]    <= 0;                           
					a0_wr[1352]    <= 0;                           
					a0_wr[1353]    <= 0;                           
					a0_wr[1354]    <= 0;                           
					a0_wr[1355]    <= 0;                           
					a0_wr[1356]    <= 0;                           
					a0_wr[1357]    <= 0;                           
					a0_wr[1358]    <= 0;                           
					a0_wr[1359]    <= 0;                           
					a0_wr[1360]    <= 0;                           
					a0_wr[1361]    <= 0;                           
					a0_wr[1362]    <= 0;                           
					a0_wr[1363]    <= 0;                           
					a0_wr[1364]    <= 0;                           
					a0_wr[1365]    <= 0;                           
					a0_wr[1366]    <= 0;                           
					a0_wr[1367]    <= 0;                           
					a0_wr[1368]    <= 0;                           
					a0_wr[1369]    <= 0;                           
					a0_wr[1370]    <= 0;                           
					a0_wr[1371]    <= 0;                           
					a0_wr[1372]    <= 0;                           
					a0_wr[1373]    <= 0;                           
					a0_wr[1374]    <= 0;                           
					a0_wr[1375]    <= 0;                           
					a0_wr[1376]    <= 0;                           
					a0_wr[1377]    <= 0;                           
					a0_wr[1378]    <= 0;                           
					a0_wr[1379]    <= 0;                           
					a0_wr[1380]    <= 0;                           
					a0_wr[1381]    <= 0;                           
					a0_wr[1382]    <= 0;                           
					a0_wr[1383]    <= 0;                           
					a0_wr[1384]    <= 0;                           
					a0_wr[1385]    <= 0;                           
					a0_wr[1386]    <= 0;                           
					a0_wr[1387]    <= 0;                           
					a0_wr[1388]    <= 0;                           
					a0_wr[1389]    <= 0;                           
					a0_wr[1390]    <= 0;                           
					a0_wr[1391]    <= 0;                           
					a0_wr[1392]    <= 0;                           
					a0_wr[1393]    <= 0;                           
					a0_wr[1394]    <= 0;                           
					a0_wr[1395]    <= 0;                           
					a0_wr[1396]    <= 0;                           
					a0_wr[1397]    <= 0;                           
					a0_wr[1398]    <= 0;                           
					a0_wr[1399]    <= 0;                           
					a0_wr[1400]    <= 0;                           
					a0_wr[1401]    <= 0;                           
					a0_wr[1402]    <= 0;                           
					a0_wr[1403]    <= 0;                           
					a0_wr[1404]    <= 0;                           
					a0_wr[1405]    <= 0;                           
					a0_wr[1406]    <= 0;                           
					a0_wr[1407]    <= 0;                           
					a0_wr[1408]    <= 0;                           
					a0_wr[1409]    <= 0;                           
					a0_wr[1410]    <= 0;                           
					a0_wr[1411]    <= 0;                           
					a0_wr[1412]    <= 0;                           
					a0_wr[1413]    <= 0;                           
					a0_wr[1414]    <= 0;                           
					a0_wr[1415]    <= 0;                           
					a0_wr[1416]    <= 0;                           
					a0_wr[1417]    <= 0;                           
					a0_wr[1418]    <= 0;                           
					a0_wr[1419]    <= 0;                           
					a0_wr[1420]    <= 0;                           
					a0_wr[1421]    <= 0;                           
					a0_wr[1422]    <= 0;                           
					a0_wr[1423]    <= 0;                           
					a0_wr[1424]    <= 0;                           
					a0_wr[1425]    <= 0;                           
					a0_wr[1426]    <= 0;                           
					a0_wr[1427]    <= 0;                           
					a0_wr[1428]    <= 0;                           
					a0_wr[1429]    <= 0;                           
					a0_wr[1430]    <= 0;                           
					a0_wr[1431]    <= 0;                           
					a0_wr[1432]    <= 0;                           
					a0_wr[1433]    <= 0;                           
					a0_wr[1434]    <= 0;                           
					a0_wr[1435]    <= 0;                           
					a0_wr[1436]    <= 0;                           
					a0_wr[1437]    <= 0;                           
					a0_wr[1438]    <= 0;                           
					a0_wr[1439]    <= 0;                           
					a0_wr[1440]    <= 0;                           
					a0_wr[1441]    <= 0;                           
					a0_wr[1442]    <= 0;                           
					a0_wr[1443]    <= 0;                           
					a0_wr[1444]    <= 0;                           
					a0_wr[1445]    <= 0;                           
					a0_wr[1446]    <= 0;                           
					a0_wr[1447]    <= 0;                           
					a0_wr[1448]    <= 0;                           
					a0_wr[1449]    <= 0;                           
					a0_wr[1450]    <= 0;                           
					a0_wr[1451]    <= 0;                           
					a0_wr[1452]    <= 0;                           
					a0_wr[1453]    <= 0;                           
					a0_wr[1454]    <= 0;                           
					a0_wr[1455]    <= 0;                           
					a0_wr[1456]    <= 0;                           
					a0_wr[1457]    <= 0;                           
					a0_wr[1458]    <= 0;                           
					a0_wr[1459]    <= 0;                           
					a0_wr[1460]    <= 0;                           
					a0_wr[1461]    <= 0;                           
					a0_wr[1462]    <= 0;                           
					a0_wr[1463]    <= 0;                           
					a0_wr[1464]    <= 0;                           
					a0_wr[1465]    <= 0;                           
					a0_wr[1466]    <= 0;                           
					a0_wr[1467]    <= 0;                           
					a0_wr[1468]    <= 0;                           
					a0_wr[1469]    <= 0;                           
					a0_wr[1470]    <= 0;                           
					a0_wr[1471]    <= 0;                           
					a0_wr[1472]    <= 0;                           
					a0_wr[1473]    <= 0;                           
					a0_wr[1474]    <= 0;                           
					a0_wr[1475]    <= 0;                           
					a0_wr[1476]    <= 0;                           
					a0_wr[1477]    <= 0;                           
					a0_wr[1478]    <= 0;                           
					a0_wr[1479]    <= 0;                           
					a0_wr[1480]    <= 0;                           
					a0_wr[1481]    <= 0;                           
					a0_wr[1482]    <= 0;                           
					a0_wr[1483]    <= 0;                           
					a0_wr[1484]    <= 0;                           
					a0_wr[1485]    <= 0;                           
					a0_wr[1486]    <= 0;                           
					a0_wr[1487]    <= 0;                           
					a0_wr[1488]    <= 0;                           
					a0_wr[1489]    <= 0;                           
					a0_wr[1490]    <= 0;                           
					a0_wr[1491]    <= 0;                           
					a0_wr[1492]    <= 0;                           
					a0_wr[1493]    <= 0;                           
					a0_wr[1494]    <= 0;                           
					a0_wr[1495]    <= 0;                           
					a0_wr[1496]    <= 0;                           
					a0_wr[1497]    <= 0;                           
					a0_wr[1498]    <= 0;                           
					a0_wr[1499]    <= 0;                           
					a0_wr[1500]    <= 0;                           
					a0_wr[1501]    <= 0;                           
					a0_wr[1502]    <= 0;                           
					a0_wr[1503]    <= 0;                           
					a0_wr[1504]    <= 0;                           
					a0_wr[1505]    <= 0;                           
					a0_wr[1506]    <= 0;                           
					a0_wr[1507]    <= 0;                           
					a0_wr[1508]    <= 0;                           
					a0_wr[1509]    <= 0;                           
					a0_wr[1510]    <= 0;                           
					a0_wr[1511]    <= 0;                           
					a0_wr[1512]    <= 0;                           
					a0_wr[1513]    <= 0;                           
					a0_wr[1514]    <= 0;                           
					a0_wr[1515]    <= 0;                           
					a0_wr[1516]    <= 0;                           
					a0_wr[1517]    <= 0;                           
					a0_wr[1518]    <= 0;                           
					a0_wr[1519]    <= 0;                           
					a0_wr[1520]    <= 0;                           
					a0_wr[1521]    <= 0;                           
					a0_wr[1522]    <= 0;                           
					a0_wr[1523]    <= 0;                           
					a0_wr[1524]    <= 0;                           
					a0_wr[1525]    <= 0;                           
					a0_wr[1526]    <= 0;                           
					a0_wr[1527]    <= 0;                           
					a0_wr[1528]    <= 0;                           
					a0_wr[1529]    <= 0;                           
					a0_wr[1530]    <= 0;                           
					a0_wr[1531]    <= 0;                           
					a0_wr[1532]    <= 0;                           
					a0_wr[1533]    <= 0;                           
					a0_wr[1534]    <= 0;                           
					a0_wr[1535]    <= 0;                           
					a0_wr[1536]    <= 0;                           
					a0_wr[1537]    <= 0;                           
					a0_wr[1538]    <= 0;                           
					a0_wr[1539]    <= 0;                           
					a0_wr[1540]    <= 0;                           
					a0_wr[1541]    <= 0;                           
					a0_wr[1542]    <= 0;                           
					a0_wr[1543]    <= 0;                           
					a0_wr[1544]    <= 0;                           
					a0_wr[1545]    <= 0;                           
					a0_wr[1546]    <= 0;                           
					a0_wr[1547]    <= 0;                           
					a0_wr[1548]    <= 0;                           
					a0_wr[1549]    <= 0;                           
					a0_wr[1550]    <= 0;                           
					a0_wr[1551]    <= 0;                           
					a0_wr[1552]    <= 0;                           
					a0_wr[1553]    <= 0;                           
					a0_wr[1554]    <= 0;                           
					a0_wr[1555]    <= 0;                           
					a0_wr[1556]    <= 0;                           
					a0_wr[1557]    <= 0;                           
					a0_wr[1558]    <= 0;                           
					a0_wr[1559]    <= 0;                           
					a0_wr[1560]    <= 0;                           
					a0_wr[1561]    <= 0;                           
					a0_wr[1562]    <= 0;                           
					a0_wr[1563]    <= 0;                           
					a0_wr[1564]    <= 0;                           
					a0_wr[1565]    <= 0;                           
					a0_wr[1566]    <= 0;                           
					a0_wr[1567]    <= 0;                           
					a0_wr[1568]    <= 0;                           
					a0_wr[1569]    <= 0;                           
					a0_wr[1570]    <= 0;                           
					a0_wr[1571]    <= 0;                           
					a0_wr[1572]    <= 0;                           
					a0_wr[1573]    <= 0;                           
					a0_wr[1574]    <= 0;                           
					a0_wr[1575]    <= 0;                           
					a0_wr[1576]    <= 0;                           
					a0_wr[1577]    <= 0;                           
					a0_wr[1578]    <= 0;                           
					a0_wr[1579]    <= 0;                           
					a0_wr[1580]    <= 0;                           
					a0_wr[1581]    <= 0;                           
					a0_wr[1582]    <= 0;                           
					a0_wr[1583]    <= 0;                           
					a0_wr[1584]    <= 0;                           
					a0_wr[1585]    <= 0;                           
					a0_wr[1586]    <= 0;                           
					a0_wr[1587]    <= 0;                           
					a0_wr[1588]    <= 0;                           
					a0_wr[1589]    <= 0;                           
					a0_wr[1590]    <= 0;                           
					a0_wr[1591]    <= 0;                           
					a0_wr[1592]    <= 0;                           
					a0_wr[1593]    <= 0;                           
					a0_wr[1594]    <= 0;                           
					a0_wr[1595]    <= 0;                           
					a0_wr[1596]    <= 0;                           
					a0_wr[1597]    <= 0;                           
					a0_wr[1598]    <= 0;                           
					a0_wr[1599]    <= 0;                           
					a0_wr[1600]    <= 0;                           
					a0_wr[1601]    <= 0;                           
					a0_wr[1602]    <= 0;                           
					a0_wr[1603]    <= 0;                           
					a0_wr[1604]    <= 0;                           
					a0_wr[1605]    <= 0;                           
					a0_wr[1606]    <= 0;                           
					a0_wr[1607]    <= 0;                           
					a0_wr[1608]    <= 0;                           
					a0_wr[1609]    <= 0;                           
					a0_wr[1610]    <= 0;                           
					a0_wr[1611]    <= 0;                           
					a0_wr[1612]    <= 0;                           
					a0_wr[1613]    <= 0;                           
					a0_wr[1614]    <= 0;                           
					a0_wr[1615]    <= 0;                           
					a0_wr[1616]    <= 0;                           
					a0_wr[1617]    <= 0;                           
					a0_wr[1618]    <= 0;                           
					a0_wr[1619]    <= 0;                           
					a0_wr[1620]    <= 0;                           
					a0_wr[1621]    <= 0;                           
					a0_wr[1622]    <= 0;                           
					a0_wr[1623]    <= 0;                           
					a0_wr[1624]    <= 0;                           
					a0_wr[1625]    <= 0;                           
					a0_wr[1626]    <= 0;                           
					a0_wr[1627]    <= 0;                           
					a0_wr[1628]    <= 0;                           
					a0_wr[1629]    <= 0;                           
					a0_wr[1630]    <= 0;                           
					a0_wr[1631]    <= 0;                           
					a0_wr[1632]    <= 0;                           
					a0_wr[1633]    <= 0;                           
					a0_wr[1634]    <= 0;                           
					a0_wr[1635]    <= 0;                           
					a0_wr[1636]    <= 0;                           
					a0_wr[1637]    <= 0;                           
					a0_wr[1638]    <= 0;                           
					a0_wr[1639]    <= 0;                           
					a0_wr[1640]    <= 0;                           
					a0_wr[1641]    <= 0;                           
					a0_wr[1642]    <= 0;                           
					a0_wr[1643]    <= 0;                           
					a0_wr[1644]    <= 0;                           
					a0_wr[1645]    <= 0;                           
					a0_wr[1646]    <= 0;                           
					a0_wr[1647]    <= 0;                           
					a0_wr[1648]    <= 0;                           
					a0_wr[1649]    <= 0;                           
					a0_wr[1650]    <= 0;                           
					a0_wr[1651]    <= 0;                           
					a0_wr[1652]    <= 0;                           
					a0_wr[1653]    <= 0;                           
					a0_wr[1654]    <= 0;                           
					a0_wr[1655]    <= 0;                           
					a0_wr[1656]    <= 0;                           
					a0_wr[1657]    <= 0;                           
					a0_wr[1658]    <= 0;                           
					a0_wr[1659]    <= 0;                           
					a0_wr[1660]    <= 0;                           
					a0_wr[1661]    <= 0;                           
					a0_wr[1662]    <= 0;                           
					a0_wr[1663]    <= 0;                           
					a0_wr[1664]    <= 0;                           
					a0_wr[1665]    <= 0;                           
					a0_wr[1666]    <= 0;                           
					a0_wr[1667]    <= 0;                           
					a0_wr[1668]    <= 0;                           
					a0_wr[1669]    <= 0;                           
					a0_wr[1670]    <= 0;                           
					a0_wr[1671]    <= 0;                           
					a0_wr[1672]    <= 0;                           
					a0_wr[1673]    <= 0;                           
					a0_wr[1674]    <= 0;                           
					a0_wr[1675]    <= 0;                           
					a0_wr[1676]    <= 0;                           
					a0_wr[1677]    <= 0;                           
					a0_wr[1678]    <= 0;                           
					a0_wr[1679]    <= 0;                           
					a0_wr[1680]    <= 0;                           
					a0_wr[1681]    <= 0;                           
					a0_wr[1682]    <= 0;                           
					a0_wr[1683]    <= 0;                           
					a0_wr[1684]    <= 0;                           
					a0_wr[1685]    <= 0;                           
					a0_wr[1686]    <= 0;                           
					a0_wr[1687]    <= 0;                           
					a0_wr[1688]    <= 0;                           
					a0_wr[1689]    <= 0;                           
					a0_wr[1690]    <= 0;                           
					a0_wr[1691]    <= 0;                           
					a0_wr[1692]    <= 0;                           
					a0_wr[1693]    <= 0;                           
					a0_wr[1694]    <= 0;                           
					a0_wr[1695]    <= 0;                           
					a0_wr[1696]    <= 0;                           
					a0_wr[1697]    <= 0;                           
					a0_wr[1698]    <= 0;                           
					a0_wr[1699]    <= 0;                           
					a0_wr[1700]    <= 0;                           
					a0_wr[1701]    <= 0;                           
					a0_wr[1702]    <= 0;                           
					a0_wr[1703]    <= 0;                           
					a0_wr[1704]    <= 0;                           
					a0_wr[1705]    <= 0;                           
					a0_wr[1706]    <= 0;                           
					a0_wr[1707]    <= 0;                           
					a0_wr[1708]    <= 0;                           
					a0_wr[1709]    <= 0;                           
					a0_wr[1710]    <= 0;                           
					a0_wr[1711]    <= 0;                           
					a0_wr[1712]    <= 0;                           
					a0_wr[1713]    <= 0;                           
					a0_wr[1714]    <= 0;                           
					a0_wr[1715]    <= 0;                           
					a0_wr[1716]    <= 0;                           
					a0_wr[1717]    <= 0;                           
					a0_wr[1718]    <= 0;                           
					a0_wr[1719]    <= 0;                           
					a0_wr[1720]    <= 0;                           
					a0_wr[1721]    <= 0;                           
					a0_wr[1722]    <= 0;                           
					a0_wr[1723]    <= 0;                           
					a0_wr[1724]    <= 0;                           
					a0_wr[1725]    <= 0;                           
					a0_wr[1726]    <= 0;                           
					a0_wr[1727]    <= 0;                           
					a0_wr[1728]    <= 0;                           
					a0_wr[1729]    <= 0;                           
					a0_wr[1730]    <= 0;                           
					a0_wr[1731]    <= 0;                           
					a0_wr[1732]    <= 0;                           
					a0_wr[1733]    <= 0;                           
					a0_wr[1734]    <= 0;                           
					a0_wr[1735]    <= 0;                           
					a0_wr[1736]    <= 0;                           
					a0_wr[1737]    <= 0;                           
					a0_wr[1738]    <= 0;                           
					a0_wr[1739]    <= 0;                           
					a0_wr[1740]    <= 0;                           
					a0_wr[1741]    <= 0;                           
					a0_wr[1742]    <= 0;                           
					a0_wr[1743]    <= 0;                           
					a0_wr[1744]    <= 0;                           
					a0_wr[1745]    <= 0;                           
					a0_wr[1746]    <= 0;                           
					a0_wr[1747]    <= 0;                           
					a0_wr[1748]    <= 0;                           
					a0_wr[1749]    <= 0;                           
					a0_wr[1750]    <= 0;                           
					a0_wr[1751]    <= 0;                           
					a0_wr[1752]    <= 0;                           
					a0_wr[1753]    <= 0;                           
					a0_wr[1754]    <= 0;                           
					a0_wr[1755]    <= 0;                           
					a0_wr[1756]    <= 0;                           
					a0_wr[1757]    <= 0;                           
					a0_wr[1758]    <= 0;                           
					a0_wr[1759]    <= 0;                           
					a0_wr[1760]    <= 0;                           
					a0_wr[1761]    <= 0;                           
					a0_wr[1762]    <= 0;                           
					a0_wr[1763]    <= 0;                           
					a0_wr[1764]    <= 0;                           
					a0_wr[1765]    <= 0;                           
					a0_wr[1766]    <= 0;                           
					a0_wr[1767]    <= 0;                           
					a0_wr[1768]    <= 0;                           
					a0_wr[1769]    <= 0;                           
					a0_wr[1770]    <= 0;                           
					a0_wr[1771]    <= 0;                           
					a0_wr[1772]    <= 0;                           
					a0_wr[1773]    <= 0;                           
					a0_wr[1774]    <= 0;                           
					a0_wr[1775]    <= 0;                           
					a0_wr[1776]    <= 0;                           
					a0_wr[1777]    <= 0;                           
					a0_wr[1778]    <= 0;                           
					a0_wr[1779]    <= 0;                           
					a0_wr[1780]    <= 0;                           
					a0_wr[1781]    <= 0;                           
					a0_wr[1782]    <= 0;                           
					a0_wr[1783]    <= 0;                           
					a0_wr[1784]    <= 0;                           
					a0_wr[1785]    <= 0;                           
					a0_wr[1786]    <= 0;                           
					a0_wr[1787]    <= 0;                           
					a0_wr[1788]    <= 0;                           
					a0_wr[1789]    <= 0;                           
					a0_wr[1790]    <= 0;                           
					a0_wr[1791]    <= 0;                           
					a0_wr[1792]    <= 0;                           
					a0_wr[1793]    <= 0;                           
					a0_wr[1794]    <= 0;                           
					a0_wr[1795]    <= 0;                           
					a0_wr[1796]    <= 0;                           
					a0_wr[1797]    <= 0;                           
					a0_wr[1798]    <= 0;                           
					a0_wr[1799]    <= 0;                           
					a0_wr[1800]    <= 0;                           
					a0_wr[1801]    <= 0;                           
					a0_wr[1802]    <= 0;                           
					a0_wr[1803]    <= 0;                           
					a0_wr[1804]    <= 0;                           
					a0_wr[1805]    <= 0;                           
					a0_wr[1806]    <= 0;                           
					a0_wr[1807]    <= 0;                           
					a0_wr[1808]    <= 0;                           
					a0_wr[1809]    <= 0;                           
					a0_wr[1810]    <= 0;                           
					a0_wr[1811]    <= 0;                           
					a0_wr[1812]    <= 0;                           
					a0_wr[1813]    <= 0;                           
					a0_wr[1814]    <= 0;                           
					a0_wr[1815]    <= 0;                           
					a0_wr[1816]    <= 0;                           
					a0_wr[1817]    <= 0;                           
					a0_wr[1818]    <= 0;                           
					a0_wr[1819]    <= 0;                           
					a0_wr[1820]    <= 0;                           
					a0_wr[1821]    <= 0;                           
					a0_wr[1822]    <= 0;                           
					a0_wr[1823]    <= 0;                           
					a0_wr[1824]    <= 0;                           
					a0_wr[1825]    <= 0;                           
					a0_wr[1826]    <= 0;                           
					a0_wr[1827]    <= 0;                           
					a0_wr[1828]    <= 0;                           
					a0_wr[1829]    <= 0;                           
					a0_wr[1830]    <= 0;                           
					a0_wr[1831]    <= 0;                           
					a0_wr[1832]    <= 0;                           
					a0_wr[1833]    <= 0;                           
					a0_wr[1834]    <= 0;                           
					a0_wr[1835]    <= 0;                           
					a0_wr[1836]    <= 0;                           
					a0_wr[1837]    <= 0;                           
					a0_wr[1838]    <= 0;                           
					a0_wr[1839]    <= 0;                           
					a0_wr[1840]    <= 0;                           
					a0_wr[1841]    <= 0;                           
					a0_wr[1842]    <= 0;                           
					a0_wr[1843]    <= 0;                           
					a0_wr[1844]    <= 0;                           
					a0_wr[1845]    <= 0;                           
					a0_wr[1846]    <= 0;                           
					a0_wr[1847]    <= 0;                           
					a0_wr[1848]    <= 0;                           
					a0_wr[1849]    <= 0;                           
					a0_wr[1850]    <= 0;                           
					a0_wr[1851]    <= 0;                           
					a0_wr[1852]    <= 0;                           
					a0_wr[1853]    <= 0;                           
					a0_wr[1854]    <= 0;                           
					a0_wr[1855]    <= 0;                           
					a0_wr[1856]    <= 0;                           
					a0_wr[1857]    <= 0;                           
					a0_wr[1858]    <= 0;                           
					a0_wr[1859]    <= 0;                           
					a0_wr[1860]    <= 0;                           
					a0_wr[1861]    <= 0;                           
					a0_wr[1862]    <= 0;                           
					a0_wr[1863]    <= 0;                           
					a0_wr[1864]    <= 0;                           
					a0_wr[1865]    <= 0;                           
					a0_wr[1866]    <= 0;                           
					a0_wr[1867]    <= 0;                           
					a0_wr[1868]    <= 0;                           
					a0_wr[1869]    <= 0;                           
					a0_wr[1870]    <= 0;                           
					a0_wr[1871]    <= 0;                           
					a0_wr[1872]    <= 0;                           
					a0_wr[1873]    <= 0;                           
					a0_wr[1874]    <= 0;                           
					a0_wr[1875]    <= 0;                           
					a0_wr[1876]    <= 0;                           
					a0_wr[1877]    <= 0;                           
					a0_wr[1878]    <= 0;                           
					a0_wr[1879]    <= 0;                           
					a0_wr[1880]    <= 0;                           
					a0_wr[1881]    <= 0;                           
					a0_wr[1882]    <= 0;                           
					a0_wr[1883]    <= 0;                           
					a0_wr[1884]    <= 0;                           
					a0_wr[1885]    <= 0;                           
					a0_wr[1886]    <= 0;                           
					a0_wr[1887]    <= 0;                           
					a0_wr[1888]    <= 0;                           
					a0_wr[1889]    <= 0;                           
					a0_wr[1890]    <= 0;                           
					a0_wr[1891]    <= 0;                           
					a0_wr[1892]    <= 0;                           
					a0_wr[1893]    <= 0;                           
					a0_wr[1894]    <= 0;                           
					a0_wr[1895]    <= 0;                           
					a0_wr[1896]    <= 0;                           
					a0_wr[1897]    <= 0;                           
					a0_wr[1898]    <= 0;                           
					a0_wr[1899]    <= 0;                           
					a0_wr[1900]    <= 0;                           
					a0_wr[1901]    <= 0;                           
					a0_wr[1902]    <= 0;                           
					a0_wr[1903]    <= 0;                           
					a0_wr[1904]    <= 0;                           
					a0_wr[1905]    <= 0;                           
					a0_wr[1906]    <= 0;                           
					a0_wr[1907]    <= 0;                           
					a0_wr[1908]    <= 0;                           
					a0_wr[1909]    <= 0;                           
					a0_wr[1910]    <= 0;                           
					a0_wr[1911]    <= 0;                           
					a0_wr[1912]    <= 0;                           
					a0_wr[1913]    <= 0;                           
					a0_wr[1914]    <= 0;                           
					a0_wr[1915]    <= 0;                           
					a0_wr[1916]    <= 0;                           
					a0_wr[1917]    <= 0;                           
					a0_wr[1918]    <= 0;                           
					a0_wr[1919]    <= 0;                           
					a0_wr[1920]    <= 0;                           
					a0_wr[1921]    <= 0;                           
					a0_wr[1922]    <= 0;                           
					a0_wr[1923]    <= 0;                           
					a0_wr[1924]    <= 0;                           
					a0_wr[1925]    <= 0;                           
					a0_wr[1926]    <= 0;                           
					a0_wr[1927]    <= 0;                           
					a0_wr[1928]    <= 0;                           
					a0_wr[1929]    <= 0;                           
					a0_wr[1930]    <= 0;                           
					a0_wr[1931]    <= 0;                           
					a0_wr[1932]    <= 0;                           
					a0_wr[1933]    <= 0;                           
					a0_wr[1934]    <= 0;                           
					a0_wr[1935]    <= 0;                           
					a0_wr[1936]    <= 0;                           
					a0_wr[1937]    <= 0;                           
					a0_wr[1938]    <= 0;                           
					a0_wr[1939]    <= 0;                           
					a0_wr[1940]    <= 0;                           
					a0_wr[1941]    <= 0;                           
					a0_wr[1942]    <= 0;                           
					a0_wr[1943]    <= 0;                           
					a0_wr[1944]    <= 0;                           
					a0_wr[1945]    <= 0;                           
					a0_wr[1946]    <= 0;                           
					a0_wr[1947]    <= 0;                           
					a0_wr[1948]    <= 0;                           
					a0_wr[1949]    <= 0;                           
					a0_wr[1950]    <= 0;                           
					a0_wr[1951]    <= 0;                           
					a0_wr[1952]    <= 0;                           
					a0_wr[1953]    <= 0;                           
					a0_wr[1954]    <= 0;                           
					a0_wr[1955]    <= 0;                           
					a0_wr[1956]    <= 0;                           
					a0_wr[1957]    <= 0;                           
					a0_wr[1958]    <= 0;                           
					a0_wr[1959]    <= 0;                           
					a0_wr[1960]    <= 0;                           
					a0_wr[1961]    <= 0;                           
					a0_wr[1962]    <= 0;                           
					a0_wr[1963]    <= 0;                           
					a0_wr[1964]    <= 0;                           
					a0_wr[1965]    <= 0;                           
					a0_wr[1966]    <= 0;                           
					a0_wr[1967]    <= 0;                           
					a0_wr[1968]    <= 0;                           
					a0_wr[1969]    <= 0;                           
					a0_wr[1970]    <= 0;                           
					a0_wr[1971]    <= 0;                           
					a0_wr[1972]    <= 0;                           
					a0_wr[1973]    <= 0;                           
					a0_wr[1974]    <= 0;                           
					a0_wr[1975]    <= 0;                           
					a0_wr[1976]    <= 0;                           
					a0_wr[1977]    <= 0;                           
					a0_wr[1978]    <= 0;                           
					a0_wr[1979]    <= 0;                           
					a0_wr[1980]    <= 0;                           
					a0_wr[1981]    <= 0;                           
					a0_wr[1982]    <= 0;                           
					a0_wr[1983]    <= 0;                           
					a0_wr[1984]    <= 0;                           
					a0_wr[1985]    <= 0;                           
					a0_wr[1986]    <= 0;                           
					a0_wr[1987]    <= 0;                           
					a0_wr[1988]    <= 0;                           
					a0_wr[1989]    <= 0;                           
					a0_wr[1990]    <= 0;                           
					a0_wr[1991]    <= 0;                           
					a0_wr[1992]    <= 0;                           
					a0_wr[1993]    <= 0;                           
					a0_wr[1994]    <= 0;                           
					a0_wr[1995]    <= 0;                           
					a0_wr[1996]    <= 0;                           
					a0_wr[1997]    <= 0;                           
					a0_wr[1998]    <= 0;                           
					a0_wr[1999]    <= 0;                           
					a0_wr[2000]    <= 0;                           
					a0_wr[2001]    <= 0;                           
					a0_wr[2002]    <= 0;                           
					a0_wr[2003]    <= 0;                           
					a0_wr[2004]    <= 0;                           
					a0_wr[2005]    <= 0;                           
					a0_wr[2006]    <= 0;                           
					a0_wr[2007]    <= 0;                           
					a0_wr[2008]    <= 0;                           
					a0_wr[2009]    <= 0;                           
					a0_wr[2010]    <= 0;                           
					a0_wr[2011]    <= 0;                           
					a0_wr[2012]    <= 0;                           
					a0_wr[2013]    <= 0;                           
					a0_wr[2014]    <= 0;                           
					a0_wr[2015]    <= 0;                           
					a0_wr[2016]    <= 0;                           
					a0_wr[2017]    <= 0;                           
					a0_wr[2018]    <= 0;                           
					a0_wr[2019]    <= 0;                           
					a0_wr[2020]    <= 0;                           
					a0_wr[2021]    <= 0;                           
					a0_wr[2022]    <= 0;                           
					a0_wr[2023]    <= 0;                           
					a0_wr[2024]    <= 0;                           
					a0_wr[2025]    <= 0;                           
					a0_wr[2026]    <= 0;                           
					a0_wr[2027]    <= 0;                           
					a0_wr[2028]    <= 0;                           
					a0_wr[2029]    <= 0;                           
					a0_wr[2030]    <= 0;                           
					a0_wr[2031]    <= 0;                           
					a0_wr[2032]    <= 0;                           
					a0_wr[2033]    <= 0;                           
					a0_wr[2034]    <= 0;                           
					a0_wr[2035]    <= 0;                           
					a0_wr[2036]    <= 0;                           
					a0_wr[2037]    <= 0;                           
					a0_wr[2038]    <= 0;                           
					a0_wr[2039]    <= 0;                           
					a0_wr[2040]    <= 0;                           
					a0_wr[2041]    <= 0;                           
					a0_wr[2042]    <= 0;                           
					a0_wr[2043]    <= 0;                           
					a0_wr[2044]    <= 0;                           
					a0_wr[2045]    <= 0;                           
					a0_wr[2046]    <= 0;                           
					a0_wr[2047]    <= 0;                           
				end
				else begin
					if (!stall) begin
						a0_wr[0]      <= x0_in;                       
						a0_wr[1]      <= x1_in;                       
						a0_wr[2]      <= x2_in;                       
						a0_wr[3]      <= x3_in;                       
						a0_wr[4]      <= x4_in;                       
						a0_wr[5]      <= x5_in;                       
						a0_wr[6]      <= x6_in;                       
						a0_wr[7]      <= x7_in;                       
						a0_wr[8]      <= x8_in;                       
						a0_wr[9]      <= x9_in;                       
						a0_wr[10]     <= x10_in;                      
						a0_wr[11]     <= x11_in;                      
						a0_wr[12]     <= x12_in;                      
						a0_wr[13]     <= x13_in;                      
						a0_wr[14]     <= x14_in;                      
						a0_wr[15]     <= x15_in;                      
						a0_wr[16]     <= x16_in;                      
						a0_wr[17]     <= x17_in;                      
						a0_wr[18]     <= x18_in;                      
						a0_wr[19]     <= x19_in;                      
						a0_wr[20]     <= x20_in;                      
						a0_wr[21]     <= x21_in;                      
						a0_wr[22]     <= x22_in;                      
						a0_wr[23]     <= x23_in;                      
						a0_wr[24]     <= x24_in;                      
						a0_wr[25]     <= x25_in;                      
						a0_wr[26]     <= x26_in;                      
						a0_wr[27]     <= x27_in;                      
						a0_wr[28]     <= x28_in;                      
						a0_wr[29]     <= x29_in;                      
						a0_wr[30]     <= x30_in;                      
						a0_wr[31]     <= x31_in;                      
						a0_wr[32]     <= x32_in;                      
						a0_wr[33]     <= x33_in;                      
						a0_wr[34]     <= x34_in;                      
						a0_wr[35]     <= x35_in;                      
						a0_wr[36]     <= x36_in;                      
						a0_wr[37]     <= x37_in;                      
						a0_wr[38]     <= x38_in;                      
						a0_wr[39]     <= x39_in;                      
						a0_wr[40]     <= x40_in;                      
						a0_wr[41]     <= x41_in;                      
						a0_wr[42]     <= x42_in;                      
						a0_wr[43]     <= x43_in;                      
						a0_wr[44]     <= x44_in;                      
						a0_wr[45]     <= x45_in;                      
						a0_wr[46]     <= x46_in;                      
						a0_wr[47]     <= x47_in;                      
						a0_wr[48]     <= x48_in;                      
						a0_wr[49]     <= x49_in;                      
						a0_wr[50]     <= x50_in;                      
						a0_wr[51]     <= x51_in;                      
						a0_wr[52]     <= x52_in;                      
						a0_wr[53]     <= x53_in;                      
						a0_wr[54]     <= x54_in;                      
						a0_wr[55]     <= x55_in;                      
						a0_wr[56]     <= x56_in;                      
						a0_wr[57]     <= x57_in;                      
						a0_wr[58]     <= x58_in;                      
						a0_wr[59]     <= x59_in;                      
						a0_wr[60]     <= x60_in;                      
						a0_wr[61]     <= x61_in;                      
						a0_wr[62]     <= x62_in;                      
						a0_wr[63]     <= x63_in;                      
						a0_wr[64]     <= x64_in;                      
						a0_wr[65]     <= x65_in;                      
						a0_wr[66]     <= x66_in;                      
						a0_wr[67]     <= x67_in;                      
						a0_wr[68]     <= x68_in;                      
						a0_wr[69]     <= x69_in;                      
						a0_wr[70]     <= x70_in;                      
						a0_wr[71]     <= x71_in;                      
						a0_wr[72]     <= x72_in;                      
						a0_wr[73]     <= x73_in;                      
						a0_wr[74]     <= x74_in;                      
						a0_wr[75]     <= x75_in;                      
						a0_wr[76]     <= x76_in;                      
						a0_wr[77]     <= x77_in;                      
						a0_wr[78]     <= x78_in;                      
						a0_wr[79]     <= x79_in;                      
						a0_wr[80]     <= x80_in;                      
						a0_wr[81]     <= x81_in;                      
						a0_wr[82]     <= x82_in;                      
						a0_wr[83]     <= x83_in;                      
						a0_wr[84]     <= x84_in;                      
						a0_wr[85]     <= x85_in;                      
						a0_wr[86]     <= x86_in;                      
						a0_wr[87]     <= x87_in;                      
						a0_wr[88]     <= x88_in;                      
						a0_wr[89]     <= x89_in;                      
						a0_wr[90]     <= x90_in;                      
						a0_wr[91]     <= x91_in;                      
						a0_wr[92]     <= x92_in;                      
						a0_wr[93]     <= x93_in;                      
						a0_wr[94]     <= x94_in;                      
						a0_wr[95]     <= x95_in;                      
						a0_wr[96]     <= x96_in;                      
						a0_wr[97]     <= x97_in;                      
						a0_wr[98]     <= x98_in;                      
						a0_wr[99]     <= x99_in;                      
						a0_wr[100]    <= x100_in;                     
						a0_wr[101]    <= x101_in;                     
						a0_wr[102]    <= x102_in;                     
						a0_wr[103]    <= x103_in;                     
						a0_wr[104]    <= x104_in;                     
						a0_wr[105]    <= x105_in;                     
						a0_wr[106]    <= x106_in;                     
						a0_wr[107]    <= x107_in;                     
						a0_wr[108]    <= x108_in;                     
						a0_wr[109]    <= x109_in;                     
						a0_wr[110]    <= x110_in;                     
						a0_wr[111]    <= x111_in;                     
						a0_wr[112]    <= x112_in;                     
						a0_wr[113]    <= x113_in;                     
						a0_wr[114]    <= x114_in;                     
						a0_wr[115]    <= x115_in;                     
						a0_wr[116]    <= x116_in;                     
						a0_wr[117]    <= x117_in;                     
						a0_wr[118]    <= x118_in;                     
						a0_wr[119]    <= x119_in;                     
						a0_wr[120]    <= x120_in;                     
						a0_wr[121]    <= x121_in;                     
						a0_wr[122]    <= x122_in;                     
						a0_wr[123]    <= x123_in;                     
						a0_wr[124]    <= x124_in;                     
						a0_wr[125]    <= x125_in;                     
						a0_wr[126]    <= x126_in;                     
						a0_wr[127]    <= x127_in;                     
						a0_wr[128]    <= x128_in;                     
						a0_wr[129]    <= x129_in;                     
						a0_wr[130]    <= x130_in;                     
						a0_wr[131]    <= x131_in;                     
						a0_wr[132]    <= x132_in;                     
						a0_wr[133]    <= x133_in;                     
						a0_wr[134]    <= x134_in;                     
						a0_wr[135]    <= x135_in;                     
						a0_wr[136]    <= x136_in;                     
						a0_wr[137]    <= x137_in;                     
						a0_wr[138]    <= x138_in;                     
						a0_wr[139]    <= x139_in;                     
						a0_wr[140]    <= x140_in;                     
						a0_wr[141]    <= x141_in;                     
						a0_wr[142]    <= x142_in;                     
						a0_wr[143]    <= x143_in;                     
						a0_wr[144]    <= x144_in;                     
						a0_wr[145]    <= x145_in;                     
						a0_wr[146]    <= x146_in;                     
						a0_wr[147]    <= x147_in;                     
						a0_wr[148]    <= x148_in;                     
						a0_wr[149]    <= x149_in;                     
						a0_wr[150]    <= x150_in;                     
						a0_wr[151]    <= x151_in;                     
						a0_wr[152]    <= x152_in;                     
						a0_wr[153]    <= x153_in;                     
						a0_wr[154]    <= x154_in;                     
						a0_wr[155]    <= x155_in;                     
						a0_wr[156]    <= x156_in;                     
						a0_wr[157]    <= x157_in;                     
						a0_wr[158]    <= x158_in;                     
						a0_wr[159]    <= x159_in;                     
						a0_wr[160]    <= x160_in;                     
						a0_wr[161]    <= x161_in;                     
						a0_wr[162]    <= x162_in;                     
						a0_wr[163]    <= x163_in;                     
						a0_wr[164]    <= x164_in;                     
						a0_wr[165]    <= x165_in;                     
						a0_wr[166]    <= x166_in;                     
						a0_wr[167]    <= x167_in;                     
						a0_wr[168]    <= x168_in;                     
						a0_wr[169]    <= x169_in;                     
						a0_wr[170]    <= x170_in;                     
						a0_wr[171]    <= x171_in;                     
						a0_wr[172]    <= x172_in;                     
						a0_wr[173]    <= x173_in;                     
						a0_wr[174]    <= x174_in;                     
						a0_wr[175]    <= x175_in;                     
						a0_wr[176]    <= x176_in;                     
						a0_wr[177]    <= x177_in;                     
						a0_wr[178]    <= x178_in;                     
						a0_wr[179]    <= x179_in;                     
						a0_wr[180]    <= x180_in;                     
						a0_wr[181]    <= x181_in;                     
						a0_wr[182]    <= x182_in;                     
						a0_wr[183]    <= x183_in;                     
						a0_wr[184]    <= x184_in;                     
						a0_wr[185]    <= x185_in;                     
						a0_wr[186]    <= x186_in;                     
						a0_wr[187]    <= x187_in;                     
						a0_wr[188]    <= x188_in;                     
						a0_wr[189]    <= x189_in;                     
						a0_wr[190]    <= x190_in;                     
						a0_wr[191]    <= x191_in;                     
						a0_wr[192]    <= x192_in;                     
						a0_wr[193]    <= x193_in;                     
						a0_wr[194]    <= x194_in;                     
						a0_wr[195]    <= x195_in;                     
						a0_wr[196]    <= x196_in;                     
						a0_wr[197]    <= x197_in;                     
						a0_wr[198]    <= x198_in;                     
						a0_wr[199]    <= x199_in;                     
						a0_wr[200]    <= x200_in;                     
						a0_wr[201]    <= x201_in;                     
						a0_wr[202]    <= x202_in;                     
						a0_wr[203]    <= x203_in;                     
						a0_wr[204]    <= x204_in;                     
						a0_wr[205]    <= x205_in;                     
						a0_wr[206]    <= x206_in;                     
						a0_wr[207]    <= x207_in;                     
						a0_wr[208]    <= x208_in;                     
						a0_wr[209]    <= x209_in;                     
						a0_wr[210]    <= x210_in;                     
						a0_wr[211]    <= x211_in;                     
						a0_wr[212]    <= x212_in;                     
						a0_wr[213]    <= x213_in;                     
						a0_wr[214]    <= x214_in;                     
						a0_wr[215]    <= x215_in;                     
						a0_wr[216]    <= x216_in;                     
						a0_wr[217]    <= x217_in;                     
						a0_wr[218]    <= x218_in;                     
						a0_wr[219]    <= x219_in;                     
						a0_wr[220]    <= x220_in;                     
						a0_wr[221]    <= x221_in;                     
						a0_wr[222]    <= x222_in;                     
						a0_wr[223]    <= x223_in;                     
						a0_wr[224]    <= x224_in;                     
						a0_wr[225]    <= x225_in;                     
						a0_wr[226]    <= x226_in;                     
						a0_wr[227]    <= x227_in;                     
						a0_wr[228]    <= x228_in;                     
						a0_wr[229]    <= x229_in;                     
						a0_wr[230]    <= x230_in;                     
						a0_wr[231]    <= x231_in;                     
						a0_wr[232]    <= x232_in;                     
						a0_wr[233]    <= x233_in;                     
						a0_wr[234]    <= x234_in;                     
						a0_wr[235]    <= x235_in;                     
						a0_wr[236]    <= x236_in;                     
						a0_wr[237]    <= x237_in;                     
						a0_wr[238]    <= x238_in;                     
						a0_wr[239]    <= x239_in;                     
						a0_wr[240]    <= x240_in;                     
						a0_wr[241]    <= x241_in;                     
						a0_wr[242]    <= x242_in;                     
						a0_wr[243]    <= x243_in;                     
						a0_wr[244]    <= x244_in;                     
						a0_wr[245]    <= x245_in;                     
						a0_wr[246]    <= x246_in;                     
						a0_wr[247]    <= x247_in;                     
						a0_wr[248]    <= x248_in;                     
						a0_wr[249]    <= x249_in;                     
						a0_wr[250]    <= x250_in;                     
						a0_wr[251]    <= x251_in;                     
						a0_wr[252]    <= x252_in;                     
						a0_wr[253]    <= x253_in;                     
						a0_wr[254]    <= x254_in;                     
						a0_wr[255]    <= x255_in;                     
						a0_wr[256]    <= x256_in;                     
						a0_wr[257]    <= x257_in;                     
						a0_wr[258]    <= x258_in;                     
						a0_wr[259]    <= x259_in;                     
						a0_wr[260]    <= x260_in;                     
						a0_wr[261]    <= x261_in;                     
						a0_wr[262]    <= x262_in;                     
						a0_wr[263]    <= x263_in;                     
						a0_wr[264]    <= x264_in;                     
						a0_wr[265]    <= x265_in;                     
						a0_wr[266]    <= x266_in;                     
						a0_wr[267]    <= x267_in;                     
						a0_wr[268]    <= x268_in;                     
						a0_wr[269]    <= x269_in;                     
						a0_wr[270]    <= x270_in;                     
						a0_wr[271]    <= x271_in;                     
						a0_wr[272]    <= x272_in;                     
						a0_wr[273]    <= x273_in;                     
						a0_wr[274]    <= x274_in;                     
						a0_wr[275]    <= x275_in;                     
						a0_wr[276]    <= x276_in;                     
						a0_wr[277]    <= x277_in;                     
						a0_wr[278]    <= x278_in;                     
						a0_wr[279]    <= x279_in;                     
						a0_wr[280]    <= x280_in;                     
						a0_wr[281]    <= x281_in;                     
						a0_wr[282]    <= x282_in;                     
						a0_wr[283]    <= x283_in;                     
						a0_wr[284]    <= x284_in;                     
						a0_wr[285]    <= x285_in;                     
						a0_wr[286]    <= x286_in;                     
						a0_wr[287]    <= x287_in;                     
						a0_wr[288]    <= x288_in;                     
						a0_wr[289]    <= x289_in;                     
						a0_wr[290]    <= x290_in;                     
						a0_wr[291]    <= x291_in;                     
						a0_wr[292]    <= x292_in;                     
						a0_wr[293]    <= x293_in;                     
						a0_wr[294]    <= x294_in;                     
						a0_wr[295]    <= x295_in;                     
						a0_wr[296]    <= x296_in;                     
						a0_wr[297]    <= x297_in;                     
						a0_wr[298]    <= x298_in;                     
						a0_wr[299]    <= x299_in;                     
						a0_wr[300]    <= x300_in;                     
						a0_wr[301]    <= x301_in;                     
						a0_wr[302]    <= x302_in;                     
						a0_wr[303]    <= x303_in;                     
						a0_wr[304]    <= x304_in;                     
						a0_wr[305]    <= x305_in;                     
						a0_wr[306]    <= x306_in;                     
						a0_wr[307]    <= x307_in;                     
						a0_wr[308]    <= x308_in;                     
						a0_wr[309]    <= x309_in;                     
						a0_wr[310]    <= x310_in;                     
						a0_wr[311]    <= x311_in;                     
						a0_wr[312]    <= x312_in;                     
						a0_wr[313]    <= x313_in;                     
						a0_wr[314]    <= x314_in;                     
						a0_wr[315]    <= x315_in;                     
						a0_wr[316]    <= x316_in;                     
						a0_wr[317]    <= x317_in;                     
						a0_wr[318]    <= x318_in;                     
						a0_wr[319]    <= x319_in;                     
						a0_wr[320]    <= x320_in;                     
						a0_wr[321]    <= x321_in;                     
						a0_wr[322]    <= x322_in;                     
						a0_wr[323]    <= x323_in;                     
						a0_wr[324]    <= x324_in;                     
						a0_wr[325]    <= x325_in;                     
						a0_wr[326]    <= x326_in;                     
						a0_wr[327]    <= x327_in;                     
						a0_wr[328]    <= x328_in;                     
						a0_wr[329]    <= x329_in;                     
						a0_wr[330]    <= x330_in;                     
						a0_wr[331]    <= x331_in;                     
						a0_wr[332]    <= x332_in;                     
						a0_wr[333]    <= x333_in;                     
						a0_wr[334]    <= x334_in;                     
						a0_wr[335]    <= x335_in;                     
						a0_wr[336]    <= x336_in;                     
						a0_wr[337]    <= x337_in;                     
						a0_wr[338]    <= x338_in;                     
						a0_wr[339]    <= x339_in;                     
						a0_wr[340]    <= x340_in;                     
						a0_wr[341]    <= x341_in;                     
						a0_wr[342]    <= x342_in;                     
						a0_wr[343]    <= x343_in;                     
						a0_wr[344]    <= x344_in;                     
						a0_wr[345]    <= x345_in;                     
						a0_wr[346]    <= x346_in;                     
						a0_wr[347]    <= x347_in;                     
						a0_wr[348]    <= x348_in;                     
						a0_wr[349]    <= x349_in;                     
						a0_wr[350]    <= x350_in;                     
						a0_wr[351]    <= x351_in;                     
						a0_wr[352]    <= x352_in;                     
						a0_wr[353]    <= x353_in;                     
						a0_wr[354]    <= x354_in;                     
						a0_wr[355]    <= x355_in;                     
						a0_wr[356]    <= x356_in;                     
						a0_wr[357]    <= x357_in;                     
						a0_wr[358]    <= x358_in;                     
						a0_wr[359]    <= x359_in;                     
						a0_wr[360]    <= x360_in;                     
						a0_wr[361]    <= x361_in;                     
						a0_wr[362]    <= x362_in;                     
						a0_wr[363]    <= x363_in;                     
						a0_wr[364]    <= x364_in;                     
						a0_wr[365]    <= x365_in;                     
						a0_wr[366]    <= x366_in;                     
						a0_wr[367]    <= x367_in;                     
						a0_wr[368]    <= x368_in;                     
						a0_wr[369]    <= x369_in;                     
						a0_wr[370]    <= x370_in;                     
						a0_wr[371]    <= x371_in;                     
						a0_wr[372]    <= x372_in;                     
						a0_wr[373]    <= x373_in;                     
						a0_wr[374]    <= x374_in;                     
						a0_wr[375]    <= x375_in;                     
						a0_wr[376]    <= x376_in;                     
						a0_wr[377]    <= x377_in;                     
						a0_wr[378]    <= x378_in;                     
						a0_wr[379]    <= x379_in;                     
						a0_wr[380]    <= x380_in;                     
						a0_wr[381]    <= x381_in;                     
						a0_wr[382]    <= x382_in;                     
						a0_wr[383]    <= x383_in;                     
						a0_wr[384]    <= x384_in;                     
						a0_wr[385]    <= x385_in;                     
						a0_wr[386]    <= x386_in;                     
						a0_wr[387]    <= x387_in;                     
						a0_wr[388]    <= x388_in;                     
						a0_wr[389]    <= x389_in;                     
						a0_wr[390]    <= x390_in;                     
						a0_wr[391]    <= x391_in;                     
						a0_wr[392]    <= x392_in;                     
						a0_wr[393]    <= x393_in;                     
						a0_wr[394]    <= x394_in;                     
						a0_wr[395]    <= x395_in;                     
						a0_wr[396]    <= x396_in;                     
						a0_wr[397]    <= x397_in;                     
						a0_wr[398]    <= x398_in;                     
						a0_wr[399]    <= x399_in;                     
						a0_wr[400]    <= x400_in;                     
						a0_wr[401]    <= x401_in;                     
						a0_wr[402]    <= x402_in;                     
						a0_wr[403]    <= x403_in;                     
						a0_wr[404]    <= x404_in;                     
						a0_wr[405]    <= x405_in;                     
						a0_wr[406]    <= x406_in;                     
						a0_wr[407]    <= x407_in;                     
						a0_wr[408]    <= x408_in;                     
						a0_wr[409]    <= x409_in;                     
						a0_wr[410]    <= x410_in;                     
						a0_wr[411]    <= x411_in;                     
						a0_wr[412]    <= x412_in;                     
						a0_wr[413]    <= x413_in;                     
						a0_wr[414]    <= x414_in;                     
						a0_wr[415]    <= x415_in;                     
						a0_wr[416]    <= x416_in;                     
						a0_wr[417]    <= x417_in;                     
						a0_wr[418]    <= x418_in;                     
						a0_wr[419]    <= x419_in;                     
						a0_wr[420]    <= x420_in;                     
						a0_wr[421]    <= x421_in;                     
						a0_wr[422]    <= x422_in;                     
						a0_wr[423]    <= x423_in;                     
						a0_wr[424]    <= x424_in;                     
						a0_wr[425]    <= x425_in;                     
						a0_wr[426]    <= x426_in;                     
						a0_wr[427]    <= x427_in;                     
						a0_wr[428]    <= x428_in;                     
						a0_wr[429]    <= x429_in;                     
						a0_wr[430]    <= x430_in;                     
						a0_wr[431]    <= x431_in;                     
						a0_wr[432]    <= x432_in;                     
						a0_wr[433]    <= x433_in;                     
						a0_wr[434]    <= x434_in;                     
						a0_wr[435]    <= x435_in;                     
						a0_wr[436]    <= x436_in;                     
						a0_wr[437]    <= x437_in;                     
						a0_wr[438]    <= x438_in;                     
						a0_wr[439]    <= x439_in;                     
						a0_wr[440]    <= x440_in;                     
						a0_wr[441]    <= x441_in;                     
						a0_wr[442]    <= x442_in;                     
						a0_wr[443]    <= x443_in;                     
						a0_wr[444]    <= x444_in;                     
						a0_wr[445]    <= x445_in;                     
						a0_wr[446]    <= x446_in;                     
						a0_wr[447]    <= x447_in;                     
						a0_wr[448]    <= x448_in;                     
						a0_wr[449]    <= x449_in;                     
						a0_wr[450]    <= x450_in;                     
						a0_wr[451]    <= x451_in;                     
						a0_wr[452]    <= x452_in;                     
						a0_wr[453]    <= x453_in;                     
						a0_wr[454]    <= x454_in;                     
						a0_wr[455]    <= x455_in;                     
						a0_wr[456]    <= x456_in;                     
						a0_wr[457]    <= x457_in;                     
						a0_wr[458]    <= x458_in;                     
						a0_wr[459]    <= x459_in;                     
						a0_wr[460]    <= x460_in;                     
						a0_wr[461]    <= x461_in;                     
						a0_wr[462]    <= x462_in;                     
						a0_wr[463]    <= x463_in;                     
						a0_wr[464]    <= x464_in;                     
						a0_wr[465]    <= x465_in;                     
						a0_wr[466]    <= x466_in;                     
						a0_wr[467]    <= x467_in;                     
						a0_wr[468]    <= x468_in;                     
						a0_wr[469]    <= x469_in;                     
						a0_wr[470]    <= x470_in;                     
						a0_wr[471]    <= x471_in;                     
						a0_wr[472]    <= x472_in;                     
						a0_wr[473]    <= x473_in;                     
						a0_wr[474]    <= x474_in;                     
						a0_wr[475]    <= x475_in;                     
						a0_wr[476]    <= x476_in;                     
						a0_wr[477]    <= x477_in;                     
						a0_wr[478]    <= x478_in;                     
						a0_wr[479]    <= x479_in;                     
						a0_wr[480]    <= x480_in;                     
						a0_wr[481]    <= x481_in;                     
						a0_wr[482]    <= x482_in;                     
						a0_wr[483]    <= x483_in;                     
						a0_wr[484]    <= x484_in;                     
						a0_wr[485]    <= x485_in;                     
						a0_wr[486]    <= x486_in;                     
						a0_wr[487]    <= x487_in;                     
						a0_wr[488]    <= x488_in;                     
						a0_wr[489]    <= x489_in;                     
						a0_wr[490]    <= x490_in;                     
						a0_wr[491]    <= x491_in;                     
						a0_wr[492]    <= x492_in;                     
						a0_wr[493]    <= x493_in;                     
						a0_wr[494]    <= x494_in;                     
						a0_wr[495]    <= x495_in;                     
						a0_wr[496]    <= x496_in;                     
						a0_wr[497]    <= x497_in;                     
						a0_wr[498]    <= x498_in;                     
						a0_wr[499]    <= x499_in;                     
						a0_wr[500]    <= x500_in;                     
						a0_wr[501]    <= x501_in;                     
						a0_wr[502]    <= x502_in;                     
						a0_wr[503]    <= x503_in;                     
						a0_wr[504]    <= x504_in;                     
						a0_wr[505]    <= x505_in;                     
						a0_wr[506]    <= x506_in;                     
						a0_wr[507]    <= x507_in;                     
						a0_wr[508]    <= x508_in;                     
						a0_wr[509]    <= x509_in;                     
						a0_wr[510]    <= x510_in;                     
						a0_wr[511]    <= x511_in;                     
						a0_wr[512]    <= x512_in;                     
						a0_wr[513]    <= x513_in;                     
						a0_wr[514]    <= x514_in;                     
						a0_wr[515]    <= x515_in;                     
						a0_wr[516]    <= x516_in;                     
						a0_wr[517]    <= x517_in;                     
						a0_wr[518]    <= x518_in;                     
						a0_wr[519]    <= x519_in;                     
						a0_wr[520]    <= x520_in;                     
						a0_wr[521]    <= x521_in;                     
						a0_wr[522]    <= x522_in;                     
						a0_wr[523]    <= x523_in;                     
						a0_wr[524]    <= x524_in;                     
						a0_wr[525]    <= x525_in;                     
						a0_wr[526]    <= x526_in;                     
						a0_wr[527]    <= x527_in;                     
						a0_wr[528]    <= x528_in;                     
						a0_wr[529]    <= x529_in;                     
						a0_wr[530]    <= x530_in;                     
						a0_wr[531]    <= x531_in;                     
						a0_wr[532]    <= x532_in;                     
						a0_wr[533]    <= x533_in;                     
						a0_wr[534]    <= x534_in;                     
						a0_wr[535]    <= x535_in;                     
						a0_wr[536]    <= x536_in;                     
						a0_wr[537]    <= x537_in;                     
						a0_wr[538]    <= x538_in;                     
						a0_wr[539]    <= x539_in;                     
						a0_wr[540]    <= x540_in;                     
						a0_wr[541]    <= x541_in;                     
						a0_wr[542]    <= x542_in;                     
						a0_wr[543]    <= x543_in;                     
						a0_wr[544]    <= x544_in;                     
						a0_wr[545]    <= x545_in;                     
						a0_wr[546]    <= x546_in;                     
						a0_wr[547]    <= x547_in;                     
						a0_wr[548]    <= x548_in;                     
						a0_wr[549]    <= x549_in;                     
						a0_wr[550]    <= x550_in;                     
						a0_wr[551]    <= x551_in;                     
						a0_wr[552]    <= x552_in;                     
						a0_wr[553]    <= x553_in;                     
						a0_wr[554]    <= x554_in;                     
						a0_wr[555]    <= x555_in;                     
						a0_wr[556]    <= x556_in;                     
						a0_wr[557]    <= x557_in;                     
						a0_wr[558]    <= x558_in;                     
						a0_wr[559]    <= x559_in;                     
						a0_wr[560]    <= x560_in;                     
						a0_wr[561]    <= x561_in;                     
						a0_wr[562]    <= x562_in;                     
						a0_wr[563]    <= x563_in;                     
						a0_wr[564]    <= x564_in;                     
						a0_wr[565]    <= x565_in;                     
						a0_wr[566]    <= x566_in;                     
						a0_wr[567]    <= x567_in;                     
						a0_wr[568]    <= x568_in;                     
						a0_wr[569]    <= x569_in;                     
						a0_wr[570]    <= x570_in;                     
						a0_wr[571]    <= x571_in;                     
						a0_wr[572]    <= x572_in;                     
						a0_wr[573]    <= x573_in;                     
						a0_wr[574]    <= x574_in;                     
						a0_wr[575]    <= x575_in;                     
						a0_wr[576]    <= x576_in;                     
						a0_wr[577]    <= x577_in;                     
						a0_wr[578]    <= x578_in;                     
						a0_wr[579]    <= x579_in;                     
						a0_wr[580]    <= x580_in;                     
						a0_wr[581]    <= x581_in;                     
						a0_wr[582]    <= x582_in;                     
						a0_wr[583]    <= x583_in;                     
						a0_wr[584]    <= x584_in;                     
						a0_wr[585]    <= x585_in;                     
						a0_wr[586]    <= x586_in;                     
						a0_wr[587]    <= x587_in;                     
						a0_wr[588]    <= x588_in;                     
						a0_wr[589]    <= x589_in;                     
						a0_wr[590]    <= x590_in;                     
						a0_wr[591]    <= x591_in;                     
						a0_wr[592]    <= x592_in;                     
						a0_wr[593]    <= x593_in;                     
						a0_wr[594]    <= x594_in;                     
						a0_wr[595]    <= x595_in;                     
						a0_wr[596]    <= x596_in;                     
						a0_wr[597]    <= x597_in;                     
						a0_wr[598]    <= x598_in;                     
						a0_wr[599]    <= x599_in;                     
						a0_wr[600]    <= x600_in;                     
						a0_wr[601]    <= x601_in;                     
						a0_wr[602]    <= x602_in;                     
						a0_wr[603]    <= x603_in;                     
						a0_wr[604]    <= x604_in;                     
						a0_wr[605]    <= x605_in;                     
						a0_wr[606]    <= x606_in;                     
						a0_wr[607]    <= x607_in;                     
						a0_wr[608]    <= x608_in;                     
						a0_wr[609]    <= x609_in;                     
						a0_wr[610]    <= x610_in;                     
						a0_wr[611]    <= x611_in;                     
						a0_wr[612]    <= x612_in;                     
						a0_wr[613]    <= x613_in;                     
						a0_wr[614]    <= x614_in;                     
						a0_wr[615]    <= x615_in;                     
						a0_wr[616]    <= x616_in;                     
						a0_wr[617]    <= x617_in;                     
						a0_wr[618]    <= x618_in;                     
						a0_wr[619]    <= x619_in;                     
						a0_wr[620]    <= x620_in;                     
						a0_wr[621]    <= x621_in;                     
						a0_wr[622]    <= x622_in;                     
						a0_wr[623]    <= x623_in;                     
						a0_wr[624]    <= x624_in;                     
						a0_wr[625]    <= x625_in;                     
						a0_wr[626]    <= x626_in;                     
						a0_wr[627]    <= x627_in;                     
						a0_wr[628]    <= x628_in;                     
						a0_wr[629]    <= x629_in;                     
						a0_wr[630]    <= x630_in;                     
						a0_wr[631]    <= x631_in;                     
						a0_wr[632]    <= x632_in;                     
						a0_wr[633]    <= x633_in;                     
						a0_wr[634]    <= x634_in;                     
						a0_wr[635]    <= x635_in;                     
						a0_wr[636]    <= x636_in;                     
						a0_wr[637]    <= x637_in;                     
						a0_wr[638]    <= x638_in;                     
						a0_wr[639]    <= x639_in;                     
						a0_wr[640]    <= x640_in;                     
						a0_wr[641]    <= x641_in;                     
						a0_wr[642]    <= x642_in;                     
						a0_wr[643]    <= x643_in;                     
						a0_wr[644]    <= x644_in;                     
						a0_wr[645]    <= x645_in;                     
						a0_wr[646]    <= x646_in;                     
						a0_wr[647]    <= x647_in;                     
						a0_wr[648]    <= x648_in;                     
						a0_wr[649]    <= x649_in;                     
						a0_wr[650]    <= x650_in;                     
						a0_wr[651]    <= x651_in;                     
						a0_wr[652]    <= x652_in;                     
						a0_wr[653]    <= x653_in;                     
						a0_wr[654]    <= x654_in;                     
						a0_wr[655]    <= x655_in;                     
						a0_wr[656]    <= x656_in;                     
						a0_wr[657]    <= x657_in;                     
						a0_wr[658]    <= x658_in;                     
						a0_wr[659]    <= x659_in;                     
						a0_wr[660]    <= x660_in;                     
						a0_wr[661]    <= x661_in;                     
						a0_wr[662]    <= x662_in;                     
						a0_wr[663]    <= x663_in;                     
						a0_wr[664]    <= x664_in;                     
						a0_wr[665]    <= x665_in;                     
						a0_wr[666]    <= x666_in;                     
						a0_wr[667]    <= x667_in;                     
						a0_wr[668]    <= x668_in;                     
						a0_wr[669]    <= x669_in;                     
						a0_wr[670]    <= x670_in;                     
						a0_wr[671]    <= x671_in;                     
						a0_wr[672]    <= x672_in;                     
						a0_wr[673]    <= x673_in;                     
						a0_wr[674]    <= x674_in;                     
						a0_wr[675]    <= x675_in;                     
						a0_wr[676]    <= x676_in;                     
						a0_wr[677]    <= x677_in;                     
						a0_wr[678]    <= x678_in;                     
						a0_wr[679]    <= x679_in;                     
						a0_wr[680]    <= x680_in;                     
						a0_wr[681]    <= x681_in;                     
						a0_wr[682]    <= x682_in;                     
						a0_wr[683]    <= x683_in;                     
						a0_wr[684]    <= x684_in;                     
						a0_wr[685]    <= x685_in;                     
						a0_wr[686]    <= x686_in;                     
						a0_wr[687]    <= x687_in;                     
						a0_wr[688]    <= x688_in;                     
						a0_wr[689]    <= x689_in;                     
						a0_wr[690]    <= x690_in;                     
						a0_wr[691]    <= x691_in;                     
						a0_wr[692]    <= x692_in;                     
						a0_wr[693]    <= x693_in;                     
						a0_wr[694]    <= x694_in;                     
						a0_wr[695]    <= x695_in;                     
						a0_wr[696]    <= x696_in;                     
						a0_wr[697]    <= x697_in;                     
						a0_wr[698]    <= x698_in;                     
						a0_wr[699]    <= x699_in;                     
						a0_wr[700]    <= x700_in;                     
						a0_wr[701]    <= x701_in;                     
						a0_wr[702]    <= x702_in;                     
						a0_wr[703]    <= x703_in;                     
						a0_wr[704]    <= x704_in;                     
						a0_wr[705]    <= x705_in;                     
						a0_wr[706]    <= x706_in;                     
						a0_wr[707]    <= x707_in;                     
						a0_wr[708]    <= x708_in;                     
						a0_wr[709]    <= x709_in;                     
						a0_wr[710]    <= x710_in;                     
						a0_wr[711]    <= x711_in;                     
						a0_wr[712]    <= x712_in;                     
						a0_wr[713]    <= x713_in;                     
						a0_wr[714]    <= x714_in;                     
						a0_wr[715]    <= x715_in;                     
						a0_wr[716]    <= x716_in;                     
						a0_wr[717]    <= x717_in;                     
						a0_wr[718]    <= x718_in;                     
						a0_wr[719]    <= x719_in;                     
						a0_wr[720]    <= x720_in;                     
						a0_wr[721]    <= x721_in;                     
						a0_wr[722]    <= x722_in;                     
						a0_wr[723]    <= x723_in;                     
						a0_wr[724]    <= x724_in;                     
						a0_wr[725]    <= x725_in;                     
						a0_wr[726]    <= x726_in;                     
						a0_wr[727]    <= x727_in;                     
						a0_wr[728]    <= x728_in;                     
						a0_wr[729]    <= x729_in;                     
						a0_wr[730]    <= x730_in;                     
						a0_wr[731]    <= x731_in;                     
						a0_wr[732]    <= x732_in;                     
						a0_wr[733]    <= x733_in;                     
						a0_wr[734]    <= x734_in;                     
						a0_wr[735]    <= x735_in;                     
						a0_wr[736]    <= x736_in;                     
						a0_wr[737]    <= x737_in;                     
						a0_wr[738]    <= x738_in;                     
						a0_wr[739]    <= x739_in;                     
						a0_wr[740]    <= x740_in;                     
						a0_wr[741]    <= x741_in;                     
						a0_wr[742]    <= x742_in;                     
						a0_wr[743]    <= x743_in;                     
						a0_wr[744]    <= x744_in;                     
						a0_wr[745]    <= x745_in;                     
						a0_wr[746]    <= x746_in;                     
						a0_wr[747]    <= x747_in;                     
						a0_wr[748]    <= x748_in;                     
						a0_wr[749]    <= x749_in;                     
						a0_wr[750]    <= x750_in;                     
						a0_wr[751]    <= x751_in;                     
						a0_wr[752]    <= x752_in;                     
						a0_wr[753]    <= x753_in;                     
						a0_wr[754]    <= x754_in;                     
						a0_wr[755]    <= x755_in;                     
						a0_wr[756]    <= x756_in;                     
						a0_wr[757]    <= x757_in;                     
						a0_wr[758]    <= x758_in;                     
						a0_wr[759]    <= x759_in;                     
						a0_wr[760]    <= x760_in;                     
						a0_wr[761]    <= x761_in;                     
						a0_wr[762]    <= x762_in;                     
						a0_wr[763]    <= x763_in;                     
						a0_wr[764]    <= x764_in;                     
						a0_wr[765]    <= x765_in;                     
						a0_wr[766]    <= x766_in;                     
						a0_wr[767]    <= x767_in;                     
						a0_wr[768]    <= x768_in;                     
						a0_wr[769]    <= x769_in;                     
						a0_wr[770]    <= x770_in;                     
						a0_wr[771]    <= x771_in;                     
						a0_wr[772]    <= x772_in;                     
						a0_wr[773]    <= x773_in;                     
						a0_wr[774]    <= x774_in;                     
						a0_wr[775]    <= x775_in;                     
						a0_wr[776]    <= x776_in;                     
						a0_wr[777]    <= x777_in;                     
						a0_wr[778]    <= x778_in;                     
						a0_wr[779]    <= x779_in;                     
						a0_wr[780]    <= x780_in;                     
						a0_wr[781]    <= x781_in;                     
						a0_wr[782]    <= x782_in;                     
						a0_wr[783]    <= x783_in;                     
						a0_wr[784]    <= x784_in;                     
						a0_wr[785]    <= x785_in;                     
						a0_wr[786]    <= x786_in;                     
						a0_wr[787]    <= x787_in;                     
						a0_wr[788]    <= x788_in;                     
						a0_wr[789]    <= x789_in;                     
						a0_wr[790]    <= x790_in;                     
						a0_wr[791]    <= x791_in;                     
						a0_wr[792]    <= x792_in;                     
						a0_wr[793]    <= x793_in;                     
						a0_wr[794]    <= x794_in;                     
						a0_wr[795]    <= x795_in;                     
						a0_wr[796]    <= x796_in;                     
						a0_wr[797]    <= x797_in;                     
						a0_wr[798]    <= x798_in;                     
						a0_wr[799]    <= x799_in;                     
						a0_wr[800]    <= x800_in;                     
						a0_wr[801]    <= x801_in;                     
						a0_wr[802]    <= x802_in;                     
						a0_wr[803]    <= x803_in;                     
						a0_wr[804]    <= x804_in;                     
						a0_wr[805]    <= x805_in;                     
						a0_wr[806]    <= x806_in;                     
						a0_wr[807]    <= x807_in;                     
						a0_wr[808]    <= x808_in;                     
						a0_wr[809]    <= x809_in;                     
						a0_wr[810]    <= x810_in;                     
						a0_wr[811]    <= x811_in;                     
						a0_wr[812]    <= x812_in;                     
						a0_wr[813]    <= x813_in;                     
						a0_wr[814]    <= x814_in;                     
						a0_wr[815]    <= x815_in;                     
						a0_wr[816]    <= x816_in;                     
						a0_wr[817]    <= x817_in;                     
						a0_wr[818]    <= x818_in;                     
						a0_wr[819]    <= x819_in;                     
						a0_wr[820]    <= x820_in;                     
						a0_wr[821]    <= x821_in;                     
						a0_wr[822]    <= x822_in;                     
						a0_wr[823]    <= x823_in;                     
						a0_wr[824]    <= x824_in;                     
						a0_wr[825]    <= x825_in;                     
						a0_wr[826]    <= x826_in;                     
						a0_wr[827]    <= x827_in;                     
						a0_wr[828]    <= x828_in;                     
						a0_wr[829]    <= x829_in;                     
						a0_wr[830]    <= x830_in;                     
						a0_wr[831]    <= x831_in;                     
						a0_wr[832]    <= x832_in;                     
						a0_wr[833]    <= x833_in;                     
						a0_wr[834]    <= x834_in;                     
						a0_wr[835]    <= x835_in;                     
						a0_wr[836]    <= x836_in;                     
						a0_wr[837]    <= x837_in;                     
						a0_wr[838]    <= x838_in;                     
						a0_wr[839]    <= x839_in;                     
						a0_wr[840]    <= x840_in;                     
						a0_wr[841]    <= x841_in;                     
						a0_wr[842]    <= x842_in;                     
						a0_wr[843]    <= x843_in;                     
						a0_wr[844]    <= x844_in;                     
						a0_wr[845]    <= x845_in;                     
						a0_wr[846]    <= x846_in;                     
						a0_wr[847]    <= x847_in;                     
						a0_wr[848]    <= x848_in;                     
						a0_wr[849]    <= x849_in;                     
						a0_wr[850]    <= x850_in;                     
						a0_wr[851]    <= x851_in;                     
						a0_wr[852]    <= x852_in;                     
						a0_wr[853]    <= x853_in;                     
						a0_wr[854]    <= x854_in;                     
						a0_wr[855]    <= x855_in;                     
						a0_wr[856]    <= x856_in;                     
						a0_wr[857]    <= x857_in;                     
						a0_wr[858]    <= x858_in;                     
						a0_wr[859]    <= x859_in;                     
						a0_wr[860]    <= x860_in;                     
						a0_wr[861]    <= x861_in;                     
						a0_wr[862]    <= x862_in;                     
						a0_wr[863]    <= x863_in;                     
						a0_wr[864]    <= x864_in;                     
						a0_wr[865]    <= x865_in;                     
						a0_wr[866]    <= x866_in;                     
						a0_wr[867]    <= x867_in;                     
						a0_wr[868]    <= x868_in;                     
						a0_wr[869]    <= x869_in;                     
						a0_wr[870]    <= x870_in;                     
						a0_wr[871]    <= x871_in;                     
						a0_wr[872]    <= x872_in;                     
						a0_wr[873]    <= x873_in;                     
						a0_wr[874]    <= x874_in;                     
						a0_wr[875]    <= x875_in;                     
						a0_wr[876]    <= x876_in;                     
						a0_wr[877]    <= x877_in;                     
						a0_wr[878]    <= x878_in;                     
						a0_wr[879]    <= x879_in;                     
						a0_wr[880]    <= x880_in;                     
						a0_wr[881]    <= x881_in;                     
						a0_wr[882]    <= x882_in;                     
						a0_wr[883]    <= x883_in;                     
						a0_wr[884]    <= x884_in;                     
						a0_wr[885]    <= x885_in;                     
						a0_wr[886]    <= x886_in;                     
						a0_wr[887]    <= x887_in;                     
						a0_wr[888]    <= x888_in;                     
						a0_wr[889]    <= x889_in;                     
						a0_wr[890]    <= x890_in;                     
						a0_wr[891]    <= x891_in;                     
						a0_wr[892]    <= x892_in;                     
						a0_wr[893]    <= x893_in;                     
						a0_wr[894]    <= x894_in;                     
						a0_wr[895]    <= x895_in;                     
						a0_wr[896]    <= x896_in;                     
						a0_wr[897]    <= x897_in;                     
						a0_wr[898]    <= x898_in;                     
						a0_wr[899]    <= x899_in;                     
						a0_wr[900]    <= x900_in;                     
						a0_wr[901]    <= x901_in;                     
						a0_wr[902]    <= x902_in;                     
						a0_wr[903]    <= x903_in;                     
						a0_wr[904]    <= x904_in;                     
						a0_wr[905]    <= x905_in;                     
						a0_wr[906]    <= x906_in;                     
						a0_wr[907]    <= x907_in;                     
						a0_wr[908]    <= x908_in;                     
						a0_wr[909]    <= x909_in;                     
						a0_wr[910]    <= x910_in;                     
						a0_wr[911]    <= x911_in;                     
						a0_wr[912]    <= x912_in;                     
						a0_wr[913]    <= x913_in;                     
						a0_wr[914]    <= x914_in;                     
						a0_wr[915]    <= x915_in;                     
						a0_wr[916]    <= x916_in;                     
						a0_wr[917]    <= x917_in;                     
						a0_wr[918]    <= x918_in;                     
						a0_wr[919]    <= x919_in;                     
						a0_wr[920]    <= x920_in;                     
						a0_wr[921]    <= x921_in;                     
						a0_wr[922]    <= x922_in;                     
						a0_wr[923]    <= x923_in;                     
						a0_wr[924]    <= x924_in;                     
						a0_wr[925]    <= x925_in;                     
						a0_wr[926]    <= x926_in;                     
						a0_wr[927]    <= x927_in;                     
						a0_wr[928]    <= x928_in;                     
						a0_wr[929]    <= x929_in;                     
						a0_wr[930]    <= x930_in;                     
						a0_wr[931]    <= x931_in;                     
						a0_wr[932]    <= x932_in;                     
						a0_wr[933]    <= x933_in;                     
						a0_wr[934]    <= x934_in;                     
						a0_wr[935]    <= x935_in;                     
						a0_wr[936]    <= x936_in;                     
						a0_wr[937]    <= x937_in;                     
						a0_wr[938]    <= x938_in;                     
						a0_wr[939]    <= x939_in;                     
						a0_wr[940]    <= x940_in;                     
						a0_wr[941]    <= x941_in;                     
						a0_wr[942]    <= x942_in;                     
						a0_wr[943]    <= x943_in;                     
						a0_wr[944]    <= x944_in;                     
						a0_wr[945]    <= x945_in;                     
						a0_wr[946]    <= x946_in;                     
						a0_wr[947]    <= x947_in;                     
						a0_wr[948]    <= x948_in;                     
						a0_wr[949]    <= x949_in;                     
						a0_wr[950]    <= x950_in;                     
						a0_wr[951]    <= x951_in;                     
						a0_wr[952]    <= x952_in;                     
						a0_wr[953]    <= x953_in;                     
						a0_wr[954]    <= x954_in;                     
						a0_wr[955]    <= x955_in;                     
						a0_wr[956]    <= x956_in;                     
						a0_wr[957]    <= x957_in;                     
						a0_wr[958]    <= x958_in;                     
						a0_wr[959]    <= x959_in;                     
						a0_wr[960]    <= x960_in;                     
						a0_wr[961]    <= x961_in;                     
						a0_wr[962]    <= x962_in;                     
						a0_wr[963]    <= x963_in;                     
						a0_wr[964]    <= x964_in;                     
						a0_wr[965]    <= x965_in;                     
						a0_wr[966]    <= x966_in;                     
						a0_wr[967]    <= x967_in;                     
						a0_wr[968]    <= x968_in;                     
						a0_wr[969]    <= x969_in;                     
						a0_wr[970]    <= x970_in;                     
						a0_wr[971]    <= x971_in;                     
						a0_wr[972]    <= x972_in;                     
						a0_wr[973]    <= x973_in;                     
						a0_wr[974]    <= x974_in;                     
						a0_wr[975]    <= x975_in;                     
						a0_wr[976]    <= x976_in;                     
						a0_wr[977]    <= x977_in;                     
						a0_wr[978]    <= x978_in;                     
						a0_wr[979]    <= x979_in;                     
						a0_wr[980]    <= x980_in;                     
						a0_wr[981]    <= x981_in;                     
						a0_wr[982]    <= x982_in;                     
						a0_wr[983]    <= x983_in;                     
						a0_wr[984]    <= x984_in;                     
						a0_wr[985]    <= x985_in;                     
						a0_wr[986]    <= x986_in;                     
						a0_wr[987]    <= x987_in;                     
						a0_wr[988]    <= x988_in;                     
						a0_wr[989]    <= x989_in;                     
						a0_wr[990]    <= x990_in;                     
						a0_wr[991]    <= x991_in;                     
						a0_wr[992]    <= x992_in;                     
						a0_wr[993]    <= x993_in;                     
						a0_wr[994]    <= x994_in;                     
						a0_wr[995]    <= x995_in;                     
						a0_wr[996]    <= x996_in;                     
						a0_wr[997]    <= x997_in;                     
						a0_wr[998]    <= x998_in;                     
						a0_wr[999]    <= x999_in;                     
						a0_wr[1000]   <= x1000_in;                    
						a0_wr[1001]   <= x1001_in;                    
						a0_wr[1002]   <= x1002_in;                    
						a0_wr[1003]   <= x1003_in;                    
						a0_wr[1004]   <= x1004_in;                    
						a0_wr[1005]   <= x1005_in;                    
						a0_wr[1006]   <= x1006_in;                    
						a0_wr[1007]   <= x1007_in;                    
						a0_wr[1008]   <= x1008_in;                    
						a0_wr[1009]   <= x1009_in;                    
						a0_wr[1010]   <= x1010_in;                    
						a0_wr[1011]   <= x1011_in;                    
						a0_wr[1012]   <= x1012_in;                    
						a0_wr[1013]   <= x1013_in;                    
						a0_wr[1014]   <= x1014_in;                    
						a0_wr[1015]   <= x1015_in;                    
						a0_wr[1016]   <= x1016_in;                    
						a0_wr[1017]   <= x1017_in;                    
						a0_wr[1018]   <= x1018_in;                    
						a0_wr[1019]   <= x1019_in;                    
						a0_wr[1020]   <= x1020_in;                    
						a0_wr[1021]   <= x1021_in;                    
						a0_wr[1022]   <= x1022_in;                    
						a0_wr[1023]   <= x1023_in;                    
						a0_wr[1024]   <= x1024_in;                    
						a0_wr[1025]   <= x1025_in;                    
						a0_wr[1026]   <= x1026_in;                    
						a0_wr[1027]   <= x1027_in;                    
						a0_wr[1028]   <= x1028_in;                    
						a0_wr[1029]   <= x1029_in;                    
						a0_wr[1030]   <= x1030_in;                    
						a0_wr[1031]   <= x1031_in;                    
						a0_wr[1032]   <= x1032_in;                    
						a0_wr[1033]   <= x1033_in;                    
						a0_wr[1034]   <= x1034_in;                    
						a0_wr[1035]   <= x1035_in;                    
						a0_wr[1036]   <= x1036_in;                    
						a0_wr[1037]   <= x1037_in;                    
						a0_wr[1038]   <= x1038_in;                    
						a0_wr[1039]   <= x1039_in;                    
						a0_wr[1040]   <= x1040_in;                    
						a0_wr[1041]   <= x1041_in;                    
						a0_wr[1042]   <= x1042_in;                    
						a0_wr[1043]   <= x1043_in;                    
						a0_wr[1044]   <= x1044_in;                    
						a0_wr[1045]   <= x1045_in;                    
						a0_wr[1046]   <= x1046_in;                    
						a0_wr[1047]   <= x1047_in;                    
						a0_wr[1048]   <= x1048_in;                    
						a0_wr[1049]   <= x1049_in;                    
						a0_wr[1050]   <= x1050_in;                    
						a0_wr[1051]   <= x1051_in;                    
						a0_wr[1052]   <= x1052_in;                    
						a0_wr[1053]   <= x1053_in;                    
						a0_wr[1054]   <= x1054_in;                    
						a0_wr[1055]   <= x1055_in;                    
						a0_wr[1056]   <= x1056_in;                    
						a0_wr[1057]   <= x1057_in;                    
						a0_wr[1058]   <= x1058_in;                    
						a0_wr[1059]   <= x1059_in;                    
						a0_wr[1060]   <= x1060_in;                    
						a0_wr[1061]   <= x1061_in;                    
						a0_wr[1062]   <= x1062_in;                    
						a0_wr[1063]   <= x1063_in;                    
						a0_wr[1064]   <= x1064_in;                    
						a0_wr[1065]   <= x1065_in;                    
						a0_wr[1066]   <= x1066_in;                    
						a0_wr[1067]   <= x1067_in;                    
						a0_wr[1068]   <= x1068_in;                    
						a0_wr[1069]   <= x1069_in;                    
						a0_wr[1070]   <= x1070_in;                    
						a0_wr[1071]   <= x1071_in;                    
						a0_wr[1072]   <= x1072_in;                    
						a0_wr[1073]   <= x1073_in;                    
						a0_wr[1074]   <= x1074_in;                    
						a0_wr[1075]   <= x1075_in;                    
						a0_wr[1076]   <= x1076_in;                    
						a0_wr[1077]   <= x1077_in;                    
						a0_wr[1078]   <= x1078_in;                    
						a0_wr[1079]   <= x1079_in;                    
						a0_wr[1080]   <= x1080_in;                    
						a0_wr[1081]   <= x1081_in;                    
						a0_wr[1082]   <= x1082_in;                    
						a0_wr[1083]   <= x1083_in;                    
						a0_wr[1084]   <= x1084_in;                    
						a0_wr[1085]   <= x1085_in;                    
						a0_wr[1086]   <= x1086_in;                    
						a0_wr[1087]   <= x1087_in;                    
						a0_wr[1088]   <= x1088_in;                    
						a0_wr[1089]   <= x1089_in;                    
						a0_wr[1090]   <= x1090_in;                    
						a0_wr[1091]   <= x1091_in;                    
						a0_wr[1092]   <= x1092_in;                    
						a0_wr[1093]   <= x1093_in;                    
						a0_wr[1094]   <= x1094_in;                    
						a0_wr[1095]   <= x1095_in;                    
						a0_wr[1096]   <= x1096_in;                    
						a0_wr[1097]   <= x1097_in;                    
						a0_wr[1098]   <= x1098_in;                    
						a0_wr[1099]   <= x1099_in;                    
						a0_wr[1100]   <= x1100_in;                    
						a0_wr[1101]   <= x1101_in;                    
						a0_wr[1102]   <= x1102_in;                    
						a0_wr[1103]   <= x1103_in;                    
						a0_wr[1104]   <= x1104_in;                    
						a0_wr[1105]   <= x1105_in;                    
						a0_wr[1106]   <= x1106_in;                    
						a0_wr[1107]   <= x1107_in;                    
						a0_wr[1108]   <= x1108_in;                    
						a0_wr[1109]   <= x1109_in;                    
						a0_wr[1110]   <= x1110_in;                    
						a0_wr[1111]   <= x1111_in;                    
						a0_wr[1112]   <= x1112_in;                    
						a0_wr[1113]   <= x1113_in;                    
						a0_wr[1114]   <= x1114_in;                    
						a0_wr[1115]   <= x1115_in;                    
						a0_wr[1116]   <= x1116_in;                    
						a0_wr[1117]   <= x1117_in;                    
						a0_wr[1118]   <= x1118_in;                    
						a0_wr[1119]   <= x1119_in;                    
						a0_wr[1120]   <= x1120_in;                    
						a0_wr[1121]   <= x1121_in;                    
						a0_wr[1122]   <= x1122_in;                    
						a0_wr[1123]   <= x1123_in;                    
						a0_wr[1124]   <= x1124_in;                    
						a0_wr[1125]   <= x1125_in;                    
						a0_wr[1126]   <= x1126_in;                    
						a0_wr[1127]   <= x1127_in;                    
						a0_wr[1128]   <= x1128_in;                    
						a0_wr[1129]   <= x1129_in;                    
						a0_wr[1130]   <= x1130_in;                    
						a0_wr[1131]   <= x1131_in;                    
						a0_wr[1132]   <= x1132_in;                    
						a0_wr[1133]   <= x1133_in;                    
						a0_wr[1134]   <= x1134_in;                    
						a0_wr[1135]   <= x1135_in;                    
						a0_wr[1136]   <= x1136_in;                    
						a0_wr[1137]   <= x1137_in;                    
						a0_wr[1138]   <= x1138_in;                    
						a0_wr[1139]   <= x1139_in;                    
						a0_wr[1140]   <= x1140_in;                    
						a0_wr[1141]   <= x1141_in;                    
						a0_wr[1142]   <= x1142_in;                    
						a0_wr[1143]   <= x1143_in;                    
						a0_wr[1144]   <= x1144_in;                    
						a0_wr[1145]   <= x1145_in;                    
						a0_wr[1146]   <= x1146_in;                    
						a0_wr[1147]   <= x1147_in;                    
						a0_wr[1148]   <= x1148_in;                    
						a0_wr[1149]   <= x1149_in;                    
						a0_wr[1150]   <= x1150_in;                    
						a0_wr[1151]   <= x1151_in;                    
						a0_wr[1152]   <= x1152_in;                    
						a0_wr[1153]   <= x1153_in;                    
						a0_wr[1154]   <= x1154_in;                    
						a0_wr[1155]   <= x1155_in;                    
						a0_wr[1156]   <= x1156_in;                    
						a0_wr[1157]   <= x1157_in;                    
						a0_wr[1158]   <= x1158_in;                    
						a0_wr[1159]   <= x1159_in;                    
						a0_wr[1160]   <= x1160_in;                    
						a0_wr[1161]   <= x1161_in;                    
						a0_wr[1162]   <= x1162_in;                    
						a0_wr[1163]   <= x1163_in;                    
						a0_wr[1164]   <= x1164_in;                    
						a0_wr[1165]   <= x1165_in;                    
						a0_wr[1166]   <= x1166_in;                    
						a0_wr[1167]   <= x1167_in;                    
						a0_wr[1168]   <= x1168_in;                    
						a0_wr[1169]   <= x1169_in;                    
						a0_wr[1170]   <= x1170_in;                    
						a0_wr[1171]   <= x1171_in;                    
						a0_wr[1172]   <= x1172_in;                    
						a0_wr[1173]   <= x1173_in;                    
						a0_wr[1174]   <= x1174_in;                    
						a0_wr[1175]   <= x1175_in;                    
						a0_wr[1176]   <= x1176_in;                    
						a0_wr[1177]   <= x1177_in;                    
						a0_wr[1178]   <= x1178_in;                    
						a0_wr[1179]   <= x1179_in;                    
						a0_wr[1180]   <= x1180_in;                    
						a0_wr[1181]   <= x1181_in;                    
						a0_wr[1182]   <= x1182_in;                    
						a0_wr[1183]   <= x1183_in;                    
						a0_wr[1184]   <= x1184_in;                    
						a0_wr[1185]   <= x1185_in;                    
						a0_wr[1186]   <= x1186_in;                    
						a0_wr[1187]   <= x1187_in;                    
						a0_wr[1188]   <= x1188_in;                    
						a0_wr[1189]   <= x1189_in;                    
						a0_wr[1190]   <= x1190_in;                    
						a0_wr[1191]   <= x1191_in;                    
						a0_wr[1192]   <= x1192_in;                    
						a0_wr[1193]   <= x1193_in;                    
						a0_wr[1194]   <= x1194_in;                    
						a0_wr[1195]   <= x1195_in;                    
						a0_wr[1196]   <= x1196_in;                    
						a0_wr[1197]   <= x1197_in;                    
						a0_wr[1198]   <= x1198_in;                    
						a0_wr[1199]   <= x1199_in;                    
						a0_wr[1200]   <= x1200_in;                    
						a0_wr[1201]   <= x1201_in;                    
						a0_wr[1202]   <= x1202_in;                    
						a0_wr[1203]   <= x1203_in;                    
						a0_wr[1204]   <= x1204_in;                    
						a0_wr[1205]   <= x1205_in;                    
						a0_wr[1206]   <= x1206_in;                    
						a0_wr[1207]   <= x1207_in;                    
						a0_wr[1208]   <= x1208_in;                    
						a0_wr[1209]   <= x1209_in;                    
						a0_wr[1210]   <= x1210_in;                    
						a0_wr[1211]   <= x1211_in;                    
						a0_wr[1212]   <= x1212_in;                    
						a0_wr[1213]   <= x1213_in;                    
						a0_wr[1214]   <= x1214_in;                    
						a0_wr[1215]   <= x1215_in;                    
						a0_wr[1216]   <= x1216_in;                    
						a0_wr[1217]   <= x1217_in;                    
						a0_wr[1218]   <= x1218_in;                    
						a0_wr[1219]   <= x1219_in;                    
						a0_wr[1220]   <= x1220_in;                    
						a0_wr[1221]   <= x1221_in;                    
						a0_wr[1222]   <= x1222_in;                    
						a0_wr[1223]   <= x1223_in;                    
						a0_wr[1224]   <= x1224_in;                    
						a0_wr[1225]   <= x1225_in;                    
						a0_wr[1226]   <= x1226_in;                    
						a0_wr[1227]   <= x1227_in;                    
						a0_wr[1228]   <= x1228_in;                    
						a0_wr[1229]   <= x1229_in;                    
						a0_wr[1230]   <= x1230_in;                    
						a0_wr[1231]   <= x1231_in;                    
						a0_wr[1232]   <= x1232_in;                    
						a0_wr[1233]   <= x1233_in;                    
						a0_wr[1234]   <= x1234_in;                    
						a0_wr[1235]   <= x1235_in;                    
						a0_wr[1236]   <= x1236_in;                    
						a0_wr[1237]   <= x1237_in;                    
						a0_wr[1238]   <= x1238_in;                    
						a0_wr[1239]   <= x1239_in;                    
						a0_wr[1240]   <= x1240_in;                    
						a0_wr[1241]   <= x1241_in;                    
						a0_wr[1242]   <= x1242_in;                    
						a0_wr[1243]   <= x1243_in;                    
						a0_wr[1244]   <= x1244_in;                    
						a0_wr[1245]   <= x1245_in;                    
						a0_wr[1246]   <= x1246_in;                    
						a0_wr[1247]   <= x1247_in;                    
						a0_wr[1248]   <= x1248_in;                    
						a0_wr[1249]   <= x1249_in;                    
						a0_wr[1250]   <= x1250_in;                    
						a0_wr[1251]   <= x1251_in;                    
						a0_wr[1252]   <= x1252_in;                    
						a0_wr[1253]   <= x1253_in;                    
						a0_wr[1254]   <= x1254_in;                    
						a0_wr[1255]   <= x1255_in;                    
						a0_wr[1256]   <= x1256_in;                    
						a0_wr[1257]   <= x1257_in;                    
						a0_wr[1258]   <= x1258_in;                    
						a0_wr[1259]   <= x1259_in;                    
						a0_wr[1260]   <= x1260_in;                    
						a0_wr[1261]   <= x1261_in;                    
						a0_wr[1262]   <= x1262_in;                    
						a0_wr[1263]   <= x1263_in;                    
						a0_wr[1264]   <= x1264_in;                    
						a0_wr[1265]   <= x1265_in;                    
						a0_wr[1266]   <= x1266_in;                    
						a0_wr[1267]   <= x1267_in;                    
						a0_wr[1268]   <= x1268_in;                    
						a0_wr[1269]   <= x1269_in;                    
						a0_wr[1270]   <= x1270_in;                    
						a0_wr[1271]   <= x1271_in;                    
						a0_wr[1272]   <= x1272_in;                    
						a0_wr[1273]   <= x1273_in;                    
						a0_wr[1274]   <= x1274_in;                    
						a0_wr[1275]   <= x1275_in;                    
						a0_wr[1276]   <= x1276_in;                    
						a0_wr[1277]   <= x1277_in;                    
						a0_wr[1278]   <= x1278_in;                    
						a0_wr[1279]   <= x1279_in;                    
						a0_wr[1280]   <= x1280_in;                    
						a0_wr[1281]   <= x1281_in;                    
						a0_wr[1282]   <= x1282_in;                    
						a0_wr[1283]   <= x1283_in;                    
						a0_wr[1284]   <= x1284_in;                    
						a0_wr[1285]   <= x1285_in;                    
						a0_wr[1286]   <= x1286_in;                    
						a0_wr[1287]   <= x1287_in;                    
						a0_wr[1288]   <= x1288_in;                    
						a0_wr[1289]   <= x1289_in;                    
						a0_wr[1290]   <= x1290_in;                    
						a0_wr[1291]   <= x1291_in;                    
						a0_wr[1292]   <= x1292_in;                    
						a0_wr[1293]   <= x1293_in;                    
						a0_wr[1294]   <= x1294_in;                    
						a0_wr[1295]   <= x1295_in;                    
						a0_wr[1296]   <= x1296_in;                    
						a0_wr[1297]   <= x1297_in;                    
						a0_wr[1298]   <= x1298_in;                    
						a0_wr[1299]   <= x1299_in;                    
						a0_wr[1300]   <= x1300_in;                    
						a0_wr[1301]   <= x1301_in;                    
						a0_wr[1302]   <= x1302_in;                    
						a0_wr[1303]   <= x1303_in;                    
						a0_wr[1304]   <= x1304_in;                    
						a0_wr[1305]   <= x1305_in;                    
						a0_wr[1306]   <= x1306_in;                    
						a0_wr[1307]   <= x1307_in;                    
						a0_wr[1308]   <= x1308_in;                    
						a0_wr[1309]   <= x1309_in;                    
						a0_wr[1310]   <= x1310_in;                    
						a0_wr[1311]   <= x1311_in;                    
						a0_wr[1312]   <= x1312_in;                    
						a0_wr[1313]   <= x1313_in;                    
						a0_wr[1314]   <= x1314_in;                    
						a0_wr[1315]   <= x1315_in;                    
						a0_wr[1316]   <= x1316_in;                    
						a0_wr[1317]   <= x1317_in;                    
						a0_wr[1318]   <= x1318_in;                    
						a0_wr[1319]   <= x1319_in;                    
						a0_wr[1320]   <= x1320_in;                    
						a0_wr[1321]   <= x1321_in;                    
						a0_wr[1322]   <= x1322_in;                    
						a0_wr[1323]   <= x1323_in;                    
						a0_wr[1324]   <= x1324_in;                    
						a0_wr[1325]   <= x1325_in;                    
						a0_wr[1326]   <= x1326_in;                    
						a0_wr[1327]   <= x1327_in;                    
						a0_wr[1328]   <= x1328_in;                    
						a0_wr[1329]   <= x1329_in;                    
						a0_wr[1330]   <= x1330_in;                    
						a0_wr[1331]   <= x1331_in;                    
						a0_wr[1332]   <= x1332_in;                    
						a0_wr[1333]   <= x1333_in;                    
						a0_wr[1334]   <= x1334_in;                    
						a0_wr[1335]   <= x1335_in;                    
						a0_wr[1336]   <= x1336_in;                    
						a0_wr[1337]   <= x1337_in;                    
						a0_wr[1338]   <= x1338_in;                    
						a0_wr[1339]   <= x1339_in;                    
						a0_wr[1340]   <= x1340_in;                    
						a0_wr[1341]   <= x1341_in;                    
						a0_wr[1342]   <= x1342_in;                    
						a0_wr[1343]   <= x1343_in;                    
						a0_wr[1344]   <= x1344_in;                    
						a0_wr[1345]   <= x1345_in;                    
						a0_wr[1346]   <= x1346_in;                    
						a0_wr[1347]   <= x1347_in;                    
						a0_wr[1348]   <= x1348_in;                    
						a0_wr[1349]   <= x1349_in;                    
						a0_wr[1350]   <= x1350_in;                    
						a0_wr[1351]   <= x1351_in;                    
						a0_wr[1352]   <= x1352_in;                    
						a0_wr[1353]   <= x1353_in;                    
						a0_wr[1354]   <= x1354_in;                    
						a0_wr[1355]   <= x1355_in;                    
						a0_wr[1356]   <= x1356_in;                    
						a0_wr[1357]   <= x1357_in;                    
						a0_wr[1358]   <= x1358_in;                    
						a0_wr[1359]   <= x1359_in;                    
						a0_wr[1360]   <= x1360_in;                    
						a0_wr[1361]   <= x1361_in;                    
						a0_wr[1362]   <= x1362_in;                    
						a0_wr[1363]   <= x1363_in;                    
						a0_wr[1364]   <= x1364_in;                    
						a0_wr[1365]   <= x1365_in;                    
						a0_wr[1366]   <= x1366_in;                    
						a0_wr[1367]   <= x1367_in;                    
						a0_wr[1368]   <= x1368_in;                    
						a0_wr[1369]   <= x1369_in;                    
						a0_wr[1370]   <= x1370_in;                    
						a0_wr[1371]   <= x1371_in;                    
						a0_wr[1372]   <= x1372_in;                    
						a0_wr[1373]   <= x1373_in;                    
						a0_wr[1374]   <= x1374_in;                    
						a0_wr[1375]   <= x1375_in;                    
						a0_wr[1376]   <= x1376_in;                    
						a0_wr[1377]   <= x1377_in;                    
						a0_wr[1378]   <= x1378_in;                    
						a0_wr[1379]   <= x1379_in;                    
						a0_wr[1380]   <= x1380_in;                    
						a0_wr[1381]   <= x1381_in;                    
						a0_wr[1382]   <= x1382_in;                    
						a0_wr[1383]   <= x1383_in;                    
						a0_wr[1384]   <= x1384_in;                    
						a0_wr[1385]   <= x1385_in;                    
						a0_wr[1386]   <= x1386_in;                    
						a0_wr[1387]   <= x1387_in;                    
						a0_wr[1388]   <= x1388_in;                    
						a0_wr[1389]   <= x1389_in;                    
						a0_wr[1390]   <= x1390_in;                    
						a0_wr[1391]   <= x1391_in;                    
						a0_wr[1392]   <= x1392_in;                    
						a0_wr[1393]   <= x1393_in;                    
						a0_wr[1394]   <= x1394_in;                    
						a0_wr[1395]   <= x1395_in;                    
						a0_wr[1396]   <= x1396_in;                    
						a0_wr[1397]   <= x1397_in;                    
						a0_wr[1398]   <= x1398_in;                    
						a0_wr[1399]   <= x1399_in;                    
						a0_wr[1400]   <= x1400_in;                    
						a0_wr[1401]   <= x1401_in;                    
						a0_wr[1402]   <= x1402_in;                    
						a0_wr[1403]   <= x1403_in;                    
						a0_wr[1404]   <= x1404_in;                    
						a0_wr[1405]   <= x1405_in;                    
						a0_wr[1406]   <= x1406_in;                    
						a0_wr[1407]   <= x1407_in;                    
						a0_wr[1408]   <= x1408_in;                    
						a0_wr[1409]   <= x1409_in;                    
						a0_wr[1410]   <= x1410_in;                    
						a0_wr[1411]   <= x1411_in;                    
						a0_wr[1412]   <= x1412_in;                    
						a0_wr[1413]   <= x1413_in;                    
						a0_wr[1414]   <= x1414_in;                    
						a0_wr[1415]   <= x1415_in;                    
						a0_wr[1416]   <= x1416_in;                    
						a0_wr[1417]   <= x1417_in;                    
						a0_wr[1418]   <= x1418_in;                    
						a0_wr[1419]   <= x1419_in;                    
						a0_wr[1420]   <= x1420_in;                    
						a0_wr[1421]   <= x1421_in;                    
						a0_wr[1422]   <= x1422_in;                    
						a0_wr[1423]   <= x1423_in;                    
						a0_wr[1424]   <= x1424_in;                    
						a0_wr[1425]   <= x1425_in;                    
						a0_wr[1426]   <= x1426_in;                    
						a0_wr[1427]   <= x1427_in;                    
						a0_wr[1428]   <= x1428_in;                    
						a0_wr[1429]   <= x1429_in;                    
						a0_wr[1430]   <= x1430_in;                    
						a0_wr[1431]   <= x1431_in;                    
						a0_wr[1432]   <= x1432_in;                    
						a0_wr[1433]   <= x1433_in;                    
						a0_wr[1434]   <= x1434_in;                    
						a0_wr[1435]   <= x1435_in;                    
						a0_wr[1436]   <= x1436_in;                    
						a0_wr[1437]   <= x1437_in;                    
						a0_wr[1438]   <= x1438_in;                    
						a0_wr[1439]   <= x1439_in;                    
						a0_wr[1440]   <= x1440_in;                    
						a0_wr[1441]   <= x1441_in;                    
						a0_wr[1442]   <= x1442_in;                    
						a0_wr[1443]   <= x1443_in;                    
						a0_wr[1444]   <= x1444_in;                    
						a0_wr[1445]   <= x1445_in;                    
						a0_wr[1446]   <= x1446_in;                    
						a0_wr[1447]   <= x1447_in;                    
						a0_wr[1448]   <= x1448_in;                    
						a0_wr[1449]   <= x1449_in;                    
						a0_wr[1450]   <= x1450_in;                    
						a0_wr[1451]   <= x1451_in;                    
						a0_wr[1452]   <= x1452_in;                    
						a0_wr[1453]   <= x1453_in;                    
						a0_wr[1454]   <= x1454_in;                    
						a0_wr[1455]   <= x1455_in;                    
						a0_wr[1456]   <= x1456_in;                    
						a0_wr[1457]   <= x1457_in;                    
						a0_wr[1458]   <= x1458_in;                    
						a0_wr[1459]   <= x1459_in;                    
						a0_wr[1460]   <= x1460_in;                    
						a0_wr[1461]   <= x1461_in;                    
						a0_wr[1462]   <= x1462_in;                    
						a0_wr[1463]   <= x1463_in;                    
						a0_wr[1464]   <= x1464_in;                    
						a0_wr[1465]   <= x1465_in;                    
						a0_wr[1466]   <= x1466_in;                    
						a0_wr[1467]   <= x1467_in;                    
						a0_wr[1468]   <= x1468_in;                    
						a0_wr[1469]   <= x1469_in;                    
						a0_wr[1470]   <= x1470_in;                    
						a0_wr[1471]   <= x1471_in;                    
						a0_wr[1472]   <= x1472_in;                    
						a0_wr[1473]   <= x1473_in;                    
						a0_wr[1474]   <= x1474_in;                    
						a0_wr[1475]   <= x1475_in;                    
						a0_wr[1476]   <= x1476_in;                    
						a0_wr[1477]   <= x1477_in;                    
						a0_wr[1478]   <= x1478_in;                    
						a0_wr[1479]   <= x1479_in;                    
						a0_wr[1480]   <= x1480_in;                    
						a0_wr[1481]   <= x1481_in;                    
						a0_wr[1482]   <= x1482_in;                    
						a0_wr[1483]   <= x1483_in;                    
						a0_wr[1484]   <= x1484_in;                    
						a0_wr[1485]   <= x1485_in;                    
						a0_wr[1486]   <= x1486_in;                    
						a0_wr[1487]   <= x1487_in;                    
						a0_wr[1488]   <= x1488_in;                    
						a0_wr[1489]   <= x1489_in;                    
						a0_wr[1490]   <= x1490_in;                    
						a0_wr[1491]   <= x1491_in;                    
						a0_wr[1492]   <= x1492_in;                    
						a0_wr[1493]   <= x1493_in;                    
						a0_wr[1494]   <= x1494_in;                    
						a0_wr[1495]   <= x1495_in;                    
						a0_wr[1496]   <= x1496_in;                    
						a0_wr[1497]   <= x1497_in;                    
						a0_wr[1498]   <= x1498_in;                    
						a0_wr[1499]   <= x1499_in;                    
						a0_wr[1500]   <= x1500_in;                    
						a0_wr[1501]   <= x1501_in;                    
						a0_wr[1502]   <= x1502_in;                    
						a0_wr[1503]   <= x1503_in;                    
						a0_wr[1504]   <= x1504_in;                    
						a0_wr[1505]   <= x1505_in;                    
						a0_wr[1506]   <= x1506_in;                    
						a0_wr[1507]   <= x1507_in;                    
						a0_wr[1508]   <= x1508_in;                    
						a0_wr[1509]   <= x1509_in;                    
						a0_wr[1510]   <= x1510_in;                    
						a0_wr[1511]   <= x1511_in;                    
						a0_wr[1512]   <= x1512_in;                    
						a0_wr[1513]   <= x1513_in;                    
						a0_wr[1514]   <= x1514_in;                    
						a0_wr[1515]   <= x1515_in;                    
						a0_wr[1516]   <= x1516_in;                    
						a0_wr[1517]   <= x1517_in;                    
						a0_wr[1518]   <= x1518_in;                    
						a0_wr[1519]   <= x1519_in;                    
						a0_wr[1520]   <= x1520_in;                    
						a0_wr[1521]   <= x1521_in;                    
						a0_wr[1522]   <= x1522_in;                    
						a0_wr[1523]   <= x1523_in;                    
						a0_wr[1524]   <= x1524_in;                    
						a0_wr[1525]   <= x1525_in;                    
						a0_wr[1526]   <= x1526_in;                    
						a0_wr[1527]   <= x1527_in;                    
						a0_wr[1528]   <= x1528_in;                    
						a0_wr[1529]   <= x1529_in;                    
						a0_wr[1530]   <= x1530_in;                    
						a0_wr[1531]   <= x1531_in;                    
						a0_wr[1532]   <= x1532_in;                    
						a0_wr[1533]   <= x1533_in;                    
						a0_wr[1534]   <= x1534_in;                    
						a0_wr[1535]   <= x1535_in;                    
						a0_wr[1536]   <= x1536_in;                    
						a0_wr[1537]   <= x1537_in;                    
						a0_wr[1538]   <= x1538_in;                    
						a0_wr[1539]   <= x1539_in;                    
						a0_wr[1540]   <= x1540_in;                    
						a0_wr[1541]   <= x1541_in;                    
						a0_wr[1542]   <= x1542_in;                    
						a0_wr[1543]   <= x1543_in;                    
						a0_wr[1544]   <= x1544_in;                    
						a0_wr[1545]   <= x1545_in;                    
						a0_wr[1546]   <= x1546_in;                    
						a0_wr[1547]   <= x1547_in;                    
						a0_wr[1548]   <= x1548_in;                    
						a0_wr[1549]   <= x1549_in;                    
						a0_wr[1550]   <= x1550_in;                    
						a0_wr[1551]   <= x1551_in;                    
						a0_wr[1552]   <= x1552_in;                    
						a0_wr[1553]   <= x1553_in;                    
						a0_wr[1554]   <= x1554_in;                    
						a0_wr[1555]   <= x1555_in;                    
						a0_wr[1556]   <= x1556_in;                    
						a0_wr[1557]   <= x1557_in;                    
						a0_wr[1558]   <= x1558_in;                    
						a0_wr[1559]   <= x1559_in;                    
						a0_wr[1560]   <= x1560_in;                    
						a0_wr[1561]   <= x1561_in;                    
						a0_wr[1562]   <= x1562_in;                    
						a0_wr[1563]   <= x1563_in;                    
						a0_wr[1564]   <= x1564_in;                    
						a0_wr[1565]   <= x1565_in;                    
						a0_wr[1566]   <= x1566_in;                    
						a0_wr[1567]   <= x1567_in;                    
						a0_wr[1568]   <= x1568_in;                    
						a0_wr[1569]   <= x1569_in;                    
						a0_wr[1570]   <= x1570_in;                    
						a0_wr[1571]   <= x1571_in;                    
						a0_wr[1572]   <= x1572_in;                    
						a0_wr[1573]   <= x1573_in;                    
						a0_wr[1574]   <= x1574_in;                    
						a0_wr[1575]   <= x1575_in;                    
						a0_wr[1576]   <= x1576_in;                    
						a0_wr[1577]   <= x1577_in;                    
						a0_wr[1578]   <= x1578_in;                    
						a0_wr[1579]   <= x1579_in;                    
						a0_wr[1580]   <= x1580_in;                    
						a0_wr[1581]   <= x1581_in;                    
						a0_wr[1582]   <= x1582_in;                    
						a0_wr[1583]   <= x1583_in;                    
						a0_wr[1584]   <= x1584_in;                    
						a0_wr[1585]   <= x1585_in;                    
						a0_wr[1586]   <= x1586_in;                    
						a0_wr[1587]   <= x1587_in;                    
						a0_wr[1588]   <= x1588_in;                    
						a0_wr[1589]   <= x1589_in;                    
						a0_wr[1590]   <= x1590_in;                    
						a0_wr[1591]   <= x1591_in;                    
						a0_wr[1592]   <= x1592_in;                    
						a0_wr[1593]   <= x1593_in;                    
						a0_wr[1594]   <= x1594_in;                    
						a0_wr[1595]   <= x1595_in;                    
						a0_wr[1596]   <= x1596_in;                    
						a0_wr[1597]   <= x1597_in;                    
						a0_wr[1598]   <= x1598_in;                    
						a0_wr[1599]   <= x1599_in;                    
						a0_wr[1600]   <= x1600_in;                    
						a0_wr[1601]   <= x1601_in;                    
						a0_wr[1602]   <= x1602_in;                    
						a0_wr[1603]   <= x1603_in;                    
						a0_wr[1604]   <= x1604_in;                    
						a0_wr[1605]   <= x1605_in;                    
						a0_wr[1606]   <= x1606_in;                    
						a0_wr[1607]   <= x1607_in;                    
						a0_wr[1608]   <= x1608_in;                    
						a0_wr[1609]   <= x1609_in;                    
						a0_wr[1610]   <= x1610_in;                    
						a0_wr[1611]   <= x1611_in;                    
						a0_wr[1612]   <= x1612_in;                    
						a0_wr[1613]   <= x1613_in;                    
						a0_wr[1614]   <= x1614_in;                    
						a0_wr[1615]   <= x1615_in;                    
						a0_wr[1616]   <= x1616_in;                    
						a0_wr[1617]   <= x1617_in;                    
						a0_wr[1618]   <= x1618_in;                    
						a0_wr[1619]   <= x1619_in;                    
						a0_wr[1620]   <= x1620_in;                    
						a0_wr[1621]   <= x1621_in;                    
						a0_wr[1622]   <= x1622_in;                    
						a0_wr[1623]   <= x1623_in;                    
						a0_wr[1624]   <= x1624_in;                    
						a0_wr[1625]   <= x1625_in;                    
						a0_wr[1626]   <= x1626_in;                    
						a0_wr[1627]   <= x1627_in;                    
						a0_wr[1628]   <= x1628_in;                    
						a0_wr[1629]   <= x1629_in;                    
						a0_wr[1630]   <= x1630_in;                    
						a0_wr[1631]   <= x1631_in;                    
						a0_wr[1632]   <= x1632_in;                    
						a0_wr[1633]   <= x1633_in;                    
						a0_wr[1634]   <= x1634_in;                    
						a0_wr[1635]   <= x1635_in;                    
						a0_wr[1636]   <= x1636_in;                    
						a0_wr[1637]   <= x1637_in;                    
						a0_wr[1638]   <= x1638_in;                    
						a0_wr[1639]   <= x1639_in;                    
						a0_wr[1640]   <= x1640_in;                    
						a0_wr[1641]   <= x1641_in;                    
						a0_wr[1642]   <= x1642_in;                    
						a0_wr[1643]   <= x1643_in;                    
						a0_wr[1644]   <= x1644_in;                    
						a0_wr[1645]   <= x1645_in;                    
						a0_wr[1646]   <= x1646_in;                    
						a0_wr[1647]   <= x1647_in;                    
						a0_wr[1648]   <= x1648_in;                    
						a0_wr[1649]   <= x1649_in;                    
						a0_wr[1650]   <= x1650_in;                    
						a0_wr[1651]   <= x1651_in;                    
						a0_wr[1652]   <= x1652_in;                    
						a0_wr[1653]   <= x1653_in;                    
						a0_wr[1654]   <= x1654_in;                    
						a0_wr[1655]   <= x1655_in;                    
						a0_wr[1656]   <= x1656_in;                    
						a0_wr[1657]   <= x1657_in;                    
						a0_wr[1658]   <= x1658_in;                    
						a0_wr[1659]   <= x1659_in;                    
						a0_wr[1660]   <= x1660_in;                    
						a0_wr[1661]   <= x1661_in;                    
						a0_wr[1662]   <= x1662_in;                    
						a0_wr[1663]   <= x1663_in;                    
						a0_wr[1664]   <= x1664_in;                    
						a0_wr[1665]   <= x1665_in;                    
						a0_wr[1666]   <= x1666_in;                    
						a0_wr[1667]   <= x1667_in;                    
						a0_wr[1668]   <= x1668_in;                    
						a0_wr[1669]   <= x1669_in;                    
						a0_wr[1670]   <= x1670_in;                    
						a0_wr[1671]   <= x1671_in;                    
						a0_wr[1672]   <= x1672_in;                    
						a0_wr[1673]   <= x1673_in;                    
						a0_wr[1674]   <= x1674_in;                    
						a0_wr[1675]   <= x1675_in;                    
						a0_wr[1676]   <= x1676_in;                    
						a0_wr[1677]   <= x1677_in;                    
						a0_wr[1678]   <= x1678_in;                    
						a0_wr[1679]   <= x1679_in;                    
						a0_wr[1680]   <= x1680_in;                    
						a0_wr[1681]   <= x1681_in;                    
						a0_wr[1682]   <= x1682_in;                    
						a0_wr[1683]   <= x1683_in;                    
						a0_wr[1684]   <= x1684_in;                    
						a0_wr[1685]   <= x1685_in;                    
						a0_wr[1686]   <= x1686_in;                    
						a0_wr[1687]   <= x1687_in;                    
						a0_wr[1688]   <= x1688_in;                    
						a0_wr[1689]   <= x1689_in;                    
						a0_wr[1690]   <= x1690_in;                    
						a0_wr[1691]   <= x1691_in;                    
						a0_wr[1692]   <= x1692_in;                    
						a0_wr[1693]   <= x1693_in;                    
						a0_wr[1694]   <= x1694_in;                    
						a0_wr[1695]   <= x1695_in;                    
						a0_wr[1696]   <= x1696_in;                    
						a0_wr[1697]   <= x1697_in;                    
						a0_wr[1698]   <= x1698_in;                    
						a0_wr[1699]   <= x1699_in;                    
						a0_wr[1700]   <= x1700_in;                    
						a0_wr[1701]   <= x1701_in;                    
						a0_wr[1702]   <= x1702_in;                    
						a0_wr[1703]   <= x1703_in;                    
						a0_wr[1704]   <= x1704_in;                    
						a0_wr[1705]   <= x1705_in;                    
						a0_wr[1706]   <= x1706_in;                    
						a0_wr[1707]   <= x1707_in;                    
						a0_wr[1708]   <= x1708_in;                    
						a0_wr[1709]   <= x1709_in;                    
						a0_wr[1710]   <= x1710_in;                    
						a0_wr[1711]   <= x1711_in;                    
						a0_wr[1712]   <= x1712_in;                    
						a0_wr[1713]   <= x1713_in;                    
						a0_wr[1714]   <= x1714_in;                    
						a0_wr[1715]   <= x1715_in;                    
						a0_wr[1716]   <= x1716_in;                    
						a0_wr[1717]   <= x1717_in;                    
						a0_wr[1718]   <= x1718_in;                    
						a0_wr[1719]   <= x1719_in;                    
						a0_wr[1720]   <= x1720_in;                    
						a0_wr[1721]   <= x1721_in;                    
						a0_wr[1722]   <= x1722_in;                    
						a0_wr[1723]   <= x1723_in;                    
						a0_wr[1724]   <= x1724_in;                    
						a0_wr[1725]   <= x1725_in;                    
						a0_wr[1726]   <= x1726_in;                    
						a0_wr[1727]   <= x1727_in;                    
						a0_wr[1728]   <= x1728_in;                    
						a0_wr[1729]   <= x1729_in;                    
						a0_wr[1730]   <= x1730_in;                    
						a0_wr[1731]   <= x1731_in;                    
						a0_wr[1732]   <= x1732_in;                    
						a0_wr[1733]   <= x1733_in;                    
						a0_wr[1734]   <= x1734_in;                    
						a0_wr[1735]   <= x1735_in;                    
						a0_wr[1736]   <= x1736_in;                    
						a0_wr[1737]   <= x1737_in;                    
						a0_wr[1738]   <= x1738_in;                    
						a0_wr[1739]   <= x1739_in;                    
						a0_wr[1740]   <= x1740_in;                    
						a0_wr[1741]   <= x1741_in;                    
						a0_wr[1742]   <= x1742_in;                    
						a0_wr[1743]   <= x1743_in;                    
						a0_wr[1744]   <= x1744_in;                    
						a0_wr[1745]   <= x1745_in;                    
						a0_wr[1746]   <= x1746_in;                    
						a0_wr[1747]   <= x1747_in;                    
						a0_wr[1748]   <= x1748_in;                    
						a0_wr[1749]   <= x1749_in;                    
						a0_wr[1750]   <= x1750_in;                    
						a0_wr[1751]   <= x1751_in;                    
						a0_wr[1752]   <= x1752_in;                    
						a0_wr[1753]   <= x1753_in;                    
						a0_wr[1754]   <= x1754_in;                    
						a0_wr[1755]   <= x1755_in;                    
						a0_wr[1756]   <= x1756_in;                    
						a0_wr[1757]   <= x1757_in;                    
						a0_wr[1758]   <= x1758_in;                    
						a0_wr[1759]   <= x1759_in;                    
						a0_wr[1760]   <= x1760_in;                    
						a0_wr[1761]   <= x1761_in;                    
						a0_wr[1762]   <= x1762_in;                    
						a0_wr[1763]   <= x1763_in;                    
						a0_wr[1764]   <= x1764_in;                    
						a0_wr[1765]   <= x1765_in;                    
						a0_wr[1766]   <= x1766_in;                    
						a0_wr[1767]   <= x1767_in;                    
						a0_wr[1768]   <= x1768_in;                    
						a0_wr[1769]   <= x1769_in;                    
						a0_wr[1770]   <= x1770_in;                    
						a0_wr[1771]   <= x1771_in;                    
						a0_wr[1772]   <= x1772_in;                    
						a0_wr[1773]   <= x1773_in;                    
						a0_wr[1774]   <= x1774_in;                    
						a0_wr[1775]   <= x1775_in;                    
						a0_wr[1776]   <= x1776_in;                    
						a0_wr[1777]   <= x1777_in;                    
						a0_wr[1778]   <= x1778_in;                    
						a0_wr[1779]   <= x1779_in;                    
						a0_wr[1780]   <= x1780_in;                    
						a0_wr[1781]   <= x1781_in;                    
						a0_wr[1782]   <= x1782_in;                    
						a0_wr[1783]   <= x1783_in;                    
						a0_wr[1784]   <= x1784_in;                    
						a0_wr[1785]   <= x1785_in;                    
						a0_wr[1786]   <= x1786_in;                    
						a0_wr[1787]   <= x1787_in;                    
						a0_wr[1788]   <= x1788_in;                    
						a0_wr[1789]   <= x1789_in;                    
						a0_wr[1790]   <= x1790_in;                    
						a0_wr[1791]   <= x1791_in;                    
						a0_wr[1792]   <= x1792_in;                    
						a0_wr[1793]   <= x1793_in;                    
						a0_wr[1794]   <= x1794_in;                    
						a0_wr[1795]   <= x1795_in;                    
						a0_wr[1796]   <= x1796_in;                    
						a0_wr[1797]   <= x1797_in;                    
						a0_wr[1798]   <= x1798_in;                    
						a0_wr[1799]   <= x1799_in;                    
						a0_wr[1800]   <= x1800_in;                    
						a0_wr[1801]   <= x1801_in;                    
						a0_wr[1802]   <= x1802_in;                    
						a0_wr[1803]   <= x1803_in;                    
						a0_wr[1804]   <= x1804_in;                    
						a0_wr[1805]   <= x1805_in;                    
						a0_wr[1806]   <= x1806_in;                    
						a0_wr[1807]   <= x1807_in;                    
						a0_wr[1808]   <= x1808_in;                    
						a0_wr[1809]   <= x1809_in;                    
						a0_wr[1810]   <= x1810_in;                    
						a0_wr[1811]   <= x1811_in;                    
						a0_wr[1812]   <= x1812_in;                    
						a0_wr[1813]   <= x1813_in;                    
						a0_wr[1814]   <= x1814_in;                    
						a0_wr[1815]   <= x1815_in;                    
						a0_wr[1816]   <= x1816_in;                    
						a0_wr[1817]   <= x1817_in;                    
						a0_wr[1818]   <= x1818_in;                    
						a0_wr[1819]   <= x1819_in;                    
						a0_wr[1820]   <= x1820_in;                    
						a0_wr[1821]   <= x1821_in;                    
						a0_wr[1822]   <= x1822_in;                    
						a0_wr[1823]   <= x1823_in;                    
						a0_wr[1824]   <= x1824_in;                    
						a0_wr[1825]   <= x1825_in;                    
						a0_wr[1826]   <= x1826_in;                    
						a0_wr[1827]   <= x1827_in;                    
						a0_wr[1828]   <= x1828_in;                    
						a0_wr[1829]   <= x1829_in;                    
						a0_wr[1830]   <= x1830_in;                    
						a0_wr[1831]   <= x1831_in;                    
						a0_wr[1832]   <= x1832_in;                    
						a0_wr[1833]   <= x1833_in;                    
						a0_wr[1834]   <= x1834_in;                    
						a0_wr[1835]   <= x1835_in;                    
						a0_wr[1836]   <= x1836_in;                    
						a0_wr[1837]   <= x1837_in;                    
						a0_wr[1838]   <= x1838_in;                    
						a0_wr[1839]   <= x1839_in;                    
						a0_wr[1840]   <= x1840_in;                    
						a0_wr[1841]   <= x1841_in;                    
						a0_wr[1842]   <= x1842_in;                    
						a0_wr[1843]   <= x1843_in;                    
						a0_wr[1844]   <= x1844_in;                    
						a0_wr[1845]   <= x1845_in;                    
						a0_wr[1846]   <= x1846_in;                    
						a0_wr[1847]   <= x1847_in;                    
						a0_wr[1848]   <= x1848_in;                    
						a0_wr[1849]   <= x1849_in;                    
						a0_wr[1850]   <= x1850_in;                    
						a0_wr[1851]   <= x1851_in;                    
						a0_wr[1852]   <= x1852_in;                    
						a0_wr[1853]   <= x1853_in;                    
						a0_wr[1854]   <= x1854_in;                    
						a0_wr[1855]   <= x1855_in;                    
						a0_wr[1856]   <= x1856_in;                    
						a0_wr[1857]   <= x1857_in;                    
						a0_wr[1858]   <= x1858_in;                    
						a0_wr[1859]   <= x1859_in;                    
						a0_wr[1860]   <= x1860_in;                    
						a0_wr[1861]   <= x1861_in;                    
						a0_wr[1862]   <= x1862_in;                    
						a0_wr[1863]   <= x1863_in;                    
						a0_wr[1864]   <= x1864_in;                    
						a0_wr[1865]   <= x1865_in;                    
						a0_wr[1866]   <= x1866_in;                    
						a0_wr[1867]   <= x1867_in;                    
						a0_wr[1868]   <= x1868_in;                    
						a0_wr[1869]   <= x1869_in;                    
						a0_wr[1870]   <= x1870_in;                    
						a0_wr[1871]   <= x1871_in;                    
						a0_wr[1872]   <= x1872_in;                    
						a0_wr[1873]   <= x1873_in;                    
						a0_wr[1874]   <= x1874_in;                    
						a0_wr[1875]   <= x1875_in;                    
						a0_wr[1876]   <= x1876_in;                    
						a0_wr[1877]   <= x1877_in;                    
						a0_wr[1878]   <= x1878_in;                    
						a0_wr[1879]   <= x1879_in;                    
						a0_wr[1880]   <= x1880_in;                    
						a0_wr[1881]   <= x1881_in;                    
						a0_wr[1882]   <= x1882_in;                    
						a0_wr[1883]   <= x1883_in;                    
						a0_wr[1884]   <= x1884_in;                    
						a0_wr[1885]   <= x1885_in;                    
						a0_wr[1886]   <= x1886_in;                    
						a0_wr[1887]   <= x1887_in;                    
						a0_wr[1888]   <= x1888_in;                    
						a0_wr[1889]   <= x1889_in;                    
						a0_wr[1890]   <= x1890_in;                    
						a0_wr[1891]   <= x1891_in;                    
						a0_wr[1892]   <= x1892_in;                    
						a0_wr[1893]   <= x1893_in;                    
						a0_wr[1894]   <= x1894_in;                    
						a0_wr[1895]   <= x1895_in;                    
						a0_wr[1896]   <= x1896_in;                    
						a0_wr[1897]   <= x1897_in;                    
						a0_wr[1898]   <= x1898_in;                    
						a0_wr[1899]   <= x1899_in;                    
						a0_wr[1900]   <= x1900_in;                    
						a0_wr[1901]   <= x1901_in;                    
						a0_wr[1902]   <= x1902_in;                    
						a0_wr[1903]   <= x1903_in;                    
						a0_wr[1904]   <= x1904_in;                    
						a0_wr[1905]   <= x1905_in;                    
						a0_wr[1906]   <= x1906_in;                    
						a0_wr[1907]   <= x1907_in;                    
						a0_wr[1908]   <= x1908_in;                    
						a0_wr[1909]   <= x1909_in;                    
						a0_wr[1910]   <= x1910_in;                    
						a0_wr[1911]   <= x1911_in;                    
						a0_wr[1912]   <= x1912_in;                    
						a0_wr[1913]   <= x1913_in;                    
						a0_wr[1914]   <= x1914_in;                    
						a0_wr[1915]   <= x1915_in;                    
						a0_wr[1916]   <= x1916_in;                    
						a0_wr[1917]   <= x1917_in;                    
						a0_wr[1918]   <= x1918_in;                    
						a0_wr[1919]   <= x1919_in;                    
						a0_wr[1920]   <= x1920_in;                    
						a0_wr[1921]   <= x1921_in;                    
						a0_wr[1922]   <= x1922_in;                    
						a0_wr[1923]   <= x1923_in;                    
						a0_wr[1924]   <= x1924_in;                    
						a0_wr[1925]   <= x1925_in;                    
						a0_wr[1926]   <= x1926_in;                    
						a0_wr[1927]   <= x1927_in;                    
						a0_wr[1928]   <= x1928_in;                    
						a0_wr[1929]   <= x1929_in;                    
						a0_wr[1930]   <= x1930_in;                    
						a0_wr[1931]   <= x1931_in;                    
						a0_wr[1932]   <= x1932_in;                    
						a0_wr[1933]   <= x1933_in;                    
						a0_wr[1934]   <= x1934_in;                    
						a0_wr[1935]   <= x1935_in;                    
						a0_wr[1936]   <= x1936_in;                    
						a0_wr[1937]   <= x1937_in;                    
						a0_wr[1938]   <= x1938_in;                    
						a0_wr[1939]   <= x1939_in;                    
						a0_wr[1940]   <= x1940_in;                    
						a0_wr[1941]   <= x1941_in;                    
						a0_wr[1942]   <= x1942_in;                    
						a0_wr[1943]   <= x1943_in;                    
						a0_wr[1944]   <= x1944_in;                    
						a0_wr[1945]   <= x1945_in;                    
						a0_wr[1946]   <= x1946_in;                    
						a0_wr[1947]   <= x1947_in;                    
						a0_wr[1948]   <= x1948_in;                    
						a0_wr[1949]   <= x1949_in;                    
						a0_wr[1950]   <= x1950_in;                    
						a0_wr[1951]   <= x1951_in;                    
						a0_wr[1952]   <= x1952_in;                    
						a0_wr[1953]   <= x1953_in;                    
						a0_wr[1954]   <= x1954_in;                    
						a0_wr[1955]   <= x1955_in;                    
						a0_wr[1956]   <= x1956_in;                    
						a0_wr[1957]   <= x1957_in;                    
						a0_wr[1958]   <= x1958_in;                    
						a0_wr[1959]   <= x1959_in;                    
						a0_wr[1960]   <= x1960_in;                    
						a0_wr[1961]   <= x1961_in;                    
						a0_wr[1962]   <= x1962_in;                    
						a0_wr[1963]   <= x1963_in;                    
						a0_wr[1964]   <= x1964_in;                    
						a0_wr[1965]   <= x1965_in;                    
						a0_wr[1966]   <= x1966_in;                    
						a0_wr[1967]   <= x1967_in;                    
						a0_wr[1968]   <= x1968_in;                    
						a0_wr[1969]   <= x1969_in;                    
						a0_wr[1970]   <= x1970_in;                    
						a0_wr[1971]   <= x1971_in;                    
						a0_wr[1972]   <= x1972_in;                    
						a0_wr[1973]   <= x1973_in;                    
						a0_wr[1974]   <= x1974_in;                    
						a0_wr[1975]   <= x1975_in;                    
						a0_wr[1976]   <= x1976_in;                    
						a0_wr[1977]   <= x1977_in;                    
						a0_wr[1978]   <= x1978_in;                    
						a0_wr[1979]   <= x1979_in;                    
						a0_wr[1980]   <= x1980_in;                    
						a0_wr[1981]   <= x1981_in;                    
						a0_wr[1982]   <= x1982_in;                    
						a0_wr[1983]   <= x1983_in;                    
						a0_wr[1984]   <= x1984_in;                    
						a0_wr[1985]   <= x1985_in;                    
						a0_wr[1986]   <= x1986_in;                    
						a0_wr[1987]   <= x1987_in;                    
						a0_wr[1988]   <= x1988_in;                    
						a0_wr[1989]   <= x1989_in;                    
						a0_wr[1990]   <= x1990_in;                    
						a0_wr[1991]   <= x1991_in;                    
						a0_wr[1992]   <= x1992_in;                    
						a0_wr[1993]   <= x1993_in;                    
						a0_wr[1994]   <= x1994_in;                    
						a0_wr[1995]   <= x1995_in;                    
						a0_wr[1996]   <= x1996_in;                    
						a0_wr[1997]   <= x1997_in;                    
						a0_wr[1998]   <= x1998_in;                    
						a0_wr[1999]   <= x1999_in;                    
						a0_wr[2000]   <= x2000_in;                    
						a0_wr[2001]   <= x2001_in;                    
						a0_wr[2002]   <= x2002_in;                    
						a0_wr[2003]   <= x2003_in;                    
						a0_wr[2004]   <= x2004_in;                    
						a0_wr[2005]   <= x2005_in;                    
						a0_wr[2006]   <= x2006_in;                    
						a0_wr[2007]   <= x2007_in;                    
						a0_wr[2008]   <= x2008_in;                    
						a0_wr[2009]   <= x2009_in;                    
						a0_wr[2010]   <= x2010_in;                    
						a0_wr[2011]   <= x2011_in;                    
						a0_wr[2012]   <= x2012_in;                    
						a0_wr[2013]   <= x2013_in;                    
						a0_wr[2014]   <= x2014_in;                    
						a0_wr[2015]   <= x2015_in;                    
						a0_wr[2016]   <= x2016_in;                    
						a0_wr[2017]   <= x2017_in;                    
						a0_wr[2018]   <= x2018_in;                    
						a0_wr[2019]   <= x2019_in;                    
						a0_wr[2020]   <= x2020_in;                    
						a0_wr[2021]   <= x2021_in;                    
						a0_wr[2022]   <= x2022_in;                    
						a0_wr[2023]   <= x2023_in;                    
						a0_wr[2024]   <= x2024_in;                    
						a0_wr[2025]   <= x2025_in;                    
						a0_wr[2026]   <= x2026_in;                    
						a0_wr[2027]   <= x2027_in;                    
						a0_wr[2028]   <= x2028_in;                    
						a0_wr[2029]   <= x2029_in;                    
						a0_wr[2030]   <= x2030_in;                    
						a0_wr[2031]   <= x2031_in;                    
						a0_wr[2032]   <= x2032_in;                    
						a0_wr[2033]   <= x2033_in;                    
						a0_wr[2034]   <= x2034_in;                    
						a0_wr[2035]   <= x2035_in;                    
						a0_wr[2036]   <= x2036_in;                    
						a0_wr[2037]   <= x2037_in;                    
						a0_wr[2038]   <= x2038_in;                    
						a0_wr[2039]   <= x2039_in;                    
						a0_wr[2040]   <= x2040_in;                    
						a0_wr[2041]   <= x2041_in;                    
						a0_wr[2042]   <= x2042_in;                    
						a0_wr[2043]   <= x2043_in;                    
						a0_wr[2044]   <= x2044_in;                    
						a0_wr[2045]   <= x2045_in;                    
						a0_wr[2046]   <= x2046_in;                    
						a0_wr[2047]   <= x2047_in;                    
					end
				end
			end

		//--- radix stage 0
			radix2 #(.width(width)) rd_st0_0   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[0]), .rdlo_in(a0_wr[1024]),  .coef_in(coef[0]), .rdup_out(a1_wr[0]), .rdlo_out(a1_wr[1024]));
			radix2 #(.width(width)) rd_st0_1   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[1]), .rdlo_in(a0_wr[1025]),  .coef_in(coef[1]), .rdup_out(a1_wr[1]), .rdlo_out(a1_wr[1025]));
			radix2 #(.width(width)) rd_st0_2   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[2]), .rdlo_in(a0_wr[1026]),  .coef_in(coef[2]), .rdup_out(a1_wr[2]), .rdlo_out(a1_wr[1026]));
			radix2 #(.width(width)) rd_st0_3   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[3]), .rdlo_in(a0_wr[1027]),  .coef_in(coef[3]), .rdup_out(a1_wr[3]), .rdlo_out(a1_wr[1027]));
			radix2 #(.width(width)) rd_st0_4   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[4]), .rdlo_in(a0_wr[1028]),  .coef_in(coef[4]), .rdup_out(a1_wr[4]), .rdlo_out(a1_wr[1028]));
			radix2 #(.width(width)) rd_st0_5   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[5]), .rdlo_in(a0_wr[1029]),  .coef_in(coef[5]), .rdup_out(a1_wr[5]), .rdlo_out(a1_wr[1029]));
			radix2 #(.width(width)) rd_st0_6   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[6]), .rdlo_in(a0_wr[1030]),  .coef_in(coef[6]), .rdup_out(a1_wr[6]), .rdlo_out(a1_wr[1030]));
			radix2 #(.width(width)) rd_st0_7   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[7]), .rdlo_in(a0_wr[1031]),  .coef_in(coef[7]), .rdup_out(a1_wr[7]), .rdlo_out(a1_wr[1031]));
			radix2 #(.width(width)) rd_st0_8   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[8]), .rdlo_in(a0_wr[1032]),  .coef_in(coef[8]), .rdup_out(a1_wr[8]), .rdlo_out(a1_wr[1032]));
			radix2 #(.width(width)) rd_st0_9   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[9]), .rdlo_in(a0_wr[1033]),  .coef_in(coef[9]), .rdup_out(a1_wr[9]), .rdlo_out(a1_wr[1033]));
			radix2 #(.width(width)) rd_st0_10  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[10]), .rdlo_in(a0_wr[1034]),  .coef_in(coef[10]), .rdup_out(a1_wr[10]), .rdlo_out(a1_wr[1034]));
			radix2 #(.width(width)) rd_st0_11  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[11]), .rdlo_in(a0_wr[1035]),  .coef_in(coef[11]), .rdup_out(a1_wr[11]), .rdlo_out(a1_wr[1035]));
			radix2 #(.width(width)) rd_st0_12  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[12]), .rdlo_in(a0_wr[1036]),  .coef_in(coef[12]), .rdup_out(a1_wr[12]), .rdlo_out(a1_wr[1036]));
			radix2 #(.width(width)) rd_st0_13  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[13]), .rdlo_in(a0_wr[1037]),  .coef_in(coef[13]), .rdup_out(a1_wr[13]), .rdlo_out(a1_wr[1037]));
			radix2 #(.width(width)) rd_st0_14  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[14]), .rdlo_in(a0_wr[1038]),  .coef_in(coef[14]), .rdup_out(a1_wr[14]), .rdlo_out(a1_wr[1038]));
			radix2 #(.width(width)) rd_st0_15  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[15]), .rdlo_in(a0_wr[1039]),  .coef_in(coef[15]), .rdup_out(a1_wr[15]), .rdlo_out(a1_wr[1039]));
			radix2 #(.width(width)) rd_st0_16  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[16]), .rdlo_in(a0_wr[1040]),  .coef_in(coef[16]), .rdup_out(a1_wr[16]), .rdlo_out(a1_wr[1040]));
			radix2 #(.width(width)) rd_st0_17  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[17]), .rdlo_in(a0_wr[1041]),  .coef_in(coef[17]), .rdup_out(a1_wr[17]), .rdlo_out(a1_wr[1041]));
			radix2 #(.width(width)) rd_st0_18  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[18]), .rdlo_in(a0_wr[1042]),  .coef_in(coef[18]), .rdup_out(a1_wr[18]), .rdlo_out(a1_wr[1042]));
			radix2 #(.width(width)) rd_st0_19  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[19]), .rdlo_in(a0_wr[1043]),  .coef_in(coef[19]), .rdup_out(a1_wr[19]), .rdlo_out(a1_wr[1043]));
			radix2 #(.width(width)) rd_st0_20  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[20]), .rdlo_in(a0_wr[1044]),  .coef_in(coef[20]), .rdup_out(a1_wr[20]), .rdlo_out(a1_wr[1044]));
			radix2 #(.width(width)) rd_st0_21  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[21]), .rdlo_in(a0_wr[1045]),  .coef_in(coef[21]), .rdup_out(a1_wr[21]), .rdlo_out(a1_wr[1045]));
			radix2 #(.width(width)) rd_st0_22  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[22]), .rdlo_in(a0_wr[1046]),  .coef_in(coef[22]), .rdup_out(a1_wr[22]), .rdlo_out(a1_wr[1046]));
			radix2 #(.width(width)) rd_st0_23  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[23]), .rdlo_in(a0_wr[1047]),  .coef_in(coef[23]), .rdup_out(a1_wr[23]), .rdlo_out(a1_wr[1047]));
			radix2 #(.width(width)) rd_st0_24  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[24]), .rdlo_in(a0_wr[1048]),  .coef_in(coef[24]), .rdup_out(a1_wr[24]), .rdlo_out(a1_wr[1048]));
			radix2 #(.width(width)) rd_st0_25  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[25]), .rdlo_in(a0_wr[1049]),  .coef_in(coef[25]), .rdup_out(a1_wr[25]), .rdlo_out(a1_wr[1049]));
			radix2 #(.width(width)) rd_st0_26  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[26]), .rdlo_in(a0_wr[1050]),  .coef_in(coef[26]), .rdup_out(a1_wr[26]), .rdlo_out(a1_wr[1050]));
			radix2 #(.width(width)) rd_st0_27  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[27]), .rdlo_in(a0_wr[1051]),  .coef_in(coef[27]), .rdup_out(a1_wr[27]), .rdlo_out(a1_wr[1051]));
			radix2 #(.width(width)) rd_st0_28  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[28]), .rdlo_in(a0_wr[1052]),  .coef_in(coef[28]), .rdup_out(a1_wr[28]), .rdlo_out(a1_wr[1052]));
			radix2 #(.width(width)) rd_st0_29  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[29]), .rdlo_in(a0_wr[1053]),  .coef_in(coef[29]), .rdup_out(a1_wr[29]), .rdlo_out(a1_wr[1053]));
			radix2 #(.width(width)) rd_st0_30  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[30]), .rdlo_in(a0_wr[1054]),  .coef_in(coef[30]), .rdup_out(a1_wr[30]), .rdlo_out(a1_wr[1054]));
			radix2 #(.width(width)) rd_st0_31  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[31]), .rdlo_in(a0_wr[1055]),  .coef_in(coef[31]), .rdup_out(a1_wr[31]), .rdlo_out(a1_wr[1055]));
			radix2 #(.width(width)) rd_st0_32  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[32]), .rdlo_in(a0_wr[1056]),  .coef_in(coef[32]), .rdup_out(a1_wr[32]), .rdlo_out(a1_wr[1056]));
			radix2 #(.width(width)) rd_st0_33  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[33]), .rdlo_in(a0_wr[1057]),  .coef_in(coef[33]), .rdup_out(a1_wr[33]), .rdlo_out(a1_wr[1057]));
			radix2 #(.width(width)) rd_st0_34  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[34]), .rdlo_in(a0_wr[1058]),  .coef_in(coef[34]), .rdup_out(a1_wr[34]), .rdlo_out(a1_wr[1058]));
			radix2 #(.width(width)) rd_st0_35  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[35]), .rdlo_in(a0_wr[1059]),  .coef_in(coef[35]), .rdup_out(a1_wr[35]), .rdlo_out(a1_wr[1059]));
			radix2 #(.width(width)) rd_st0_36  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[36]), .rdlo_in(a0_wr[1060]),  .coef_in(coef[36]), .rdup_out(a1_wr[36]), .rdlo_out(a1_wr[1060]));
			radix2 #(.width(width)) rd_st0_37  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[37]), .rdlo_in(a0_wr[1061]),  .coef_in(coef[37]), .rdup_out(a1_wr[37]), .rdlo_out(a1_wr[1061]));
			radix2 #(.width(width)) rd_st0_38  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[38]), .rdlo_in(a0_wr[1062]),  .coef_in(coef[38]), .rdup_out(a1_wr[38]), .rdlo_out(a1_wr[1062]));
			radix2 #(.width(width)) rd_st0_39  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[39]), .rdlo_in(a0_wr[1063]),  .coef_in(coef[39]), .rdup_out(a1_wr[39]), .rdlo_out(a1_wr[1063]));
			radix2 #(.width(width)) rd_st0_40  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[40]), .rdlo_in(a0_wr[1064]),  .coef_in(coef[40]), .rdup_out(a1_wr[40]), .rdlo_out(a1_wr[1064]));
			radix2 #(.width(width)) rd_st0_41  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[41]), .rdlo_in(a0_wr[1065]),  .coef_in(coef[41]), .rdup_out(a1_wr[41]), .rdlo_out(a1_wr[1065]));
			radix2 #(.width(width)) rd_st0_42  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[42]), .rdlo_in(a0_wr[1066]),  .coef_in(coef[42]), .rdup_out(a1_wr[42]), .rdlo_out(a1_wr[1066]));
			radix2 #(.width(width)) rd_st0_43  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[43]), .rdlo_in(a0_wr[1067]),  .coef_in(coef[43]), .rdup_out(a1_wr[43]), .rdlo_out(a1_wr[1067]));
			radix2 #(.width(width)) rd_st0_44  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[44]), .rdlo_in(a0_wr[1068]),  .coef_in(coef[44]), .rdup_out(a1_wr[44]), .rdlo_out(a1_wr[1068]));
			radix2 #(.width(width)) rd_st0_45  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[45]), .rdlo_in(a0_wr[1069]),  .coef_in(coef[45]), .rdup_out(a1_wr[45]), .rdlo_out(a1_wr[1069]));
			radix2 #(.width(width)) rd_st0_46  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[46]), .rdlo_in(a0_wr[1070]),  .coef_in(coef[46]), .rdup_out(a1_wr[46]), .rdlo_out(a1_wr[1070]));
			radix2 #(.width(width)) rd_st0_47  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[47]), .rdlo_in(a0_wr[1071]),  .coef_in(coef[47]), .rdup_out(a1_wr[47]), .rdlo_out(a1_wr[1071]));
			radix2 #(.width(width)) rd_st0_48  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[48]), .rdlo_in(a0_wr[1072]),  .coef_in(coef[48]), .rdup_out(a1_wr[48]), .rdlo_out(a1_wr[1072]));
			radix2 #(.width(width)) rd_st0_49  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[49]), .rdlo_in(a0_wr[1073]),  .coef_in(coef[49]), .rdup_out(a1_wr[49]), .rdlo_out(a1_wr[1073]));
			radix2 #(.width(width)) rd_st0_50  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[50]), .rdlo_in(a0_wr[1074]),  .coef_in(coef[50]), .rdup_out(a1_wr[50]), .rdlo_out(a1_wr[1074]));
			radix2 #(.width(width)) rd_st0_51  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[51]), .rdlo_in(a0_wr[1075]),  .coef_in(coef[51]), .rdup_out(a1_wr[51]), .rdlo_out(a1_wr[1075]));
			radix2 #(.width(width)) rd_st0_52  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[52]), .rdlo_in(a0_wr[1076]),  .coef_in(coef[52]), .rdup_out(a1_wr[52]), .rdlo_out(a1_wr[1076]));
			radix2 #(.width(width)) rd_st0_53  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[53]), .rdlo_in(a0_wr[1077]),  .coef_in(coef[53]), .rdup_out(a1_wr[53]), .rdlo_out(a1_wr[1077]));
			radix2 #(.width(width)) rd_st0_54  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[54]), .rdlo_in(a0_wr[1078]),  .coef_in(coef[54]), .rdup_out(a1_wr[54]), .rdlo_out(a1_wr[1078]));
			radix2 #(.width(width)) rd_st0_55  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[55]), .rdlo_in(a0_wr[1079]),  .coef_in(coef[55]), .rdup_out(a1_wr[55]), .rdlo_out(a1_wr[1079]));
			radix2 #(.width(width)) rd_st0_56  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[56]), .rdlo_in(a0_wr[1080]),  .coef_in(coef[56]), .rdup_out(a1_wr[56]), .rdlo_out(a1_wr[1080]));
			radix2 #(.width(width)) rd_st0_57  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[57]), .rdlo_in(a0_wr[1081]),  .coef_in(coef[57]), .rdup_out(a1_wr[57]), .rdlo_out(a1_wr[1081]));
			radix2 #(.width(width)) rd_st0_58  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[58]), .rdlo_in(a0_wr[1082]),  .coef_in(coef[58]), .rdup_out(a1_wr[58]), .rdlo_out(a1_wr[1082]));
			radix2 #(.width(width)) rd_st0_59  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[59]), .rdlo_in(a0_wr[1083]),  .coef_in(coef[59]), .rdup_out(a1_wr[59]), .rdlo_out(a1_wr[1083]));
			radix2 #(.width(width)) rd_st0_60  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[60]), .rdlo_in(a0_wr[1084]),  .coef_in(coef[60]), .rdup_out(a1_wr[60]), .rdlo_out(a1_wr[1084]));
			radix2 #(.width(width)) rd_st0_61  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[61]), .rdlo_in(a0_wr[1085]),  .coef_in(coef[61]), .rdup_out(a1_wr[61]), .rdlo_out(a1_wr[1085]));
			radix2 #(.width(width)) rd_st0_62  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[62]), .rdlo_in(a0_wr[1086]),  .coef_in(coef[62]), .rdup_out(a1_wr[62]), .rdlo_out(a1_wr[1086]));
			radix2 #(.width(width)) rd_st0_63  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[63]), .rdlo_in(a0_wr[1087]),  .coef_in(coef[63]), .rdup_out(a1_wr[63]), .rdlo_out(a1_wr[1087]));
			radix2 #(.width(width)) rd_st0_64  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[64]), .rdlo_in(a0_wr[1088]),  .coef_in(coef[64]), .rdup_out(a1_wr[64]), .rdlo_out(a1_wr[1088]));
			radix2 #(.width(width)) rd_st0_65  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[65]), .rdlo_in(a0_wr[1089]),  .coef_in(coef[65]), .rdup_out(a1_wr[65]), .rdlo_out(a1_wr[1089]));
			radix2 #(.width(width)) rd_st0_66  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[66]), .rdlo_in(a0_wr[1090]),  .coef_in(coef[66]), .rdup_out(a1_wr[66]), .rdlo_out(a1_wr[1090]));
			radix2 #(.width(width)) rd_st0_67  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[67]), .rdlo_in(a0_wr[1091]),  .coef_in(coef[67]), .rdup_out(a1_wr[67]), .rdlo_out(a1_wr[1091]));
			radix2 #(.width(width)) rd_st0_68  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[68]), .rdlo_in(a0_wr[1092]),  .coef_in(coef[68]), .rdup_out(a1_wr[68]), .rdlo_out(a1_wr[1092]));
			radix2 #(.width(width)) rd_st0_69  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[69]), .rdlo_in(a0_wr[1093]),  .coef_in(coef[69]), .rdup_out(a1_wr[69]), .rdlo_out(a1_wr[1093]));
			radix2 #(.width(width)) rd_st0_70  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[70]), .rdlo_in(a0_wr[1094]),  .coef_in(coef[70]), .rdup_out(a1_wr[70]), .rdlo_out(a1_wr[1094]));
			radix2 #(.width(width)) rd_st0_71  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[71]), .rdlo_in(a0_wr[1095]),  .coef_in(coef[71]), .rdup_out(a1_wr[71]), .rdlo_out(a1_wr[1095]));
			radix2 #(.width(width)) rd_st0_72  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[72]), .rdlo_in(a0_wr[1096]),  .coef_in(coef[72]), .rdup_out(a1_wr[72]), .rdlo_out(a1_wr[1096]));
			radix2 #(.width(width)) rd_st0_73  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[73]), .rdlo_in(a0_wr[1097]),  .coef_in(coef[73]), .rdup_out(a1_wr[73]), .rdlo_out(a1_wr[1097]));
			radix2 #(.width(width)) rd_st0_74  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[74]), .rdlo_in(a0_wr[1098]),  .coef_in(coef[74]), .rdup_out(a1_wr[74]), .rdlo_out(a1_wr[1098]));
			radix2 #(.width(width)) rd_st0_75  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[75]), .rdlo_in(a0_wr[1099]),  .coef_in(coef[75]), .rdup_out(a1_wr[75]), .rdlo_out(a1_wr[1099]));
			radix2 #(.width(width)) rd_st0_76  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[76]), .rdlo_in(a0_wr[1100]),  .coef_in(coef[76]), .rdup_out(a1_wr[76]), .rdlo_out(a1_wr[1100]));
			radix2 #(.width(width)) rd_st0_77  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[77]), .rdlo_in(a0_wr[1101]),  .coef_in(coef[77]), .rdup_out(a1_wr[77]), .rdlo_out(a1_wr[1101]));
			radix2 #(.width(width)) rd_st0_78  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[78]), .rdlo_in(a0_wr[1102]),  .coef_in(coef[78]), .rdup_out(a1_wr[78]), .rdlo_out(a1_wr[1102]));
			radix2 #(.width(width)) rd_st0_79  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[79]), .rdlo_in(a0_wr[1103]),  .coef_in(coef[79]), .rdup_out(a1_wr[79]), .rdlo_out(a1_wr[1103]));
			radix2 #(.width(width)) rd_st0_80  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[80]), .rdlo_in(a0_wr[1104]),  .coef_in(coef[80]), .rdup_out(a1_wr[80]), .rdlo_out(a1_wr[1104]));
			radix2 #(.width(width)) rd_st0_81  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[81]), .rdlo_in(a0_wr[1105]),  .coef_in(coef[81]), .rdup_out(a1_wr[81]), .rdlo_out(a1_wr[1105]));
			radix2 #(.width(width)) rd_st0_82  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[82]), .rdlo_in(a0_wr[1106]),  .coef_in(coef[82]), .rdup_out(a1_wr[82]), .rdlo_out(a1_wr[1106]));
			radix2 #(.width(width)) rd_st0_83  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[83]), .rdlo_in(a0_wr[1107]),  .coef_in(coef[83]), .rdup_out(a1_wr[83]), .rdlo_out(a1_wr[1107]));
			radix2 #(.width(width)) rd_st0_84  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[84]), .rdlo_in(a0_wr[1108]),  .coef_in(coef[84]), .rdup_out(a1_wr[84]), .rdlo_out(a1_wr[1108]));
			radix2 #(.width(width)) rd_st0_85  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[85]), .rdlo_in(a0_wr[1109]),  .coef_in(coef[85]), .rdup_out(a1_wr[85]), .rdlo_out(a1_wr[1109]));
			radix2 #(.width(width)) rd_st0_86  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[86]), .rdlo_in(a0_wr[1110]),  .coef_in(coef[86]), .rdup_out(a1_wr[86]), .rdlo_out(a1_wr[1110]));
			radix2 #(.width(width)) rd_st0_87  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[87]), .rdlo_in(a0_wr[1111]),  .coef_in(coef[87]), .rdup_out(a1_wr[87]), .rdlo_out(a1_wr[1111]));
			radix2 #(.width(width)) rd_st0_88  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[88]), .rdlo_in(a0_wr[1112]),  .coef_in(coef[88]), .rdup_out(a1_wr[88]), .rdlo_out(a1_wr[1112]));
			radix2 #(.width(width)) rd_st0_89  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[89]), .rdlo_in(a0_wr[1113]),  .coef_in(coef[89]), .rdup_out(a1_wr[89]), .rdlo_out(a1_wr[1113]));
			radix2 #(.width(width)) rd_st0_90  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[90]), .rdlo_in(a0_wr[1114]),  .coef_in(coef[90]), .rdup_out(a1_wr[90]), .rdlo_out(a1_wr[1114]));
			radix2 #(.width(width)) rd_st0_91  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[91]), .rdlo_in(a0_wr[1115]),  .coef_in(coef[91]), .rdup_out(a1_wr[91]), .rdlo_out(a1_wr[1115]));
			radix2 #(.width(width)) rd_st0_92  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[92]), .rdlo_in(a0_wr[1116]),  .coef_in(coef[92]), .rdup_out(a1_wr[92]), .rdlo_out(a1_wr[1116]));
			radix2 #(.width(width)) rd_st0_93  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[93]), .rdlo_in(a0_wr[1117]),  .coef_in(coef[93]), .rdup_out(a1_wr[93]), .rdlo_out(a1_wr[1117]));
			radix2 #(.width(width)) rd_st0_94  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[94]), .rdlo_in(a0_wr[1118]),  .coef_in(coef[94]), .rdup_out(a1_wr[94]), .rdlo_out(a1_wr[1118]));
			radix2 #(.width(width)) rd_st0_95  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[95]), .rdlo_in(a0_wr[1119]),  .coef_in(coef[95]), .rdup_out(a1_wr[95]), .rdlo_out(a1_wr[1119]));
			radix2 #(.width(width)) rd_st0_96  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[96]), .rdlo_in(a0_wr[1120]),  .coef_in(coef[96]), .rdup_out(a1_wr[96]), .rdlo_out(a1_wr[1120]));
			radix2 #(.width(width)) rd_st0_97  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[97]), .rdlo_in(a0_wr[1121]),  .coef_in(coef[97]), .rdup_out(a1_wr[97]), .rdlo_out(a1_wr[1121]));
			radix2 #(.width(width)) rd_st0_98  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[98]), .rdlo_in(a0_wr[1122]),  .coef_in(coef[98]), .rdup_out(a1_wr[98]), .rdlo_out(a1_wr[1122]));
			radix2 #(.width(width)) rd_st0_99  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[99]), .rdlo_in(a0_wr[1123]),  .coef_in(coef[99]), .rdup_out(a1_wr[99]), .rdlo_out(a1_wr[1123]));
			radix2 #(.width(width)) rd_st0_100  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[100]), .rdlo_in(a0_wr[1124]),  .coef_in(coef[100]), .rdup_out(a1_wr[100]), .rdlo_out(a1_wr[1124]));
			radix2 #(.width(width)) rd_st0_101  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[101]), .rdlo_in(a0_wr[1125]),  .coef_in(coef[101]), .rdup_out(a1_wr[101]), .rdlo_out(a1_wr[1125]));
			radix2 #(.width(width)) rd_st0_102  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[102]), .rdlo_in(a0_wr[1126]),  .coef_in(coef[102]), .rdup_out(a1_wr[102]), .rdlo_out(a1_wr[1126]));
			radix2 #(.width(width)) rd_st0_103  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[103]), .rdlo_in(a0_wr[1127]),  .coef_in(coef[103]), .rdup_out(a1_wr[103]), .rdlo_out(a1_wr[1127]));
			radix2 #(.width(width)) rd_st0_104  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[104]), .rdlo_in(a0_wr[1128]),  .coef_in(coef[104]), .rdup_out(a1_wr[104]), .rdlo_out(a1_wr[1128]));
			radix2 #(.width(width)) rd_st0_105  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[105]), .rdlo_in(a0_wr[1129]),  .coef_in(coef[105]), .rdup_out(a1_wr[105]), .rdlo_out(a1_wr[1129]));
			radix2 #(.width(width)) rd_st0_106  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[106]), .rdlo_in(a0_wr[1130]),  .coef_in(coef[106]), .rdup_out(a1_wr[106]), .rdlo_out(a1_wr[1130]));
			radix2 #(.width(width)) rd_st0_107  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[107]), .rdlo_in(a0_wr[1131]),  .coef_in(coef[107]), .rdup_out(a1_wr[107]), .rdlo_out(a1_wr[1131]));
			radix2 #(.width(width)) rd_st0_108  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[108]), .rdlo_in(a0_wr[1132]),  .coef_in(coef[108]), .rdup_out(a1_wr[108]), .rdlo_out(a1_wr[1132]));
			radix2 #(.width(width)) rd_st0_109  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[109]), .rdlo_in(a0_wr[1133]),  .coef_in(coef[109]), .rdup_out(a1_wr[109]), .rdlo_out(a1_wr[1133]));
			radix2 #(.width(width)) rd_st0_110  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[110]), .rdlo_in(a0_wr[1134]),  .coef_in(coef[110]), .rdup_out(a1_wr[110]), .rdlo_out(a1_wr[1134]));
			radix2 #(.width(width)) rd_st0_111  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[111]), .rdlo_in(a0_wr[1135]),  .coef_in(coef[111]), .rdup_out(a1_wr[111]), .rdlo_out(a1_wr[1135]));
			radix2 #(.width(width)) rd_st0_112  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[112]), .rdlo_in(a0_wr[1136]),  .coef_in(coef[112]), .rdup_out(a1_wr[112]), .rdlo_out(a1_wr[1136]));
			radix2 #(.width(width)) rd_st0_113  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[113]), .rdlo_in(a0_wr[1137]),  .coef_in(coef[113]), .rdup_out(a1_wr[113]), .rdlo_out(a1_wr[1137]));
			radix2 #(.width(width)) rd_st0_114  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[114]), .rdlo_in(a0_wr[1138]),  .coef_in(coef[114]), .rdup_out(a1_wr[114]), .rdlo_out(a1_wr[1138]));
			radix2 #(.width(width)) rd_st0_115  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[115]), .rdlo_in(a0_wr[1139]),  .coef_in(coef[115]), .rdup_out(a1_wr[115]), .rdlo_out(a1_wr[1139]));
			radix2 #(.width(width)) rd_st0_116  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[116]), .rdlo_in(a0_wr[1140]),  .coef_in(coef[116]), .rdup_out(a1_wr[116]), .rdlo_out(a1_wr[1140]));
			radix2 #(.width(width)) rd_st0_117  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[117]), .rdlo_in(a0_wr[1141]),  .coef_in(coef[117]), .rdup_out(a1_wr[117]), .rdlo_out(a1_wr[1141]));
			radix2 #(.width(width)) rd_st0_118  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[118]), .rdlo_in(a0_wr[1142]),  .coef_in(coef[118]), .rdup_out(a1_wr[118]), .rdlo_out(a1_wr[1142]));
			radix2 #(.width(width)) rd_st0_119  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[119]), .rdlo_in(a0_wr[1143]),  .coef_in(coef[119]), .rdup_out(a1_wr[119]), .rdlo_out(a1_wr[1143]));
			radix2 #(.width(width)) rd_st0_120  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[120]), .rdlo_in(a0_wr[1144]),  .coef_in(coef[120]), .rdup_out(a1_wr[120]), .rdlo_out(a1_wr[1144]));
			radix2 #(.width(width)) rd_st0_121  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[121]), .rdlo_in(a0_wr[1145]),  .coef_in(coef[121]), .rdup_out(a1_wr[121]), .rdlo_out(a1_wr[1145]));
			radix2 #(.width(width)) rd_st0_122  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[122]), .rdlo_in(a0_wr[1146]),  .coef_in(coef[122]), .rdup_out(a1_wr[122]), .rdlo_out(a1_wr[1146]));
			radix2 #(.width(width)) rd_st0_123  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[123]), .rdlo_in(a0_wr[1147]),  .coef_in(coef[123]), .rdup_out(a1_wr[123]), .rdlo_out(a1_wr[1147]));
			radix2 #(.width(width)) rd_st0_124  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[124]), .rdlo_in(a0_wr[1148]),  .coef_in(coef[124]), .rdup_out(a1_wr[124]), .rdlo_out(a1_wr[1148]));
			radix2 #(.width(width)) rd_st0_125  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[125]), .rdlo_in(a0_wr[1149]),  .coef_in(coef[125]), .rdup_out(a1_wr[125]), .rdlo_out(a1_wr[1149]));
			radix2 #(.width(width)) rd_st0_126  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[126]), .rdlo_in(a0_wr[1150]),  .coef_in(coef[126]), .rdup_out(a1_wr[126]), .rdlo_out(a1_wr[1150]));
			radix2 #(.width(width)) rd_st0_127  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[127]), .rdlo_in(a0_wr[1151]),  .coef_in(coef[127]), .rdup_out(a1_wr[127]), .rdlo_out(a1_wr[1151]));
			radix2 #(.width(width)) rd_st0_128  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[128]), .rdlo_in(a0_wr[1152]),  .coef_in(coef[128]), .rdup_out(a1_wr[128]), .rdlo_out(a1_wr[1152]));
			radix2 #(.width(width)) rd_st0_129  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[129]), .rdlo_in(a0_wr[1153]),  .coef_in(coef[129]), .rdup_out(a1_wr[129]), .rdlo_out(a1_wr[1153]));
			radix2 #(.width(width)) rd_st0_130  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[130]), .rdlo_in(a0_wr[1154]),  .coef_in(coef[130]), .rdup_out(a1_wr[130]), .rdlo_out(a1_wr[1154]));
			radix2 #(.width(width)) rd_st0_131  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[131]), .rdlo_in(a0_wr[1155]),  .coef_in(coef[131]), .rdup_out(a1_wr[131]), .rdlo_out(a1_wr[1155]));
			radix2 #(.width(width)) rd_st0_132  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[132]), .rdlo_in(a0_wr[1156]),  .coef_in(coef[132]), .rdup_out(a1_wr[132]), .rdlo_out(a1_wr[1156]));
			radix2 #(.width(width)) rd_st0_133  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[133]), .rdlo_in(a0_wr[1157]),  .coef_in(coef[133]), .rdup_out(a1_wr[133]), .rdlo_out(a1_wr[1157]));
			radix2 #(.width(width)) rd_st0_134  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[134]), .rdlo_in(a0_wr[1158]),  .coef_in(coef[134]), .rdup_out(a1_wr[134]), .rdlo_out(a1_wr[1158]));
			radix2 #(.width(width)) rd_st0_135  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[135]), .rdlo_in(a0_wr[1159]),  .coef_in(coef[135]), .rdup_out(a1_wr[135]), .rdlo_out(a1_wr[1159]));
			radix2 #(.width(width)) rd_st0_136  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[136]), .rdlo_in(a0_wr[1160]),  .coef_in(coef[136]), .rdup_out(a1_wr[136]), .rdlo_out(a1_wr[1160]));
			radix2 #(.width(width)) rd_st0_137  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[137]), .rdlo_in(a0_wr[1161]),  .coef_in(coef[137]), .rdup_out(a1_wr[137]), .rdlo_out(a1_wr[1161]));
			radix2 #(.width(width)) rd_st0_138  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[138]), .rdlo_in(a0_wr[1162]),  .coef_in(coef[138]), .rdup_out(a1_wr[138]), .rdlo_out(a1_wr[1162]));
			radix2 #(.width(width)) rd_st0_139  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[139]), .rdlo_in(a0_wr[1163]),  .coef_in(coef[139]), .rdup_out(a1_wr[139]), .rdlo_out(a1_wr[1163]));
			radix2 #(.width(width)) rd_st0_140  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[140]), .rdlo_in(a0_wr[1164]),  .coef_in(coef[140]), .rdup_out(a1_wr[140]), .rdlo_out(a1_wr[1164]));
			radix2 #(.width(width)) rd_st0_141  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[141]), .rdlo_in(a0_wr[1165]),  .coef_in(coef[141]), .rdup_out(a1_wr[141]), .rdlo_out(a1_wr[1165]));
			radix2 #(.width(width)) rd_st0_142  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[142]), .rdlo_in(a0_wr[1166]),  .coef_in(coef[142]), .rdup_out(a1_wr[142]), .rdlo_out(a1_wr[1166]));
			radix2 #(.width(width)) rd_st0_143  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[143]), .rdlo_in(a0_wr[1167]),  .coef_in(coef[143]), .rdup_out(a1_wr[143]), .rdlo_out(a1_wr[1167]));
			radix2 #(.width(width)) rd_st0_144  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[144]), .rdlo_in(a0_wr[1168]),  .coef_in(coef[144]), .rdup_out(a1_wr[144]), .rdlo_out(a1_wr[1168]));
			radix2 #(.width(width)) rd_st0_145  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[145]), .rdlo_in(a0_wr[1169]),  .coef_in(coef[145]), .rdup_out(a1_wr[145]), .rdlo_out(a1_wr[1169]));
			radix2 #(.width(width)) rd_st0_146  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[146]), .rdlo_in(a0_wr[1170]),  .coef_in(coef[146]), .rdup_out(a1_wr[146]), .rdlo_out(a1_wr[1170]));
			radix2 #(.width(width)) rd_st0_147  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[147]), .rdlo_in(a0_wr[1171]),  .coef_in(coef[147]), .rdup_out(a1_wr[147]), .rdlo_out(a1_wr[1171]));
			radix2 #(.width(width)) rd_st0_148  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[148]), .rdlo_in(a0_wr[1172]),  .coef_in(coef[148]), .rdup_out(a1_wr[148]), .rdlo_out(a1_wr[1172]));
			radix2 #(.width(width)) rd_st0_149  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[149]), .rdlo_in(a0_wr[1173]),  .coef_in(coef[149]), .rdup_out(a1_wr[149]), .rdlo_out(a1_wr[1173]));
			radix2 #(.width(width)) rd_st0_150  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[150]), .rdlo_in(a0_wr[1174]),  .coef_in(coef[150]), .rdup_out(a1_wr[150]), .rdlo_out(a1_wr[1174]));
			radix2 #(.width(width)) rd_st0_151  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[151]), .rdlo_in(a0_wr[1175]),  .coef_in(coef[151]), .rdup_out(a1_wr[151]), .rdlo_out(a1_wr[1175]));
			radix2 #(.width(width)) rd_st0_152  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[152]), .rdlo_in(a0_wr[1176]),  .coef_in(coef[152]), .rdup_out(a1_wr[152]), .rdlo_out(a1_wr[1176]));
			radix2 #(.width(width)) rd_st0_153  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[153]), .rdlo_in(a0_wr[1177]),  .coef_in(coef[153]), .rdup_out(a1_wr[153]), .rdlo_out(a1_wr[1177]));
			radix2 #(.width(width)) rd_st0_154  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[154]), .rdlo_in(a0_wr[1178]),  .coef_in(coef[154]), .rdup_out(a1_wr[154]), .rdlo_out(a1_wr[1178]));
			radix2 #(.width(width)) rd_st0_155  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[155]), .rdlo_in(a0_wr[1179]),  .coef_in(coef[155]), .rdup_out(a1_wr[155]), .rdlo_out(a1_wr[1179]));
			radix2 #(.width(width)) rd_st0_156  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[156]), .rdlo_in(a0_wr[1180]),  .coef_in(coef[156]), .rdup_out(a1_wr[156]), .rdlo_out(a1_wr[1180]));
			radix2 #(.width(width)) rd_st0_157  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[157]), .rdlo_in(a0_wr[1181]),  .coef_in(coef[157]), .rdup_out(a1_wr[157]), .rdlo_out(a1_wr[1181]));
			radix2 #(.width(width)) rd_st0_158  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[158]), .rdlo_in(a0_wr[1182]),  .coef_in(coef[158]), .rdup_out(a1_wr[158]), .rdlo_out(a1_wr[1182]));
			radix2 #(.width(width)) rd_st0_159  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[159]), .rdlo_in(a0_wr[1183]),  .coef_in(coef[159]), .rdup_out(a1_wr[159]), .rdlo_out(a1_wr[1183]));
			radix2 #(.width(width)) rd_st0_160  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[160]), .rdlo_in(a0_wr[1184]),  .coef_in(coef[160]), .rdup_out(a1_wr[160]), .rdlo_out(a1_wr[1184]));
			radix2 #(.width(width)) rd_st0_161  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[161]), .rdlo_in(a0_wr[1185]),  .coef_in(coef[161]), .rdup_out(a1_wr[161]), .rdlo_out(a1_wr[1185]));
			radix2 #(.width(width)) rd_st0_162  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[162]), .rdlo_in(a0_wr[1186]),  .coef_in(coef[162]), .rdup_out(a1_wr[162]), .rdlo_out(a1_wr[1186]));
			radix2 #(.width(width)) rd_st0_163  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[163]), .rdlo_in(a0_wr[1187]),  .coef_in(coef[163]), .rdup_out(a1_wr[163]), .rdlo_out(a1_wr[1187]));
			radix2 #(.width(width)) rd_st0_164  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[164]), .rdlo_in(a0_wr[1188]),  .coef_in(coef[164]), .rdup_out(a1_wr[164]), .rdlo_out(a1_wr[1188]));
			radix2 #(.width(width)) rd_st0_165  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[165]), .rdlo_in(a0_wr[1189]),  .coef_in(coef[165]), .rdup_out(a1_wr[165]), .rdlo_out(a1_wr[1189]));
			radix2 #(.width(width)) rd_st0_166  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[166]), .rdlo_in(a0_wr[1190]),  .coef_in(coef[166]), .rdup_out(a1_wr[166]), .rdlo_out(a1_wr[1190]));
			radix2 #(.width(width)) rd_st0_167  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[167]), .rdlo_in(a0_wr[1191]),  .coef_in(coef[167]), .rdup_out(a1_wr[167]), .rdlo_out(a1_wr[1191]));
			radix2 #(.width(width)) rd_st0_168  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[168]), .rdlo_in(a0_wr[1192]),  .coef_in(coef[168]), .rdup_out(a1_wr[168]), .rdlo_out(a1_wr[1192]));
			radix2 #(.width(width)) rd_st0_169  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[169]), .rdlo_in(a0_wr[1193]),  .coef_in(coef[169]), .rdup_out(a1_wr[169]), .rdlo_out(a1_wr[1193]));
			radix2 #(.width(width)) rd_st0_170  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[170]), .rdlo_in(a0_wr[1194]),  .coef_in(coef[170]), .rdup_out(a1_wr[170]), .rdlo_out(a1_wr[1194]));
			radix2 #(.width(width)) rd_st0_171  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[171]), .rdlo_in(a0_wr[1195]),  .coef_in(coef[171]), .rdup_out(a1_wr[171]), .rdlo_out(a1_wr[1195]));
			radix2 #(.width(width)) rd_st0_172  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[172]), .rdlo_in(a0_wr[1196]),  .coef_in(coef[172]), .rdup_out(a1_wr[172]), .rdlo_out(a1_wr[1196]));
			radix2 #(.width(width)) rd_st0_173  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[173]), .rdlo_in(a0_wr[1197]),  .coef_in(coef[173]), .rdup_out(a1_wr[173]), .rdlo_out(a1_wr[1197]));
			radix2 #(.width(width)) rd_st0_174  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[174]), .rdlo_in(a0_wr[1198]),  .coef_in(coef[174]), .rdup_out(a1_wr[174]), .rdlo_out(a1_wr[1198]));
			radix2 #(.width(width)) rd_st0_175  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[175]), .rdlo_in(a0_wr[1199]),  .coef_in(coef[175]), .rdup_out(a1_wr[175]), .rdlo_out(a1_wr[1199]));
			radix2 #(.width(width)) rd_st0_176  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[176]), .rdlo_in(a0_wr[1200]),  .coef_in(coef[176]), .rdup_out(a1_wr[176]), .rdlo_out(a1_wr[1200]));
			radix2 #(.width(width)) rd_st0_177  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[177]), .rdlo_in(a0_wr[1201]),  .coef_in(coef[177]), .rdup_out(a1_wr[177]), .rdlo_out(a1_wr[1201]));
			radix2 #(.width(width)) rd_st0_178  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[178]), .rdlo_in(a0_wr[1202]),  .coef_in(coef[178]), .rdup_out(a1_wr[178]), .rdlo_out(a1_wr[1202]));
			radix2 #(.width(width)) rd_st0_179  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[179]), .rdlo_in(a0_wr[1203]),  .coef_in(coef[179]), .rdup_out(a1_wr[179]), .rdlo_out(a1_wr[1203]));
			radix2 #(.width(width)) rd_st0_180  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[180]), .rdlo_in(a0_wr[1204]),  .coef_in(coef[180]), .rdup_out(a1_wr[180]), .rdlo_out(a1_wr[1204]));
			radix2 #(.width(width)) rd_st0_181  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[181]), .rdlo_in(a0_wr[1205]),  .coef_in(coef[181]), .rdup_out(a1_wr[181]), .rdlo_out(a1_wr[1205]));
			radix2 #(.width(width)) rd_st0_182  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[182]), .rdlo_in(a0_wr[1206]),  .coef_in(coef[182]), .rdup_out(a1_wr[182]), .rdlo_out(a1_wr[1206]));
			radix2 #(.width(width)) rd_st0_183  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[183]), .rdlo_in(a0_wr[1207]),  .coef_in(coef[183]), .rdup_out(a1_wr[183]), .rdlo_out(a1_wr[1207]));
			radix2 #(.width(width)) rd_st0_184  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[184]), .rdlo_in(a0_wr[1208]),  .coef_in(coef[184]), .rdup_out(a1_wr[184]), .rdlo_out(a1_wr[1208]));
			radix2 #(.width(width)) rd_st0_185  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[185]), .rdlo_in(a0_wr[1209]),  .coef_in(coef[185]), .rdup_out(a1_wr[185]), .rdlo_out(a1_wr[1209]));
			radix2 #(.width(width)) rd_st0_186  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[186]), .rdlo_in(a0_wr[1210]),  .coef_in(coef[186]), .rdup_out(a1_wr[186]), .rdlo_out(a1_wr[1210]));
			radix2 #(.width(width)) rd_st0_187  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[187]), .rdlo_in(a0_wr[1211]),  .coef_in(coef[187]), .rdup_out(a1_wr[187]), .rdlo_out(a1_wr[1211]));
			radix2 #(.width(width)) rd_st0_188  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[188]), .rdlo_in(a0_wr[1212]),  .coef_in(coef[188]), .rdup_out(a1_wr[188]), .rdlo_out(a1_wr[1212]));
			radix2 #(.width(width)) rd_st0_189  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[189]), .rdlo_in(a0_wr[1213]),  .coef_in(coef[189]), .rdup_out(a1_wr[189]), .rdlo_out(a1_wr[1213]));
			radix2 #(.width(width)) rd_st0_190  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[190]), .rdlo_in(a0_wr[1214]),  .coef_in(coef[190]), .rdup_out(a1_wr[190]), .rdlo_out(a1_wr[1214]));
			radix2 #(.width(width)) rd_st0_191  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[191]), .rdlo_in(a0_wr[1215]),  .coef_in(coef[191]), .rdup_out(a1_wr[191]), .rdlo_out(a1_wr[1215]));
			radix2 #(.width(width)) rd_st0_192  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[192]), .rdlo_in(a0_wr[1216]),  .coef_in(coef[192]), .rdup_out(a1_wr[192]), .rdlo_out(a1_wr[1216]));
			radix2 #(.width(width)) rd_st0_193  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[193]), .rdlo_in(a0_wr[1217]),  .coef_in(coef[193]), .rdup_out(a1_wr[193]), .rdlo_out(a1_wr[1217]));
			radix2 #(.width(width)) rd_st0_194  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[194]), .rdlo_in(a0_wr[1218]),  .coef_in(coef[194]), .rdup_out(a1_wr[194]), .rdlo_out(a1_wr[1218]));
			radix2 #(.width(width)) rd_st0_195  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[195]), .rdlo_in(a0_wr[1219]),  .coef_in(coef[195]), .rdup_out(a1_wr[195]), .rdlo_out(a1_wr[1219]));
			radix2 #(.width(width)) rd_st0_196  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[196]), .rdlo_in(a0_wr[1220]),  .coef_in(coef[196]), .rdup_out(a1_wr[196]), .rdlo_out(a1_wr[1220]));
			radix2 #(.width(width)) rd_st0_197  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[197]), .rdlo_in(a0_wr[1221]),  .coef_in(coef[197]), .rdup_out(a1_wr[197]), .rdlo_out(a1_wr[1221]));
			radix2 #(.width(width)) rd_st0_198  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[198]), .rdlo_in(a0_wr[1222]),  .coef_in(coef[198]), .rdup_out(a1_wr[198]), .rdlo_out(a1_wr[1222]));
			radix2 #(.width(width)) rd_st0_199  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[199]), .rdlo_in(a0_wr[1223]),  .coef_in(coef[199]), .rdup_out(a1_wr[199]), .rdlo_out(a1_wr[1223]));
			radix2 #(.width(width)) rd_st0_200  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[200]), .rdlo_in(a0_wr[1224]),  .coef_in(coef[200]), .rdup_out(a1_wr[200]), .rdlo_out(a1_wr[1224]));
			radix2 #(.width(width)) rd_st0_201  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[201]), .rdlo_in(a0_wr[1225]),  .coef_in(coef[201]), .rdup_out(a1_wr[201]), .rdlo_out(a1_wr[1225]));
			radix2 #(.width(width)) rd_st0_202  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[202]), .rdlo_in(a0_wr[1226]),  .coef_in(coef[202]), .rdup_out(a1_wr[202]), .rdlo_out(a1_wr[1226]));
			radix2 #(.width(width)) rd_st0_203  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[203]), .rdlo_in(a0_wr[1227]),  .coef_in(coef[203]), .rdup_out(a1_wr[203]), .rdlo_out(a1_wr[1227]));
			radix2 #(.width(width)) rd_st0_204  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[204]), .rdlo_in(a0_wr[1228]),  .coef_in(coef[204]), .rdup_out(a1_wr[204]), .rdlo_out(a1_wr[1228]));
			radix2 #(.width(width)) rd_st0_205  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[205]), .rdlo_in(a0_wr[1229]),  .coef_in(coef[205]), .rdup_out(a1_wr[205]), .rdlo_out(a1_wr[1229]));
			radix2 #(.width(width)) rd_st0_206  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[206]), .rdlo_in(a0_wr[1230]),  .coef_in(coef[206]), .rdup_out(a1_wr[206]), .rdlo_out(a1_wr[1230]));
			radix2 #(.width(width)) rd_st0_207  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[207]), .rdlo_in(a0_wr[1231]),  .coef_in(coef[207]), .rdup_out(a1_wr[207]), .rdlo_out(a1_wr[1231]));
			radix2 #(.width(width)) rd_st0_208  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[208]), .rdlo_in(a0_wr[1232]),  .coef_in(coef[208]), .rdup_out(a1_wr[208]), .rdlo_out(a1_wr[1232]));
			radix2 #(.width(width)) rd_st0_209  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[209]), .rdlo_in(a0_wr[1233]),  .coef_in(coef[209]), .rdup_out(a1_wr[209]), .rdlo_out(a1_wr[1233]));
			radix2 #(.width(width)) rd_st0_210  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[210]), .rdlo_in(a0_wr[1234]),  .coef_in(coef[210]), .rdup_out(a1_wr[210]), .rdlo_out(a1_wr[1234]));
			radix2 #(.width(width)) rd_st0_211  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[211]), .rdlo_in(a0_wr[1235]),  .coef_in(coef[211]), .rdup_out(a1_wr[211]), .rdlo_out(a1_wr[1235]));
			radix2 #(.width(width)) rd_st0_212  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[212]), .rdlo_in(a0_wr[1236]),  .coef_in(coef[212]), .rdup_out(a1_wr[212]), .rdlo_out(a1_wr[1236]));
			radix2 #(.width(width)) rd_st0_213  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[213]), .rdlo_in(a0_wr[1237]),  .coef_in(coef[213]), .rdup_out(a1_wr[213]), .rdlo_out(a1_wr[1237]));
			radix2 #(.width(width)) rd_st0_214  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[214]), .rdlo_in(a0_wr[1238]),  .coef_in(coef[214]), .rdup_out(a1_wr[214]), .rdlo_out(a1_wr[1238]));
			radix2 #(.width(width)) rd_st0_215  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[215]), .rdlo_in(a0_wr[1239]),  .coef_in(coef[215]), .rdup_out(a1_wr[215]), .rdlo_out(a1_wr[1239]));
			radix2 #(.width(width)) rd_st0_216  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[216]), .rdlo_in(a0_wr[1240]),  .coef_in(coef[216]), .rdup_out(a1_wr[216]), .rdlo_out(a1_wr[1240]));
			radix2 #(.width(width)) rd_st0_217  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[217]), .rdlo_in(a0_wr[1241]),  .coef_in(coef[217]), .rdup_out(a1_wr[217]), .rdlo_out(a1_wr[1241]));
			radix2 #(.width(width)) rd_st0_218  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[218]), .rdlo_in(a0_wr[1242]),  .coef_in(coef[218]), .rdup_out(a1_wr[218]), .rdlo_out(a1_wr[1242]));
			radix2 #(.width(width)) rd_st0_219  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[219]), .rdlo_in(a0_wr[1243]),  .coef_in(coef[219]), .rdup_out(a1_wr[219]), .rdlo_out(a1_wr[1243]));
			radix2 #(.width(width)) rd_st0_220  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[220]), .rdlo_in(a0_wr[1244]),  .coef_in(coef[220]), .rdup_out(a1_wr[220]), .rdlo_out(a1_wr[1244]));
			radix2 #(.width(width)) rd_st0_221  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[221]), .rdlo_in(a0_wr[1245]),  .coef_in(coef[221]), .rdup_out(a1_wr[221]), .rdlo_out(a1_wr[1245]));
			radix2 #(.width(width)) rd_st0_222  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[222]), .rdlo_in(a0_wr[1246]),  .coef_in(coef[222]), .rdup_out(a1_wr[222]), .rdlo_out(a1_wr[1246]));
			radix2 #(.width(width)) rd_st0_223  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[223]), .rdlo_in(a0_wr[1247]),  .coef_in(coef[223]), .rdup_out(a1_wr[223]), .rdlo_out(a1_wr[1247]));
			radix2 #(.width(width)) rd_st0_224  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[224]), .rdlo_in(a0_wr[1248]),  .coef_in(coef[224]), .rdup_out(a1_wr[224]), .rdlo_out(a1_wr[1248]));
			radix2 #(.width(width)) rd_st0_225  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[225]), .rdlo_in(a0_wr[1249]),  .coef_in(coef[225]), .rdup_out(a1_wr[225]), .rdlo_out(a1_wr[1249]));
			radix2 #(.width(width)) rd_st0_226  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[226]), .rdlo_in(a0_wr[1250]),  .coef_in(coef[226]), .rdup_out(a1_wr[226]), .rdlo_out(a1_wr[1250]));
			radix2 #(.width(width)) rd_st0_227  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[227]), .rdlo_in(a0_wr[1251]),  .coef_in(coef[227]), .rdup_out(a1_wr[227]), .rdlo_out(a1_wr[1251]));
			radix2 #(.width(width)) rd_st0_228  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[228]), .rdlo_in(a0_wr[1252]),  .coef_in(coef[228]), .rdup_out(a1_wr[228]), .rdlo_out(a1_wr[1252]));
			radix2 #(.width(width)) rd_st0_229  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[229]), .rdlo_in(a0_wr[1253]),  .coef_in(coef[229]), .rdup_out(a1_wr[229]), .rdlo_out(a1_wr[1253]));
			radix2 #(.width(width)) rd_st0_230  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[230]), .rdlo_in(a0_wr[1254]),  .coef_in(coef[230]), .rdup_out(a1_wr[230]), .rdlo_out(a1_wr[1254]));
			radix2 #(.width(width)) rd_st0_231  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[231]), .rdlo_in(a0_wr[1255]),  .coef_in(coef[231]), .rdup_out(a1_wr[231]), .rdlo_out(a1_wr[1255]));
			radix2 #(.width(width)) rd_st0_232  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[232]), .rdlo_in(a0_wr[1256]),  .coef_in(coef[232]), .rdup_out(a1_wr[232]), .rdlo_out(a1_wr[1256]));
			radix2 #(.width(width)) rd_st0_233  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[233]), .rdlo_in(a0_wr[1257]),  .coef_in(coef[233]), .rdup_out(a1_wr[233]), .rdlo_out(a1_wr[1257]));
			radix2 #(.width(width)) rd_st0_234  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[234]), .rdlo_in(a0_wr[1258]),  .coef_in(coef[234]), .rdup_out(a1_wr[234]), .rdlo_out(a1_wr[1258]));
			radix2 #(.width(width)) rd_st0_235  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[235]), .rdlo_in(a0_wr[1259]),  .coef_in(coef[235]), .rdup_out(a1_wr[235]), .rdlo_out(a1_wr[1259]));
			radix2 #(.width(width)) rd_st0_236  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[236]), .rdlo_in(a0_wr[1260]),  .coef_in(coef[236]), .rdup_out(a1_wr[236]), .rdlo_out(a1_wr[1260]));
			radix2 #(.width(width)) rd_st0_237  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[237]), .rdlo_in(a0_wr[1261]),  .coef_in(coef[237]), .rdup_out(a1_wr[237]), .rdlo_out(a1_wr[1261]));
			radix2 #(.width(width)) rd_st0_238  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[238]), .rdlo_in(a0_wr[1262]),  .coef_in(coef[238]), .rdup_out(a1_wr[238]), .rdlo_out(a1_wr[1262]));
			radix2 #(.width(width)) rd_st0_239  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[239]), .rdlo_in(a0_wr[1263]),  .coef_in(coef[239]), .rdup_out(a1_wr[239]), .rdlo_out(a1_wr[1263]));
			radix2 #(.width(width)) rd_st0_240  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[240]), .rdlo_in(a0_wr[1264]),  .coef_in(coef[240]), .rdup_out(a1_wr[240]), .rdlo_out(a1_wr[1264]));
			radix2 #(.width(width)) rd_st0_241  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[241]), .rdlo_in(a0_wr[1265]),  .coef_in(coef[241]), .rdup_out(a1_wr[241]), .rdlo_out(a1_wr[1265]));
			radix2 #(.width(width)) rd_st0_242  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[242]), .rdlo_in(a0_wr[1266]),  .coef_in(coef[242]), .rdup_out(a1_wr[242]), .rdlo_out(a1_wr[1266]));
			radix2 #(.width(width)) rd_st0_243  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[243]), .rdlo_in(a0_wr[1267]),  .coef_in(coef[243]), .rdup_out(a1_wr[243]), .rdlo_out(a1_wr[1267]));
			radix2 #(.width(width)) rd_st0_244  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[244]), .rdlo_in(a0_wr[1268]),  .coef_in(coef[244]), .rdup_out(a1_wr[244]), .rdlo_out(a1_wr[1268]));
			radix2 #(.width(width)) rd_st0_245  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[245]), .rdlo_in(a0_wr[1269]),  .coef_in(coef[245]), .rdup_out(a1_wr[245]), .rdlo_out(a1_wr[1269]));
			radix2 #(.width(width)) rd_st0_246  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[246]), .rdlo_in(a0_wr[1270]),  .coef_in(coef[246]), .rdup_out(a1_wr[246]), .rdlo_out(a1_wr[1270]));
			radix2 #(.width(width)) rd_st0_247  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[247]), .rdlo_in(a0_wr[1271]),  .coef_in(coef[247]), .rdup_out(a1_wr[247]), .rdlo_out(a1_wr[1271]));
			radix2 #(.width(width)) rd_st0_248  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[248]), .rdlo_in(a0_wr[1272]),  .coef_in(coef[248]), .rdup_out(a1_wr[248]), .rdlo_out(a1_wr[1272]));
			radix2 #(.width(width)) rd_st0_249  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[249]), .rdlo_in(a0_wr[1273]),  .coef_in(coef[249]), .rdup_out(a1_wr[249]), .rdlo_out(a1_wr[1273]));
			radix2 #(.width(width)) rd_st0_250  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[250]), .rdlo_in(a0_wr[1274]),  .coef_in(coef[250]), .rdup_out(a1_wr[250]), .rdlo_out(a1_wr[1274]));
			radix2 #(.width(width)) rd_st0_251  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[251]), .rdlo_in(a0_wr[1275]),  .coef_in(coef[251]), .rdup_out(a1_wr[251]), .rdlo_out(a1_wr[1275]));
			radix2 #(.width(width)) rd_st0_252  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[252]), .rdlo_in(a0_wr[1276]),  .coef_in(coef[252]), .rdup_out(a1_wr[252]), .rdlo_out(a1_wr[1276]));
			radix2 #(.width(width)) rd_st0_253  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[253]), .rdlo_in(a0_wr[1277]),  .coef_in(coef[253]), .rdup_out(a1_wr[253]), .rdlo_out(a1_wr[1277]));
			radix2 #(.width(width)) rd_st0_254  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[254]), .rdlo_in(a0_wr[1278]),  .coef_in(coef[254]), .rdup_out(a1_wr[254]), .rdlo_out(a1_wr[1278]));
			radix2 #(.width(width)) rd_st0_255  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[255]), .rdlo_in(a0_wr[1279]),  .coef_in(coef[255]), .rdup_out(a1_wr[255]), .rdlo_out(a1_wr[1279]));
			radix2 #(.width(width)) rd_st0_256  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[256]), .rdlo_in(a0_wr[1280]),  .coef_in(coef[256]), .rdup_out(a1_wr[256]), .rdlo_out(a1_wr[1280]));
			radix2 #(.width(width)) rd_st0_257  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[257]), .rdlo_in(a0_wr[1281]),  .coef_in(coef[257]), .rdup_out(a1_wr[257]), .rdlo_out(a1_wr[1281]));
			radix2 #(.width(width)) rd_st0_258  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[258]), .rdlo_in(a0_wr[1282]),  .coef_in(coef[258]), .rdup_out(a1_wr[258]), .rdlo_out(a1_wr[1282]));
			radix2 #(.width(width)) rd_st0_259  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[259]), .rdlo_in(a0_wr[1283]),  .coef_in(coef[259]), .rdup_out(a1_wr[259]), .rdlo_out(a1_wr[1283]));
			radix2 #(.width(width)) rd_st0_260  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[260]), .rdlo_in(a0_wr[1284]),  .coef_in(coef[260]), .rdup_out(a1_wr[260]), .rdlo_out(a1_wr[1284]));
			radix2 #(.width(width)) rd_st0_261  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[261]), .rdlo_in(a0_wr[1285]),  .coef_in(coef[261]), .rdup_out(a1_wr[261]), .rdlo_out(a1_wr[1285]));
			radix2 #(.width(width)) rd_st0_262  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[262]), .rdlo_in(a0_wr[1286]),  .coef_in(coef[262]), .rdup_out(a1_wr[262]), .rdlo_out(a1_wr[1286]));
			radix2 #(.width(width)) rd_st0_263  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[263]), .rdlo_in(a0_wr[1287]),  .coef_in(coef[263]), .rdup_out(a1_wr[263]), .rdlo_out(a1_wr[1287]));
			radix2 #(.width(width)) rd_st0_264  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[264]), .rdlo_in(a0_wr[1288]),  .coef_in(coef[264]), .rdup_out(a1_wr[264]), .rdlo_out(a1_wr[1288]));
			radix2 #(.width(width)) rd_st0_265  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[265]), .rdlo_in(a0_wr[1289]),  .coef_in(coef[265]), .rdup_out(a1_wr[265]), .rdlo_out(a1_wr[1289]));
			radix2 #(.width(width)) rd_st0_266  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[266]), .rdlo_in(a0_wr[1290]),  .coef_in(coef[266]), .rdup_out(a1_wr[266]), .rdlo_out(a1_wr[1290]));
			radix2 #(.width(width)) rd_st0_267  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[267]), .rdlo_in(a0_wr[1291]),  .coef_in(coef[267]), .rdup_out(a1_wr[267]), .rdlo_out(a1_wr[1291]));
			radix2 #(.width(width)) rd_st0_268  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[268]), .rdlo_in(a0_wr[1292]),  .coef_in(coef[268]), .rdup_out(a1_wr[268]), .rdlo_out(a1_wr[1292]));
			radix2 #(.width(width)) rd_st0_269  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[269]), .rdlo_in(a0_wr[1293]),  .coef_in(coef[269]), .rdup_out(a1_wr[269]), .rdlo_out(a1_wr[1293]));
			radix2 #(.width(width)) rd_st0_270  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[270]), .rdlo_in(a0_wr[1294]),  .coef_in(coef[270]), .rdup_out(a1_wr[270]), .rdlo_out(a1_wr[1294]));
			radix2 #(.width(width)) rd_st0_271  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[271]), .rdlo_in(a0_wr[1295]),  .coef_in(coef[271]), .rdup_out(a1_wr[271]), .rdlo_out(a1_wr[1295]));
			radix2 #(.width(width)) rd_st0_272  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[272]), .rdlo_in(a0_wr[1296]),  .coef_in(coef[272]), .rdup_out(a1_wr[272]), .rdlo_out(a1_wr[1296]));
			radix2 #(.width(width)) rd_st0_273  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[273]), .rdlo_in(a0_wr[1297]),  .coef_in(coef[273]), .rdup_out(a1_wr[273]), .rdlo_out(a1_wr[1297]));
			radix2 #(.width(width)) rd_st0_274  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[274]), .rdlo_in(a0_wr[1298]),  .coef_in(coef[274]), .rdup_out(a1_wr[274]), .rdlo_out(a1_wr[1298]));
			radix2 #(.width(width)) rd_st0_275  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[275]), .rdlo_in(a0_wr[1299]),  .coef_in(coef[275]), .rdup_out(a1_wr[275]), .rdlo_out(a1_wr[1299]));
			radix2 #(.width(width)) rd_st0_276  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[276]), .rdlo_in(a0_wr[1300]),  .coef_in(coef[276]), .rdup_out(a1_wr[276]), .rdlo_out(a1_wr[1300]));
			radix2 #(.width(width)) rd_st0_277  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[277]), .rdlo_in(a0_wr[1301]),  .coef_in(coef[277]), .rdup_out(a1_wr[277]), .rdlo_out(a1_wr[1301]));
			radix2 #(.width(width)) rd_st0_278  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[278]), .rdlo_in(a0_wr[1302]),  .coef_in(coef[278]), .rdup_out(a1_wr[278]), .rdlo_out(a1_wr[1302]));
			radix2 #(.width(width)) rd_st0_279  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[279]), .rdlo_in(a0_wr[1303]),  .coef_in(coef[279]), .rdup_out(a1_wr[279]), .rdlo_out(a1_wr[1303]));
			radix2 #(.width(width)) rd_st0_280  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[280]), .rdlo_in(a0_wr[1304]),  .coef_in(coef[280]), .rdup_out(a1_wr[280]), .rdlo_out(a1_wr[1304]));
			radix2 #(.width(width)) rd_st0_281  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[281]), .rdlo_in(a0_wr[1305]),  .coef_in(coef[281]), .rdup_out(a1_wr[281]), .rdlo_out(a1_wr[1305]));
			radix2 #(.width(width)) rd_st0_282  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[282]), .rdlo_in(a0_wr[1306]),  .coef_in(coef[282]), .rdup_out(a1_wr[282]), .rdlo_out(a1_wr[1306]));
			radix2 #(.width(width)) rd_st0_283  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[283]), .rdlo_in(a0_wr[1307]),  .coef_in(coef[283]), .rdup_out(a1_wr[283]), .rdlo_out(a1_wr[1307]));
			radix2 #(.width(width)) rd_st0_284  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[284]), .rdlo_in(a0_wr[1308]),  .coef_in(coef[284]), .rdup_out(a1_wr[284]), .rdlo_out(a1_wr[1308]));
			radix2 #(.width(width)) rd_st0_285  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[285]), .rdlo_in(a0_wr[1309]),  .coef_in(coef[285]), .rdup_out(a1_wr[285]), .rdlo_out(a1_wr[1309]));
			radix2 #(.width(width)) rd_st0_286  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[286]), .rdlo_in(a0_wr[1310]),  .coef_in(coef[286]), .rdup_out(a1_wr[286]), .rdlo_out(a1_wr[1310]));
			radix2 #(.width(width)) rd_st0_287  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[287]), .rdlo_in(a0_wr[1311]),  .coef_in(coef[287]), .rdup_out(a1_wr[287]), .rdlo_out(a1_wr[1311]));
			radix2 #(.width(width)) rd_st0_288  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[288]), .rdlo_in(a0_wr[1312]),  .coef_in(coef[288]), .rdup_out(a1_wr[288]), .rdlo_out(a1_wr[1312]));
			radix2 #(.width(width)) rd_st0_289  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[289]), .rdlo_in(a0_wr[1313]),  .coef_in(coef[289]), .rdup_out(a1_wr[289]), .rdlo_out(a1_wr[1313]));
			radix2 #(.width(width)) rd_st0_290  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[290]), .rdlo_in(a0_wr[1314]),  .coef_in(coef[290]), .rdup_out(a1_wr[290]), .rdlo_out(a1_wr[1314]));
			radix2 #(.width(width)) rd_st0_291  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[291]), .rdlo_in(a0_wr[1315]),  .coef_in(coef[291]), .rdup_out(a1_wr[291]), .rdlo_out(a1_wr[1315]));
			radix2 #(.width(width)) rd_st0_292  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[292]), .rdlo_in(a0_wr[1316]),  .coef_in(coef[292]), .rdup_out(a1_wr[292]), .rdlo_out(a1_wr[1316]));
			radix2 #(.width(width)) rd_st0_293  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[293]), .rdlo_in(a0_wr[1317]),  .coef_in(coef[293]), .rdup_out(a1_wr[293]), .rdlo_out(a1_wr[1317]));
			radix2 #(.width(width)) rd_st0_294  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[294]), .rdlo_in(a0_wr[1318]),  .coef_in(coef[294]), .rdup_out(a1_wr[294]), .rdlo_out(a1_wr[1318]));
			radix2 #(.width(width)) rd_st0_295  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[295]), .rdlo_in(a0_wr[1319]),  .coef_in(coef[295]), .rdup_out(a1_wr[295]), .rdlo_out(a1_wr[1319]));
			radix2 #(.width(width)) rd_st0_296  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[296]), .rdlo_in(a0_wr[1320]),  .coef_in(coef[296]), .rdup_out(a1_wr[296]), .rdlo_out(a1_wr[1320]));
			radix2 #(.width(width)) rd_st0_297  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[297]), .rdlo_in(a0_wr[1321]),  .coef_in(coef[297]), .rdup_out(a1_wr[297]), .rdlo_out(a1_wr[1321]));
			radix2 #(.width(width)) rd_st0_298  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[298]), .rdlo_in(a0_wr[1322]),  .coef_in(coef[298]), .rdup_out(a1_wr[298]), .rdlo_out(a1_wr[1322]));
			radix2 #(.width(width)) rd_st0_299  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[299]), .rdlo_in(a0_wr[1323]),  .coef_in(coef[299]), .rdup_out(a1_wr[299]), .rdlo_out(a1_wr[1323]));
			radix2 #(.width(width)) rd_st0_300  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[300]), .rdlo_in(a0_wr[1324]),  .coef_in(coef[300]), .rdup_out(a1_wr[300]), .rdlo_out(a1_wr[1324]));
			radix2 #(.width(width)) rd_st0_301  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[301]), .rdlo_in(a0_wr[1325]),  .coef_in(coef[301]), .rdup_out(a1_wr[301]), .rdlo_out(a1_wr[1325]));
			radix2 #(.width(width)) rd_st0_302  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[302]), .rdlo_in(a0_wr[1326]),  .coef_in(coef[302]), .rdup_out(a1_wr[302]), .rdlo_out(a1_wr[1326]));
			radix2 #(.width(width)) rd_st0_303  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[303]), .rdlo_in(a0_wr[1327]),  .coef_in(coef[303]), .rdup_out(a1_wr[303]), .rdlo_out(a1_wr[1327]));
			radix2 #(.width(width)) rd_st0_304  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[304]), .rdlo_in(a0_wr[1328]),  .coef_in(coef[304]), .rdup_out(a1_wr[304]), .rdlo_out(a1_wr[1328]));
			radix2 #(.width(width)) rd_st0_305  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[305]), .rdlo_in(a0_wr[1329]),  .coef_in(coef[305]), .rdup_out(a1_wr[305]), .rdlo_out(a1_wr[1329]));
			radix2 #(.width(width)) rd_st0_306  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[306]), .rdlo_in(a0_wr[1330]),  .coef_in(coef[306]), .rdup_out(a1_wr[306]), .rdlo_out(a1_wr[1330]));
			radix2 #(.width(width)) rd_st0_307  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[307]), .rdlo_in(a0_wr[1331]),  .coef_in(coef[307]), .rdup_out(a1_wr[307]), .rdlo_out(a1_wr[1331]));
			radix2 #(.width(width)) rd_st0_308  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[308]), .rdlo_in(a0_wr[1332]),  .coef_in(coef[308]), .rdup_out(a1_wr[308]), .rdlo_out(a1_wr[1332]));
			radix2 #(.width(width)) rd_st0_309  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[309]), .rdlo_in(a0_wr[1333]),  .coef_in(coef[309]), .rdup_out(a1_wr[309]), .rdlo_out(a1_wr[1333]));
			radix2 #(.width(width)) rd_st0_310  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[310]), .rdlo_in(a0_wr[1334]),  .coef_in(coef[310]), .rdup_out(a1_wr[310]), .rdlo_out(a1_wr[1334]));
			radix2 #(.width(width)) rd_st0_311  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[311]), .rdlo_in(a0_wr[1335]),  .coef_in(coef[311]), .rdup_out(a1_wr[311]), .rdlo_out(a1_wr[1335]));
			radix2 #(.width(width)) rd_st0_312  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[312]), .rdlo_in(a0_wr[1336]),  .coef_in(coef[312]), .rdup_out(a1_wr[312]), .rdlo_out(a1_wr[1336]));
			radix2 #(.width(width)) rd_st0_313  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[313]), .rdlo_in(a0_wr[1337]),  .coef_in(coef[313]), .rdup_out(a1_wr[313]), .rdlo_out(a1_wr[1337]));
			radix2 #(.width(width)) rd_st0_314  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[314]), .rdlo_in(a0_wr[1338]),  .coef_in(coef[314]), .rdup_out(a1_wr[314]), .rdlo_out(a1_wr[1338]));
			radix2 #(.width(width)) rd_st0_315  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[315]), .rdlo_in(a0_wr[1339]),  .coef_in(coef[315]), .rdup_out(a1_wr[315]), .rdlo_out(a1_wr[1339]));
			radix2 #(.width(width)) rd_st0_316  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[316]), .rdlo_in(a0_wr[1340]),  .coef_in(coef[316]), .rdup_out(a1_wr[316]), .rdlo_out(a1_wr[1340]));
			radix2 #(.width(width)) rd_st0_317  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[317]), .rdlo_in(a0_wr[1341]),  .coef_in(coef[317]), .rdup_out(a1_wr[317]), .rdlo_out(a1_wr[1341]));
			radix2 #(.width(width)) rd_st0_318  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[318]), .rdlo_in(a0_wr[1342]),  .coef_in(coef[318]), .rdup_out(a1_wr[318]), .rdlo_out(a1_wr[1342]));
			radix2 #(.width(width)) rd_st0_319  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[319]), .rdlo_in(a0_wr[1343]),  .coef_in(coef[319]), .rdup_out(a1_wr[319]), .rdlo_out(a1_wr[1343]));
			radix2 #(.width(width)) rd_st0_320  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[320]), .rdlo_in(a0_wr[1344]),  .coef_in(coef[320]), .rdup_out(a1_wr[320]), .rdlo_out(a1_wr[1344]));
			radix2 #(.width(width)) rd_st0_321  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[321]), .rdlo_in(a0_wr[1345]),  .coef_in(coef[321]), .rdup_out(a1_wr[321]), .rdlo_out(a1_wr[1345]));
			radix2 #(.width(width)) rd_st0_322  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[322]), .rdlo_in(a0_wr[1346]),  .coef_in(coef[322]), .rdup_out(a1_wr[322]), .rdlo_out(a1_wr[1346]));
			radix2 #(.width(width)) rd_st0_323  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[323]), .rdlo_in(a0_wr[1347]),  .coef_in(coef[323]), .rdup_out(a1_wr[323]), .rdlo_out(a1_wr[1347]));
			radix2 #(.width(width)) rd_st0_324  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[324]), .rdlo_in(a0_wr[1348]),  .coef_in(coef[324]), .rdup_out(a1_wr[324]), .rdlo_out(a1_wr[1348]));
			radix2 #(.width(width)) rd_st0_325  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[325]), .rdlo_in(a0_wr[1349]),  .coef_in(coef[325]), .rdup_out(a1_wr[325]), .rdlo_out(a1_wr[1349]));
			radix2 #(.width(width)) rd_st0_326  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[326]), .rdlo_in(a0_wr[1350]),  .coef_in(coef[326]), .rdup_out(a1_wr[326]), .rdlo_out(a1_wr[1350]));
			radix2 #(.width(width)) rd_st0_327  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[327]), .rdlo_in(a0_wr[1351]),  .coef_in(coef[327]), .rdup_out(a1_wr[327]), .rdlo_out(a1_wr[1351]));
			radix2 #(.width(width)) rd_st0_328  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[328]), .rdlo_in(a0_wr[1352]),  .coef_in(coef[328]), .rdup_out(a1_wr[328]), .rdlo_out(a1_wr[1352]));
			radix2 #(.width(width)) rd_st0_329  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[329]), .rdlo_in(a0_wr[1353]),  .coef_in(coef[329]), .rdup_out(a1_wr[329]), .rdlo_out(a1_wr[1353]));
			radix2 #(.width(width)) rd_st0_330  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[330]), .rdlo_in(a0_wr[1354]),  .coef_in(coef[330]), .rdup_out(a1_wr[330]), .rdlo_out(a1_wr[1354]));
			radix2 #(.width(width)) rd_st0_331  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[331]), .rdlo_in(a0_wr[1355]),  .coef_in(coef[331]), .rdup_out(a1_wr[331]), .rdlo_out(a1_wr[1355]));
			radix2 #(.width(width)) rd_st0_332  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[332]), .rdlo_in(a0_wr[1356]),  .coef_in(coef[332]), .rdup_out(a1_wr[332]), .rdlo_out(a1_wr[1356]));
			radix2 #(.width(width)) rd_st0_333  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[333]), .rdlo_in(a0_wr[1357]),  .coef_in(coef[333]), .rdup_out(a1_wr[333]), .rdlo_out(a1_wr[1357]));
			radix2 #(.width(width)) rd_st0_334  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[334]), .rdlo_in(a0_wr[1358]),  .coef_in(coef[334]), .rdup_out(a1_wr[334]), .rdlo_out(a1_wr[1358]));
			radix2 #(.width(width)) rd_st0_335  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[335]), .rdlo_in(a0_wr[1359]),  .coef_in(coef[335]), .rdup_out(a1_wr[335]), .rdlo_out(a1_wr[1359]));
			radix2 #(.width(width)) rd_st0_336  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[336]), .rdlo_in(a0_wr[1360]),  .coef_in(coef[336]), .rdup_out(a1_wr[336]), .rdlo_out(a1_wr[1360]));
			radix2 #(.width(width)) rd_st0_337  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[337]), .rdlo_in(a0_wr[1361]),  .coef_in(coef[337]), .rdup_out(a1_wr[337]), .rdlo_out(a1_wr[1361]));
			radix2 #(.width(width)) rd_st0_338  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[338]), .rdlo_in(a0_wr[1362]),  .coef_in(coef[338]), .rdup_out(a1_wr[338]), .rdlo_out(a1_wr[1362]));
			radix2 #(.width(width)) rd_st0_339  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[339]), .rdlo_in(a0_wr[1363]),  .coef_in(coef[339]), .rdup_out(a1_wr[339]), .rdlo_out(a1_wr[1363]));
			radix2 #(.width(width)) rd_st0_340  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[340]), .rdlo_in(a0_wr[1364]),  .coef_in(coef[340]), .rdup_out(a1_wr[340]), .rdlo_out(a1_wr[1364]));
			radix2 #(.width(width)) rd_st0_341  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[341]), .rdlo_in(a0_wr[1365]),  .coef_in(coef[341]), .rdup_out(a1_wr[341]), .rdlo_out(a1_wr[1365]));
			radix2 #(.width(width)) rd_st0_342  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[342]), .rdlo_in(a0_wr[1366]),  .coef_in(coef[342]), .rdup_out(a1_wr[342]), .rdlo_out(a1_wr[1366]));
			radix2 #(.width(width)) rd_st0_343  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[343]), .rdlo_in(a0_wr[1367]),  .coef_in(coef[343]), .rdup_out(a1_wr[343]), .rdlo_out(a1_wr[1367]));
			radix2 #(.width(width)) rd_st0_344  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[344]), .rdlo_in(a0_wr[1368]),  .coef_in(coef[344]), .rdup_out(a1_wr[344]), .rdlo_out(a1_wr[1368]));
			radix2 #(.width(width)) rd_st0_345  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[345]), .rdlo_in(a0_wr[1369]),  .coef_in(coef[345]), .rdup_out(a1_wr[345]), .rdlo_out(a1_wr[1369]));
			radix2 #(.width(width)) rd_st0_346  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[346]), .rdlo_in(a0_wr[1370]),  .coef_in(coef[346]), .rdup_out(a1_wr[346]), .rdlo_out(a1_wr[1370]));
			radix2 #(.width(width)) rd_st0_347  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[347]), .rdlo_in(a0_wr[1371]),  .coef_in(coef[347]), .rdup_out(a1_wr[347]), .rdlo_out(a1_wr[1371]));
			radix2 #(.width(width)) rd_st0_348  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[348]), .rdlo_in(a0_wr[1372]),  .coef_in(coef[348]), .rdup_out(a1_wr[348]), .rdlo_out(a1_wr[1372]));
			radix2 #(.width(width)) rd_st0_349  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[349]), .rdlo_in(a0_wr[1373]),  .coef_in(coef[349]), .rdup_out(a1_wr[349]), .rdlo_out(a1_wr[1373]));
			radix2 #(.width(width)) rd_st0_350  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[350]), .rdlo_in(a0_wr[1374]),  .coef_in(coef[350]), .rdup_out(a1_wr[350]), .rdlo_out(a1_wr[1374]));
			radix2 #(.width(width)) rd_st0_351  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[351]), .rdlo_in(a0_wr[1375]),  .coef_in(coef[351]), .rdup_out(a1_wr[351]), .rdlo_out(a1_wr[1375]));
			radix2 #(.width(width)) rd_st0_352  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[352]), .rdlo_in(a0_wr[1376]),  .coef_in(coef[352]), .rdup_out(a1_wr[352]), .rdlo_out(a1_wr[1376]));
			radix2 #(.width(width)) rd_st0_353  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[353]), .rdlo_in(a0_wr[1377]),  .coef_in(coef[353]), .rdup_out(a1_wr[353]), .rdlo_out(a1_wr[1377]));
			radix2 #(.width(width)) rd_st0_354  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[354]), .rdlo_in(a0_wr[1378]),  .coef_in(coef[354]), .rdup_out(a1_wr[354]), .rdlo_out(a1_wr[1378]));
			radix2 #(.width(width)) rd_st0_355  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[355]), .rdlo_in(a0_wr[1379]),  .coef_in(coef[355]), .rdup_out(a1_wr[355]), .rdlo_out(a1_wr[1379]));
			radix2 #(.width(width)) rd_st0_356  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[356]), .rdlo_in(a0_wr[1380]),  .coef_in(coef[356]), .rdup_out(a1_wr[356]), .rdlo_out(a1_wr[1380]));
			radix2 #(.width(width)) rd_st0_357  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[357]), .rdlo_in(a0_wr[1381]),  .coef_in(coef[357]), .rdup_out(a1_wr[357]), .rdlo_out(a1_wr[1381]));
			radix2 #(.width(width)) rd_st0_358  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[358]), .rdlo_in(a0_wr[1382]),  .coef_in(coef[358]), .rdup_out(a1_wr[358]), .rdlo_out(a1_wr[1382]));
			radix2 #(.width(width)) rd_st0_359  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[359]), .rdlo_in(a0_wr[1383]),  .coef_in(coef[359]), .rdup_out(a1_wr[359]), .rdlo_out(a1_wr[1383]));
			radix2 #(.width(width)) rd_st0_360  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[360]), .rdlo_in(a0_wr[1384]),  .coef_in(coef[360]), .rdup_out(a1_wr[360]), .rdlo_out(a1_wr[1384]));
			radix2 #(.width(width)) rd_st0_361  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[361]), .rdlo_in(a0_wr[1385]),  .coef_in(coef[361]), .rdup_out(a1_wr[361]), .rdlo_out(a1_wr[1385]));
			radix2 #(.width(width)) rd_st0_362  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[362]), .rdlo_in(a0_wr[1386]),  .coef_in(coef[362]), .rdup_out(a1_wr[362]), .rdlo_out(a1_wr[1386]));
			radix2 #(.width(width)) rd_st0_363  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[363]), .rdlo_in(a0_wr[1387]),  .coef_in(coef[363]), .rdup_out(a1_wr[363]), .rdlo_out(a1_wr[1387]));
			radix2 #(.width(width)) rd_st0_364  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[364]), .rdlo_in(a0_wr[1388]),  .coef_in(coef[364]), .rdup_out(a1_wr[364]), .rdlo_out(a1_wr[1388]));
			radix2 #(.width(width)) rd_st0_365  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[365]), .rdlo_in(a0_wr[1389]),  .coef_in(coef[365]), .rdup_out(a1_wr[365]), .rdlo_out(a1_wr[1389]));
			radix2 #(.width(width)) rd_st0_366  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[366]), .rdlo_in(a0_wr[1390]),  .coef_in(coef[366]), .rdup_out(a1_wr[366]), .rdlo_out(a1_wr[1390]));
			radix2 #(.width(width)) rd_st0_367  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[367]), .rdlo_in(a0_wr[1391]),  .coef_in(coef[367]), .rdup_out(a1_wr[367]), .rdlo_out(a1_wr[1391]));
			radix2 #(.width(width)) rd_st0_368  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[368]), .rdlo_in(a0_wr[1392]),  .coef_in(coef[368]), .rdup_out(a1_wr[368]), .rdlo_out(a1_wr[1392]));
			radix2 #(.width(width)) rd_st0_369  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[369]), .rdlo_in(a0_wr[1393]),  .coef_in(coef[369]), .rdup_out(a1_wr[369]), .rdlo_out(a1_wr[1393]));
			radix2 #(.width(width)) rd_st0_370  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[370]), .rdlo_in(a0_wr[1394]),  .coef_in(coef[370]), .rdup_out(a1_wr[370]), .rdlo_out(a1_wr[1394]));
			radix2 #(.width(width)) rd_st0_371  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[371]), .rdlo_in(a0_wr[1395]),  .coef_in(coef[371]), .rdup_out(a1_wr[371]), .rdlo_out(a1_wr[1395]));
			radix2 #(.width(width)) rd_st0_372  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[372]), .rdlo_in(a0_wr[1396]),  .coef_in(coef[372]), .rdup_out(a1_wr[372]), .rdlo_out(a1_wr[1396]));
			radix2 #(.width(width)) rd_st0_373  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[373]), .rdlo_in(a0_wr[1397]),  .coef_in(coef[373]), .rdup_out(a1_wr[373]), .rdlo_out(a1_wr[1397]));
			radix2 #(.width(width)) rd_st0_374  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[374]), .rdlo_in(a0_wr[1398]),  .coef_in(coef[374]), .rdup_out(a1_wr[374]), .rdlo_out(a1_wr[1398]));
			radix2 #(.width(width)) rd_st0_375  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[375]), .rdlo_in(a0_wr[1399]),  .coef_in(coef[375]), .rdup_out(a1_wr[375]), .rdlo_out(a1_wr[1399]));
			radix2 #(.width(width)) rd_st0_376  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[376]), .rdlo_in(a0_wr[1400]),  .coef_in(coef[376]), .rdup_out(a1_wr[376]), .rdlo_out(a1_wr[1400]));
			radix2 #(.width(width)) rd_st0_377  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[377]), .rdlo_in(a0_wr[1401]),  .coef_in(coef[377]), .rdup_out(a1_wr[377]), .rdlo_out(a1_wr[1401]));
			radix2 #(.width(width)) rd_st0_378  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[378]), .rdlo_in(a0_wr[1402]),  .coef_in(coef[378]), .rdup_out(a1_wr[378]), .rdlo_out(a1_wr[1402]));
			radix2 #(.width(width)) rd_st0_379  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[379]), .rdlo_in(a0_wr[1403]),  .coef_in(coef[379]), .rdup_out(a1_wr[379]), .rdlo_out(a1_wr[1403]));
			radix2 #(.width(width)) rd_st0_380  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[380]), .rdlo_in(a0_wr[1404]),  .coef_in(coef[380]), .rdup_out(a1_wr[380]), .rdlo_out(a1_wr[1404]));
			radix2 #(.width(width)) rd_st0_381  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[381]), .rdlo_in(a0_wr[1405]),  .coef_in(coef[381]), .rdup_out(a1_wr[381]), .rdlo_out(a1_wr[1405]));
			radix2 #(.width(width)) rd_st0_382  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[382]), .rdlo_in(a0_wr[1406]),  .coef_in(coef[382]), .rdup_out(a1_wr[382]), .rdlo_out(a1_wr[1406]));
			radix2 #(.width(width)) rd_st0_383  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[383]), .rdlo_in(a0_wr[1407]),  .coef_in(coef[383]), .rdup_out(a1_wr[383]), .rdlo_out(a1_wr[1407]));
			radix2 #(.width(width)) rd_st0_384  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[384]), .rdlo_in(a0_wr[1408]),  .coef_in(coef[384]), .rdup_out(a1_wr[384]), .rdlo_out(a1_wr[1408]));
			radix2 #(.width(width)) rd_st0_385  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[385]), .rdlo_in(a0_wr[1409]),  .coef_in(coef[385]), .rdup_out(a1_wr[385]), .rdlo_out(a1_wr[1409]));
			radix2 #(.width(width)) rd_st0_386  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[386]), .rdlo_in(a0_wr[1410]),  .coef_in(coef[386]), .rdup_out(a1_wr[386]), .rdlo_out(a1_wr[1410]));
			radix2 #(.width(width)) rd_st0_387  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[387]), .rdlo_in(a0_wr[1411]),  .coef_in(coef[387]), .rdup_out(a1_wr[387]), .rdlo_out(a1_wr[1411]));
			radix2 #(.width(width)) rd_st0_388  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[388]), .rdlo_in(a0_wr[1412]),  .coef_in(coef[388]), .rdup_out(a1_wr[388]), .rdlo_out(a1_wr[1412]));
			radix2 #(.width(width)) rd_st0_389  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[389]), .rdlo_in(a0_wr[1413]),  .coef_in(coef[389]), .rdup_out(a1_wr[389]), .rdlo_out(a1_wr[1413]));
			radix2 #(.width(width)) rd_st0_390  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[390]), .rdlo_in(a0_wr[1414]),  .coef_in(coef[390]), .rdup_out(a1_wr[390]), .rdlo_out(a1_wr[1414]));
			radix2 #(.width(width)) rd_st0_391  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[391]), .rdlo_in(a0_wr[1415]),  .coef_in(coef[391]), .rdup_out(a1_wr[391]), .rdlo_out(a1_wr[1415]));
			radix2 #(.width(width)) rd_st0_392  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[392]), .rdlo_in(a0_wr[1416]),  .coef_in(coef[392]), .rdup_out(a1_wr[392]), .rdlo_out(a1_wr[1416]));
			radix2 #(.width(width)) rd_st0_393  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[393]), .rdlo_in(a0_wr[1417]),  .coef_in(coef[393]), .rdup_out(a1_wr[393]), .rdlo_out(a1_wr[1417]));
			radix2 #(.width(width)) rd_st0_394  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[394]), .rdlo_in(a0_wr[1418]),  .coef_in(coef[394]), .rdup_out(a1_wr[394]), .rdlo_out(a1_wr[1418]));
			radix2 #(.width(width)) rd_st0_395  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[395]), .rdlo_in(a0_wr[1419]),  .coef_in(coef[395]), .rdup_out(a1_wr[395]), .rdlo_out(a1_wr[1419]));
			radix2 #(.width(width)) rd_st0_396  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[396]), .rdlo_in(a0_wr[1420]),  .coef_in(coef[396]), .rdup_out(a1_wr[396]), .rdlo_out(a1_wr[1420]));
			radix2 #(.width(width)) rd_st0_397  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[397]), .rdlo_in(a0_wr[1421]),  .coef_in(coef[397]), .rdup_out(a1_wr[397]), .rdlo_out(a1_wr[1421]));
			radix2 #(.width(width)) rd_st0_398  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[398]), .rdlo_in(a0_wr[1422]),  .coef_in(coef[398]), .rdup_out(a1_wr[398]), .rdlo_out(a1_wr[1422]));
			radix2 #(.width(width)) rd_st0_399  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[399]), .rdlo_in(a0_wr[1423]),  .coef_in(coef[399]), .rdup_out(a1_wr[399]), .rdlo_out(a1_wr[1423]));
			radix2 #(.width(width)) rd_st0_400  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[400]), .rdlo_in(a0_wr[1424]),  .coef_in(coef[400]), .rdup_out(a1_wr[400]), .rdlo_out(a1_wr[1424]));
			radix2 #(.width(width)) rd_st0_401  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[401]), .rdlo_in(a0_wr[1425]),  .coef_in(coef[401]), .rdup_out(a1_wr[401]), .rdlo_out(a1_wr[1425]));
			radix2 #(.width(width)) rd_st0_402  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[402]), .rdlo_in(a0_wr[1426]),  .coef_in(coef[402]), .rdup_out(a1_wr[402]), .rdlo_out(a1_wr[1426]));
			radix2 #(.width(width)) rd_st0_403  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[403]), .rdlo_in(a0_wr[1427]),  .coef_in(coef[403]), .rdup_out(a1_wr[403]), .rdlo_out(a1_wr[1427]));
			radix2 #(.width(width)) rd_st0_404  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[404]), .rdlo_in(a0_wr[1428]),  .coef_in(coef[404]), .rdup_out(a1_wr[404]), .rdlo_out(a1_wr[1428]));
			radix2 #(.width(width)) rd_st0_405  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[405]), .rdlo_in(a0_wr[1429]),  .coef_in(coef[405]), .rdup_out(a1_wr[405]), .rdlo_out(a1_wr[1429]));
			radix2 #(.width(width)) rd_st0_406  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[406]), .rdlo_in(a0_wr[1430]),  .coef_in(coef[406]), .rdup_out(a1_wr[406]), .rdlo_out(a1_wr[1430]));
			radix2 #(.width(width)) rd_st0_407  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[407]), .rdlo_in(a0_wr[1431]),  .coef_in(coef[407]), .rdup_out(a1_wr[407]), .rdlo_out(a1_wr[1431]));
			radix2 #(.width(width)) rd_st0_408  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[408]), .rdlo_in(a0_wr[1432]),  .coef_in(coef[408]), .rdup_out(a1_wr[408]), .rdlo_out(a1_wr[1432]));
			radix2 #(.width(width)) rd_st0_409  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[409]), .rdlo_in(a0_wr[1433]),  .coef_in(coef[409]), .rdup_out(a1_wr[409]), .rdlo_out(a1_wr[1433]));
			radix2 #(.width(width)) rd_st0_410  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[410]), .rdlo_in(a0_wr[1434]),  .coef_in(coef[410]), .rdup_out(a1_wr[410]), .rdlo_out(a1_wr[1434]));
			radix2 #(.width(width)) rd_st0_411  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[411]), .rdlo_in(a0_wr[1435]),  .coef_in(coef[411]), .rdup_out(a1_wr[411]), .rdlo_out(a1_wr[1435]));
			radix2 #(.width(width)) rd_st0_412  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[412]), .rdlo_in(a0_wr[1436]),  .coef_in(coef[412]), .rdup_out(a1_wr[412]), .rdlo_out(a1_wr[1436]));
			radix2 #(.width(width)) rd_st0_413  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[413]), .rdlo_in(a0_wr[1437]),  .coef_in(coef[413]), .rdup_out(a1_wr[413]), .rdlo_out(a1_wr[1437]));
			radix2 #(.width(width)) rd_st0_414  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[414]), .rdlo_in(a0_wr[1438]),  .coef_in(coef[414]), .rdup_out(a1_wr[414]), .rdlo_out(a1_wr[1438]));
			radix2 #(.width(width)) rd_st0_415  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[415]), .rdlo_in(a0_wr[1439]),  .coef_in(coef[415]), .rdup_out(a1_wr[415]), .rdlo_out(a1_wr[1439]));
			radix2 #(.width(width)) rd_st0_416  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[416]), .rdlo_in(a0_wr[1440]),  .coef_in(coef[416]), .rdup_out(a1_wr[416]), .rdlo_out(a1_wr[1440]));
			radix2 #(.width(width)) rd_st0_417  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[417]), .rdlo_in(a0_wr[1441]),  .coef_in(coef[417]), .rdup_out(a1_wr[417]), .rdlo_out(a1_wr[1441]));
			radix2 #(.width(width)) rd_st0_418  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[418]), .rdlo_in(a0_wr[1442]),  .coef_in(coef[418]), .rdup_out(a1_wr[418]), .rdlo_out(a1_wr[1442]));
			radix2 #(.width(width)) rd_st0_419  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[419]), .rdlo_in(a0_wr[1443]),  .coef_in(coef[419]), .rdup_out(a1_wr[419]), .rdlo_out(a1_wr[1443]));
			radix2 #(.width(width)) rd_st0_420  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[420]), .rdlo_in(a0_wr[1444]),  .coef_in(coef[420]), .rdup_out(a1_wr[420]), .rdlo_out(a1_wr[1444]));
			radix2 #(.width(width)) rd_st0_421  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[421]), .rdlo_in(a0_wr[1445]),  .coef_in(coef[421]), .rdup_out(a1_wr[421]), .rdlo_out(a1_wr[1445]));
			radix2 #(.width(width)) rd_st0_422  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[422]), .rdlo_in(a0_wr[1446]),  .coef_in(coef[422]), .rdup_out(a1_wr[422]), .rdlo_out(a1_wr[1446]));
			radix2 #(.width(width)) rd_st0_423  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[423]), .rdlo_in(a0_wr[1447]),  .coef_in(coef[423]), .rdup_out(a1_wr[423]), .rdlo_out(a1_wr[1447]));
			radix2 #(.width(width)) rd_st0_424  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[424]), .rdlo_in(a0_wr[1448]),  .coef_in(coef[424]), .rdup_out(a1_wr[424]), .rdlo_out(a1_wr[1448]));
			radix2 #(.width(width)) rd_st0_425  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[425]), .rdlo_in(a0_wr[1449]),  .coef_in(coef[425]), .rdup_out(a1_wr[425]), .rdlo_out(a1_wr[1449]));
			radix2 #(.width(width)) rd_st0_426  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[426]), .rdlo_in(a0_wr[1450]),  .coef_in(coef[426]), .rdup_out(a1_wr[426]), .rdlo_out(a1_wr[1450]));
			radix2 #(.width(width)) rd_st0_427  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[427]), .rdlo_in(a0_wr[1451]),  .coef_in(coef[427]), .rdup_out(a1_wr[427]), .rdlo_out(a1_wr[1451]));
			radix2 #(.width(width)) rd_st0_428  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[428]), .rdlo_in(a0_wr[1452]),  .coef_in(coef[428]), .rdup_out(a1_wr[428]), .rdlo_out(a1_wr[1452]));
			radix2 #(.width(width)) rd_st0_429  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[429]), .rdlo_in(a0_wr[1453]),  .coef_in(coef[429]), .rdup_out(a1_wr[429]), .rdlo_out(a1_wr[1453]));
			radix2 #(.width(width)) rd_st0_430  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[430]), .rdlo_in(a0_wr[1454]),  .coef_in(coef[430]), .rdup_out(a1_wr[430]), .rdlo_out(a1_wr[1454]));
			radix2 #(.width(width)) rd_st0_431  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[431]), .rdlo_in(a0_wr[1455]),  .coef_in(coef[431]), .rdup_out(a1_wr[431]), .rdlo_out(a1_wr[1455]));
			radix2 #(.width(width)) rd_st0_432  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[432]), .rdlo_in(a0_wr[1456]),  .coef_in(coef[432]), .rdup_out(a1_wr[432]), .rdlo_out(a1_wr[1456]));
			radix2 #(.width(width)) rd_st0_433  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[433]), .rdlo_in(a0_wr[1457]),  .coef_in(coef[433]), .rdup_out(a1_wr[433]), .rdlo_out(a1_wr[1457]));
			radix2 #(.width(width)) rd_st0_434  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[434]), .rdlo_in(a0_wr[1458]),  .coef_in(coef[434]), .rdup_out(a1_wr[434]), .rdlo_out(a1_wr[1458]));
			radix2 #(.width(width)) rd_st0_435  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[435]), .rdlo_in(a0_wr[1459]),  .coef_in(coef[435]), .rdup_out(a1_wr[435]), .rdlo_out(a1_wr[1459]));
			radix2 #(.width(width)) rd_st0_436  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[436]), .rdlo_in(a0_wr[1460]),  .coef_in(coef[436]), .rdup_out(a1_wr[436]), .rdlo_out(a1_wr[1460]));
			radix2 #(.width(width)) rd_st0_437  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[437]), .rdlo_in(a0_wr[1461]),  .coef_in(coef[437]), .rdup_out(a1_wr[437]), .rdlo_out(a1_wr[1461]));
			radix2 #(.width(width)) rd_st0_438  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[438]), .rdlo_in(a0_wr[1462]),  .coef_in(coef[438]), .rdup_out(a1_wr[438]), .rdlo_out(a1_wr[1462]));
			radix2 #(.width(width)) rd_st0_439  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[439]), .rdlo_in(a0_wr[1463]),  .coef_in(coef[439]), .rdup_out(a1_wr[439]), .rdlo_out(a1_wr[1463]));
			radix2 #(.width(width)) rd_st0_440  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[440]), .rdlo_in(a0_wr[1464]),  .coef_in(coef[440]), .rdup_out(a1_wr[440]), .rdlo_out(a1_wr[1464]));
			radix2 #(.width(width)) rd_st0_441  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[441]), .rdlo_in(a0_wr[1465]),  .coef_in(coef[441]), .rdup_out(a1_wr[441]), .rdlo_out(a1_wr[1465]));
			radix2 #(.width(width)) rd_st0_442  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[442]), .rdlo_in(a0_wr[1466]),  .coef_in(coef[442]), .rdup_out(a1_wr[442]), .rdlo_out(a1_wr[1466]));
			radix2 #(.width(width)) rd_st0_443  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[443]), .rdlo_in(a0_wr[1467]),  .coef_in(coef[443]), .rdup_out(a1_wr[443]), .rdlo_out(a1_wr[1467]));
			radix2 #(.width(width)) rd_st0_444  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[444]), .rdlo_in(a0_wr[1468]),  .coef_in(coef[444]), .rdup_out(a1_wr[444]), .rdlo_out(a1_wr[1468]));
			radix2 #(.width(width)) rd_st0_445  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[445]), .rdlo_in(a0_wr[1469]),  .coef_in(coef[445]), .rdup_out(a1_wr[445]), .rdlo_out(a1_wr[1469]));
			radix2 #(.width(width)) rd_st0_446  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[446]), .rdlo_in(a0_wr[1470]),  .coef_in(coef[446]), .rdup_out(a1_wr[446]), .rdlo_out(a1_wr[1470]));
			radix2 #(.width(width)) rd_st0_447  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[447]), .rdlo_in(a0_wr[1471]),  .coef_in(coef[447]), .rdup_out(a1_wr[447]), .rdlo_out(a1_wr[1471]));
			radix2 #(.width(width)) rd_st0_448  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[448]), .rdlo_in(a0_wr[1472]),  .coef_in(coef[448]), .rdup_out(a1_wr[448]), .rdlo_out(a1_wr[1472]));
			radix2 #(.width(width)) rd_st0_449  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[449]), .rdlo_in(a0_wr[1473]),  .coef_in(coef[449]), .rdup_out(a1_wr[449]), .rdlo_out(a1_wr[1473]));
			radix2 #(.width(width)) rd_st0_450  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[450]), .rdlo_in(a0_wr[1474]),  .coef_in(coef[450]), .rdup_out(a1_wr[450]), .rdlo_out(a1_wr[1474]));
			radix2 #(.width(width)) rd_st0_451  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[451]), .rdlo_in(a0_wr[1475]),  .coef_in(coef[451]), .rdup_out(a1_wr[451]), .rdlo_out(a1_wr[1475]));
			radix2 #(.width(width)) rd_st0_452  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[452]), .rdlo_in(a0_wr[1476]),  .coef_in(coef[452]), .rdup_out(a1_wr[452]), .rdlo_out(a1_wr[1476]));
			radix2 #(.width(width)) rd_st0_453  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[453]), .rdlo_in(a0_wr[1477]),  .coef_in(coef[453]), .rdup_out(a1_wr[453]), .rdlo_out(a1_wr[1477]));
			radix2 #(.width(width)) rd_st0_454  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[454]), .rdlo_in(a0_wr[1478]),  .coef_in(coef[454]), .rdup_out(a1_wr[454]), .rdlo_out(a1_wr[1478]));
			radix2 #(.width(width)) rd_st0_455  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[455]), .rdlo_in(a0_wr[1479]),  .coef_in(coef[455]), .rdup_out(a1_wr[455]), .rdlo_out(a1_wr[1479]));
			radix2 #(.width(width)) rd_st0_456  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[456]), .rdlo_in(a0_wr[1480]),  .coef_in(coef[456]), .rdup_out(a1_wr[456]), .rdlo_out(a1_wr[1480]));
			radix2 #(.width(width)) rd_st0_457  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[457]), .rdlo_in(a0_wr[1481]),  .coef_in(coef[457]), .rdup_out(a1_wr[457]), .rdlo_out(a1_wr[1481]));
			radix2 #(.width(width)) rd_st0_458  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[458]), .rdlo_in(a0_wr[1482]),  .coef_in(coef[458]), .rdup_out(a1_wr[458]), .rdlo_out(a1_wr[1482]));
			radix2 #(.width(width)) rd_st0_459  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[459]), .rdlo_in(a0_wr[1483]),  .coef_in(coef[459]), .rdup_out(a1_wr[459]), .rdlo_out(a1_wr[1483]));
			radix2 #(.width(width)) rd_st0_460  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[460]), .rdlo_in(a0_wr[1484]),  .coef_in(coef[460]), .rdup_out(a1_wr[460]), .rdlo_out(a1_wr[1484]));
			radix2 #(.width(width)) rd_st0_461  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[461]), .rdlo_in(a0_wr[1485]),  .coef_in(coef[461]), .rdup_out(a1_wr[461]), .rdlo_out(a1_wr[1485]));
			radix2 #(.width(width)) rd_st0_462  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[462]), .rdlo_in(a0_wr[1486]),  .coef_in(coef[462]), .rdup_out(a1_wr[462]), .rdlo_out(a1_wr[1486]));
			radix2 #(.width(width)) rd_st0_463  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[463]), .rdlo_in(a0_wr[1487]),  .coef_in(coef[463]), .rdup_out(a1_wr[463]), .rdlo_out(a1_wr[1487]));
			radix2 #(.width(width)) rd_st0_464  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[464]), .rdlo_in(a0_wr[1488]),  .coef_in(coef[464]), .rdup_out(a1_wr[464]), .rdlo_out(a1_wr[1488]));
			radix2 #(.width(width)) rd_st0_465  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[465]), .rdlo_in(a0_wr[1489]),  .coef_in(coef[465]), .rdup_out(a1_wr[465]), .rdlo_out(a1_wr[1489]));
			radix2 #(.width(width)) rd_st0_466  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[466]), .rdlo_in(a0_wr[1490]),  .coef_in(coef[466]), .rdup_out(a1_wr[466]), .rdlo_out(a1_wr[1490]));
			radix2 #(.width(width)) rd_st0_467  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[467]), .rdlo_in(a0_wr[1491]),  .coef_in(coef[467]), .rdup_out(a1_wr[467]), .rdlo_out(a1_wr[1491]));
			radix2 #(.width(width)) rd_st0_468  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[468]), .rdlo_in(a0_wr[1492]),  .coef_in(coef[468]), .rdup_out(a1_wr[468]), .rdlo_out(a1_wr[1492]));
			radix2 #(.width(width)) rd_st0_469  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[469]), .rdlo_in(a0_wr[1493]),  .coef_in(coef[469]), .rdup_out(a1_wr[469]), .rdlo_out(a1_wr[1493]));
			radix2 #(.width(width)) rd_st0_470  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[470]), .rdlo_in(a0_wr[1494]),  .coef_in(coef[470]), .rdup_out(a1_wr[470]), .rdlo_out(a1_wr[1494]));
			radix2 #(.width(width)) rd_st0_471  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[471]), .rdlo_in(a0_wr[1495]),  .coef_in(coef[471]), .rdup_out(a1_wr[471]), .rdlo_out(a1_wr[1495]));
			radix2 #(.width(width)) rd_st0_472  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[472]), .rdlo_in(a0_wr[1496]),  .coef_in(coef[472]), .rdup_out(a1_wr[472]), .rdlo_out(a1_wr[1496]));
			radix2 #(.width(width)) rd_st0_473  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[473]), .rdlo_in(a0_wr[1497]),  .coef_in(coef[473]), .rdup_out(a1_wr[473]), .rdlo_out(a1_wr[1497]));
			radix2 #(.width(width)) rd_st0_474  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[474]), .rdlo_in(a0_wr[1498]),  .coef_in(coef[474]), .rdup_out(a1_wr[474]), .rdlo_out(a1_wr[1498]));
			radix2 #(.width(width)) rd_st0_475  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[475]), .rdlo_in(a0_wr[1499]),  .coef_in(coef[475]), .rdup_out(a1_wr[475]), .rdlo_out(a1_wr[1499]));
			radix2 #(.width(width)) rd_st0_476  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[476]), .rdlo_in(a0_wr[1500]),  .coef_in(coef[476]), .rdup_out(a1_wr[476]), .rdlo_out(a1_wr[1500]));
			radix2 #(.width(width)) rd_st0_477  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[477]), .rdlo_in(a0_wr[1501]),  .coef_in(coef[477]), .rdup_out(a1_wr[477]), .rdlo_out(a1_wr[1501]));
			radix2 #(.width(width)) rd_st0_478  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[478]), .rdlo_in(a0_wr[1502]),  .coef_in(coef[478]), .rdup_out(a1_wr[478]), .rdlo_out(a1_wr[1502]));
			radix2 #(.width(width)) rd_st0_479  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[479]), .rdlo_in(a0_wr[1503]),  .coef_in(coef[479]), .rdup_out(a1_wr[479]), .rdlo_out(a1_wr[1503]));
			radix2 #(.width(width)) rd_st0_480  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[480]), .rdlo_in(a0_wr[1504]),  .coef_in(coef[480]), .rdup_out(a1_wr[480]), .rdlo_out(a1_wr[1504]));
			radix2 #(.width(width)) rd_st0_481  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[481]), .rdlo_in(a0_wr[1505]),  .coef_in(coef[481]), .rdup_out(a1_wr[481]), .rdlo_out(a1_wr[1505]));
			radix2 #(.width(width)) rd_st0_482  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[482]), .rdlo_in(a0_wr[1506]),  .coef_in(coef[482]), .rdup_out(a1_wr[482]), .rdlo_out(a1_wr[1506]));
			radix2 #(.width(width)) rd_st0_483  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[483]), .rdlo_in(a0_wr[1507]),  .coef_in(coef[483]), .rdup_out(a1_wr[483]), .rdlo_out(a1_wr[1507]));
			radix2 #(.width(width)) rd_st0_484  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[484]), .rdlo_in(a0_wr[1508]),  .coef_in(coef[484]), .rdup_out(a1_wr[484]), .rdlo_out(a1_wr[1508]));
			radix2 #(.width(width)) rd_st0_485  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[485]), .rdlo_in(a0_wr[1509]),  .coef_in(coef[485]), .rdup_out(a1_wr[485]), .rdlo_out(a1_wr[1509]));
			radix2 #(.width(width)) rd_st0_486  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[486]), .rdlo_in(a0_wr[1510]),  .coef_in(coef[486]), .rdup_out(a1_wr[486]), .rdlo_out(a1_wr[1510]));
			radix2 #(.width(width)) rd_st0_487  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[487]), .rdlo_in(a0_wr[1511]),  .coef_in(coef[487]), .rdup_out(a1_wr[487]), .rdlo_out(a1_wr[1511]));
			radix2 #(.width(width)) rd_st0_488  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[488]), .rdlo_in(a0_wr[1512]),  .coef_in(coef[488]), .rdup_out(a1_wr[488]), .rdlo_out(a1_wr[1512]));
			radix2 #(.width(width)) rd_st0_489  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[489]), .rdlo_in(a0_wr[1513]),  .coef_in(coef[489]), .rdup_out(a1_wr[489]), .rdlo_out(a1_wr[1513]));
			radix2 #(.width(width)) rd_st0_490  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[490]), .rdlo_in(a0_wr[1514]),  .coef_in(coef[490]), .rdup_out(a1_wr[490]), .rdlo_out(a1_wr[1514]));
			radix2 #(.width(width)) rd_st0_491  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[491]), .rdlo_in(a0_wr[1515]),  .coef_in(coef[491]), .rdup_out(a1_wr[491]), .rdlo_out(a1_wr[1515]));
			radix2 #(.width(width)) rd_st0_492  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[492]), .rdlo_in(a0_wr[1516]),  .coef_in(coef[492]), .rdup_out(a1_wr[492]), .rdlo_out(a1_wr[1516]));
			radix2 #(.width(width)) rd_st0_493  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[493]), .rdlo_in(a0_wr[1517]),  .coef_in(coef[493]), .rdup_out(a1_wr[493]), .rdlo_out(a1_wr[1517]));
			radix2 #(.width(width)) rd_st0_494  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[494]), .rdlo_in(a0_wr[1518]),  .coef_in(coef[494]), .rdup_out(a1_wr[494]), .rdlo_out(a1_wr[1518]));
			radix2 #(.width(width)) rd_st0_495  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[495]), .rdlo_in(a0_wr[1519]),  .coef_in(coef[495]), .rdup_out(a1_wr[495]), .rdlo_out(a1_wr[1519]));
			radix2 #(.width(width)) rd_st0_496  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[496]), .rdlo_in(a0_wr[1520]),  .coef_in(coef[496]), .rdup_out(a1_wr[496]), .rdlo_out(a1_wr[1520]));
			radix2 #(.width(width)) rd_st0_497  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[497]), .rdlo_in(a0_wr[1521]),  .coef_in(coef[497]), .rdup_out(a1_wr[497]), .rdlo_out(a1_wr[1521]));
			radix2 #(.width(width)) rd_st0_498  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[498]), .rdlo_in(a0_wr[1522]),  .coef_in(coef[498]), .rdup_out(a1_wr[498]), .rdlo_out(a1_wr[1522]));
			radix2 #(.width(width)) rd_st0_499  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[499]), .rdlo_in(a0_wr[1523]),  .coef_in(coef[499]), .rdup_out(a1_wr[499]), .rdlo_out(a1_wr[1523]));
			radix2 #(.width(width)) rd_st0_500  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[500]), .rdlo_in(a0_wr[1524]),  .coef_in(coef[500]), .rdup_out(a1_wr[500]), .rdlo_out(a1_wr[1524]));
			radix2 #(.width(width)) rd_st0_501  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[501]), .rdlo_in(a0_wr[1525]),  .coef_in(coef[501]), .rdup_out(a1_wr[501]), .rdlo_out(a1_wr[1525]));
			radix2 #(.width(width)) rd_st0_502  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[502]), .rdlo_in(a0_wr[1526]),  .coef_in(coef[502]), .rdup_out(a1_wr[502]), .rdlo_out(a1_wr[1526]));
			radix2 #(.width(width)) rd_st0_503  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[503]), .rdlo_in(a0_wr[1527]),  .coef_in(coef[503]), .rdup_out(a1_wr[503]), .rdlo_out(a1_wr[1527]));
			radix2 #(.width(width)) rd_st0_504  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[504]), .rdlo_in(a0_wr[1528]),  .coef_in(coef[504]), .rdup_out(a1_wr[504]), .rdlo_out(a1_wr[1528]));
			radix2 #(.width(width)) rd_st0_505  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[505]), .rdlo_in(a0_wr[1529]),  .coef_in(coef[505]), .rdup_out(a1_wr[505]), .rdlo_out(a1_wr[1529]));
			radix2 #(.width(width)) rd_st0_506  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[506]), .rdlo_in(a0_wr[1530]),  .coef_in(coef[506]), .rdup_out(a1_wr[506]), .rdlo_out(a1_wr[1530]));
			radix2 #(.width(width)) rd_st0_507  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[507]), .rdlo_in(a0_wr[1531]),  .coef_in(coef[507]), .rdup_out(a1_wr[507]), .rdlo_out(a1_wr[1531]));
			radix2 #(.width(width)) rd_st0_508  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[508]), .rdlo_in(a0_wr[1532]),  .coef_in(coef[508]), .rdup_out(a1_wr[508]), .rdlo_out(a1_wr[1532]));
			radix2 #(.width(width)) rd_st0_509  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[509]), .rdlo_in(a0_wr[1533]),  .coef_in(coef[509]), .rdup_out(a1_wr[509]), .rdlo_out(a1_wr[1533]));
			radix2 #(.width(width)) rd_st0_510  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[510]), .rdlo_in(a0_wr[1534]),  .coef_in(coef[510]), .rdup_out(a1_wr[510]), .rdlo_out(a1_wr[1534]));
			radix2 #(.width(width)) rd_st0_511  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[511]), .rdlo_in(a0_wr[1535]),  .coef_in(coef[511]), .rdup_out(a1_wr[511]), .rdlo_out(a1_wr[1535]));
			radix2 #(.width(width)) rd_st0_512  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[512]), .rdlo_in(a0_wr[1536]),  .coef_in(coef[512]), .rdup_out(a1_wr[512]), .rdlo_out(a1_wr[1536]));
			radix2 #(.width(width)) rd_st0_513  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[513]), .rdlo_in(a0_wr[1537]),  .coef_in(coef[513]), .rdup_out(a1_wr[513]), .rdlo_out(a1_wr[1537]));
			radix2 #(.width(width)) rd_st0_514  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[514]), .rdlo_in(a0_wr[1538]),  .coef_in(coef[514]), .rdup_out(a1_wr[514]), .rdlo_out(a1_wr[1538]));
			radix2 #(.width(width)) rd_st0_515  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[515]), .rdlo_in(a0_wr[1539]),  .coef_in(coef[515]), .rdup_out(a1_wr[515]), .rdlo_out(a1_wr[1539]));
			radix2 #(.width(width)) rd_st0_516  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[516]), .rdlo_in(a0_wr[1540]),  .coef_in(coef[516]), .rdup_out(a1_wr[516]), .rdlo_out(a1_wr[1540]));
			radix2 #(.width(width)) rd_st0_517  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[517]), .rdlo_in(a0_wr[1541]),  .coef_in(coef[517]), .rdup_out(a1_wr[517]), .rdlo_out(a1_wr[1541]));
			radix2 #(.width(width)) rd_st0_518  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[518]), .rdlo_in(a0_wr[1542]),  .coef_in(coef[518]), .rdup_out(a1_wr[518]), .rdlo_out(a1_wr[1542]));
			radix2 #(.width(width)) rd_st0_519  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[519]), .rdlo_in(a0_wr[1543]),  .coef_in(coef[519]), .rdup_out(a1_wr[519]), .rdlo_out(a1_wr[1543]));
			radix2 #(.width(width)) rd_st0_520  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[520]), .rdlo_in(a0_wr[1544]),  .coef_in(coef[520]), .rdup_out(a1_wr[520]), .rdlo_out(a1_wr[1544]));
			radix2 #(.width(width)) rd_st0_521  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[521]), .rdlo_in(a0_wr[1545]),  .coef_in(coef[521]), .rdup_out(a1_wr[521]), .rdlo_out(a1_wr[1545]));
			radix2 #(.width(width)) rd_st0_522  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[522]), .rdlo_in(a0_wr[1546]),  .coef_in(coef[522]), .rdup_out(a1_wr[522]), .rdlo_out(a1_wr[1546]));
			radix2 #(.width(width)) rd_st0_523  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[523]), .rdlo_in(a0_wr[1547]),  .coef_in(coef[523]), .rdup_out(a1_wr[523]), .rdlo_out(a1_wr[1547]));
			radix2 #(.width(width)) rd_st0_524  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[524]), .rdlo_in(a0_wr[1548]),  .coef_in(coef[524]), .rdup_out(a1_wr[524]), .rdlo_out(a1_wr[1548]));
			radix2 #(.width(width)) rd_st0_525  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[525]), .rdlo_in(a0_wr[1549]),  .coef_in(coef[525]), .rdup_out(a1_wr[525]), .rdlo_out(a1_wr[1549]));
			radix2 #(.width(width)) rd_st0_526  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[526]), .rdlo_in(a0_wr[1550]),  .coef_in(coef[526]), .rdup_out(a1_wr[526]), .rdlo_out(a1_wr[1550]));
			radix2 #(.width(width)) rd_st0_527  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[527]), .rdlo_in(a0_wr[1551]),  .coef_in(coef[527]), .rdup_out(a1_wr[527]), .rdlo_out(a1_wr[1551]));
			radix2 #(.width(width)) rd_st0_528  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[528]), .rdlo_in(a0_wr[1552]),  .coef_in(coef[528]), .rdup_out(a1_wr[528]), .rdlo_out(a1_wr[1552]));
			radix2 #(.width(width)) rd_st0_529  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[529]), .rdlo_in(a0_wr[1553]),  .coef_in(coef[529]), .rdup_out(a1_wr[529]), .rdlo_out(a1_wr[1553]));
			radix2 #(.width(width)) rd_st0_530  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[530]), .rdlo_in(a0_wr[1554]),  .coef_in(coef[530]), .rdup_out(a1_wr[530]), .rdlo_out(a1_wr[1554]));
			radix2 #(.width(width)) rd_st0_531  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[531]), .rdlo_in(a0_wr[1555]),  .coef_in(coef[531]), .rdup_out(a1_wr[531]), .rdlo_out(a1_wr[1555]));
			radix2 #(.width(width)) rd_st0_532  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[532]), .rdlo_in(a0_wr[1556]),  .coef_in(coef[532]), .rdup_out(a1_wr[532]), .rdlo_out(a1_wr[1556]));
			radix2 #(.width(width)) rd_st0_533  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[533]), .rdlo_in(a0_wr[1557]),  .coef_in(coef[533]), .rdup_out(a1_wr[533]), .rdlo_out(a1_wr[1557]));
			radix2 #(.width(width)) rd_st0_534  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[534]), .rdlo_in(a0_wr[1558]),  .coef_in(coef[534]), .rdup_out(a1_wr[534]), .rdlo_out(a1_wr[1558]));
			radix2 #(.width(width)) rd_st0_535  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[535]), .rdlo_in(a0_wr[1559]),  .coef_in(coef[535]), .rdup_out(a1_wr[535]), .rdlo_out(a1_wr[1559]));
			radix2 #(.width(width)) rd_st0_536  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[536]), .rdlo_in(a0_wr[1560]),  .coef_in(coef[536]), .rdup_out(a1_wr[536]), .rdlo_out(a1_wr[1560]));
			radix2 #(.width(width)) rd_st0_537  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[537]), .rdlo_in(a0_wr[1561]),  .coef_in(coef[537]), .rdup_out(a1_wr[537]), .rdlo_out(a1_wr[1561]));
			radix2 #(.width(width)) rd_st0_538  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[538]), .rdlo_in(a0_wr[1562]),  .coef_in(coef[538]), .rdup_out(a1_wr[538]), .rdlo_out(a1_wr[1562]));
			radix2 #(.width(width)) rd_st0_539  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[539]), .rdlo_in(a0_wr[1563]),  .coef_in(coef[539]), .rdup_out(a1_wr[539]), .rdlo_out(a1_wr[1563]));
			radix2 #(.width(width)) rd_st0_540  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[540]), .rdlo_in(a0_wr[1564]),  .coef_in(coef[540]), .rdup_out(a1_wr[540]), .rdlo_out(a1_wr[1564]));
			radix2 #(.width(width)) rd_st0_541  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[541]), .rdlo_in(a0_wr[1565]),  .coef_in(coef[541]), .rdup_out(a1_wr[541]), .rdlo_out(a1_wr[1565]));
			radix2 #(.width(width)) rd_st0_542  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[542]), .rdlo_in(a0_wr[1566]),  .coef_in(coef[542]), .rdup_out(a1_wr[542]), .rdlo_out(a1_wr[1566]));
			radix2 #(.width(width)) rd_st0_543  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[543]), .rdlo_in(a0_wr[1567]),  .coef_in(coef[543]), .rdup_out(a1_wr[543]), .rdlo_out(a1_wr[1567]));
			radix2 #(.width(width)) rd_st0_544  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[544]), .rdlo_in(a0_wr[1568]),  .coef_in(coef[544]), .rdup_out(a1_wr[544]), .rdlo_out(a1_wr[1568]));
			radix2 #(.width(width)) rd_st0_545  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[545]), .rdlo_in(a0_wr[1569]),  .coef_in(coef[545]), .rdup_out(a1_wr[545]), .rdlo_out(a1_wr[1569]));
			radix2 #(.width(width)) rd_st0_546  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[546]), .rdlo_in(a0_wr[1570]),  .coef_in(coef[546]), .rdup_out(a1_wr[546]), .rdlo_out(a1_wr[1570]));
			radix2 #(.width(width)) rd_st0_547  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[547]), .rdlo_in(a0_wr[1571]),  .coef_in(coef[547]), .rdup_out(a1_wr[547]), .rdlo_out(a1_wr[1571]));
			radix2 #(.width(width)) rd_st0_548  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[548]), .rdlo_in(a0_wr[1572]),  .coef_in(coef[548]), .rdup_out(a1_wr[548]), .rdlo_out(a1_wr[1572]));
			radix2 #(.width(width)) rd_st0_549  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[549]), .rdlo_in(a0_wr[1573]),  .coef_in(coef[549]), .rdup_out(a1_wr[549]), .rdlo_out(a1_wr[1573]));
			radix2 #(.width(width)) rd_st0_550  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[550]), .rdlo_in(a0_wr[1574]),  .coef_in(coef[550]), .rdup_out(a1_wr[550]), .rdlo_out(a1_wr[1574]));
			radix2 #(.width(width)) rd_st0_551  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[551]), .rdlo_in(a0_wr[1575]),  .coef_in(coef[551]), .rdup_out(a1_wr[551]), .rdlo_out(a1_wr[1575]));
			radix2 #(.width(width)) rd_st0_552  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[552]), .rdlo_in(a0_wr[1576]),  .coef_in(coef[552]), .rdup_out(a1_wr[552]), .rdlo_out(a1_wr[1576]));
			radix2 #(.width(width)) rd_st0_553  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[553]), .rdlo_in(a0_wr[1577]),  .coef_in(coef[553]), .rdup_out(a1_wr[553]), .rdlo_out(a1_wr[1577]));
			radix2 #(.width(width)) rd_st0_554  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[554]), .rdlo_in(a0_wr[1578]),  .coef_in(coef[554]), .rdup_out(a1_wr[554]), .rdlo_out(a1_wr[1578]));
			radix2 #(.width(width)) rd_st0_555  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[555]), .rdlo_in(a0_wr[1579]),  .coef_in(coef[555]), .rdup_out(a1_wr[555]), .rdlo_out(a1_wr[1579]));
			radix2 #(.width(width)) rd_st0_556  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[556]), .rdlo_in(a0_wr[1580]),  .coef_in(coef[556]), .rdup_out(a1_wr[556]), .rdlo_out(a1_wr[1580]));
			radix2 #(.width(width)) rd_st0_557  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[557]), .rdlo_in(a0_wr[1581]),  .coef_in(coef[557]), .rdup_out(a1_wr[557]), .rdlo_out(a1_wr[1581]));
			radix2 #(.width(width)) rd_st0_558  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[558]), .rdlo_in(a0_wr[1582]),  .coef_in(coef[558]), .rdup_out(a1_wr[558]), .rdlo_out(a1_wr[1582]));
			radix2 #(.width(width)) rd_st0_559  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[559]), .rdlo_in(a0_wr[1583]),  .coef_in(coef[559]), .rdup_out(a1_wr[559]), .rdlo_out(a1_wr[1583]));
			radix2 #(.width(width)) rd_st0_560  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[560]), .rdlo_in(a0_wr[1584]),  .coef_in(coef[560]), .rdup_out(a1_wr[560]), .rdlo_out(a1_wr[1584]));
			radix2 #(.width(width)) rd_st0_561  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[561]), .rdlo_in(a0_wr[1585]),  .coef_in(coef[561]), .rdup_out(a1_wr[561]), .rdlo_out(a1_wr[1585]));
			radix2 #(.width(width)) rd_st0_562  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[562]), .rdlo_in(a0_wr[1586]),  .coef_in(coef[562]), .rdup_out(a1_wr[562]), .rdlo_out(a1_wr[1586]));
			radix2 #(.width(width)) rd_st0_563  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[563]), .rdlo_in(a0_wr[1587]),  .coef_in(coef[563]), .rdup_out(a1_wr[563]), .rdlo_out(a1_wr[1587]));
			radix2 #(.width(width)) rd_st0_564  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[564]), .rdlo_in(a0_wr[1588]),  .coef_in(coef[564]), .rdup_out(a1_wr[564]), .rdlo_out(a1_wr[1588]));
			radix2 #(.width(width)) rd_st0_565  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[565]), .rdlo_in(a0_wr[1589]),  .coef_in(coef[565]), .rdup_out(a1_wr[565]), .rdlo_out(a1_wr[1589]));
			radix2 #(.width(width)) rd_st0_566  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[566]), .rdlo_in(a0_wr[1590]),  .coef_in(coef[566]), .rdup_out(a1_wr[566]), .rdlo_out(a1_wr[1590]));
			radix2 #(.width(width)) rd_st0_567  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[567]), .rdlo_in(a0_wr[1591]),  .coef_in(coef[567]), .rdup_out(a1_wr[567]), .rdlo_out(a1_wr[1591]));
			radix2 #(.width(width)) rd_st0_568  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[568]), .rdlo_in(a0_wr[1592]),  .coef_in(coef[568]), .rdup_out(a1_wr[568]), .rdlo_out(a1_wr[1592]));
			radix2 #(.width(width)) rd_st0_569  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[569]), .rdlo_in(a0_wr[1593]),  .coef_in(coef[569]), .rdup_out(a1_wr[569]), .rdlo_out(a1_wr[1593]));
			radix2 #(.width(width)) rd_st0_570  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[570]), .rdlo_in(a0_wr[1594]),  .coef_in(coef[570]), .rdup_out(a1_wr[570]), .rdlo_out(a1_wr[1594]));
			radix2 #(.width(width)) rd_st0_571  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[571]), .rdlo_in(a0_wr[1595]),  .coef_in(coef[571]), .rdup_out(a1_wr[571]), .rdlo_out(a1_wr[1595]));
			radix2 #(.width(width)) rd_st0_572  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[572]), .rdlo_in(a0_wr[1596]),  .coef_in(coef[572]), .rdup_out(a1_wr[572]), .rdlo_out(a1_wr[1596]));
			radix2 #(.width(width)) rd_st0_573  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[573]), .rdlo_in(a0_wr[1597]),  .coef_in(coef[573]), .rdup_out(a1_wr[573]), .rdlo_out(a1_wr[1597]));
			radix2 #(.width(width)) rd_st0_574  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[574]), .rdlo_in(a0_wr[1598]),  .coef_in(coef[574]), .rdup_out(a1_wr[574]), .rdlo_out(a1_wr[1598]));
			radix2 #(.width(width)) rd_st0_575  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[575]), .rdlo_in(a0_wr[1599]),  .coef_in(coef[575]), .rdup_out(a1_wr[575]), .rdlo_out(a1_wr[1599]));
			radix2 #(.width(width)) rd_st0_576  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[576]), .rdlo_in(a0_wr[1600]),  .coef_in(coef[576]), .rdup_out(a1_wr[576]), .rdlo_out(a1_wr[1600]));
			radix2 #(.width(width)) rd_st0_577  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[577]), .rdlo_in(a0_wr[1601]),  .coef_in(coef[577]), .rdup_out(a1_wr[577]), .rdlo_out(a1_wr[1601]));
			radix2 #(.width(width)) rd_st0_578  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[578]), .rdlo_in(a0_wr[1602]),  .coef_in(coef[578]), .rdup_out(a1_wr[578]), .rdlo_out(a1_wr[1602]));
			radix2 #(.width(width)) rd_st0_579  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[579]), .rdlo_in(a0_wr[1603]),  .coef_in(coef[579]), .rdup_out(a1_wr[579]), .rdlo_out(a1_wr[1603]));
			radix2 #(.width(width)) rd_st0_580  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[580]), .rdlo_in(a0_wr[1604]),  .coef_in(coef[580]), .rdup_out(a1_wr[580]), .rdlo_out(a1_wr[1604]));
			radix2 #(.width(width)) rd_st0_581  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[581]), .rdlo_in(a0_wr[1605]),  .coef_in(coef[581]), .rdup_out(a1_wr[581]), .rdlo_out(a1_wr[1605]));
			radix2 #(.width(width)) rd_st0_582  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[582]), .rdlo_in(a0_wr[1606]),  .coef_in(coef[582]), .rdup_out(a1_wr[582]), .rdlo_out(a1_wr[1606]));
			radix2 #(.width(width)) rd_st0_583  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[583]), .rdlo_in(a0_wr[1607]),  .coef_in(coef[583]), .rdup_out(a1_wr[583]), .rdlo_out(a1_wr[1607]));
			radix2 #(.width(width)) rd_st0_584  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[584]), .rdlo_in(a0_wr[1608]),  .coef_in(coef[584]), .rdup_out(a1_wr[584]), .rdlo_out(a1_wr[1608]));
			radix2 #(.width(width)) rd_st0_585  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[585]), .rdlo_in(a0_wr[1609]),  .coef_in(coef[585]), .rdup_out(a1_wr[585]), .rdlo_out(a1_wr[1609]));
			radix2 #(.width(width)) rd_st0_586  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[586]), .rdlo_in(a0_wr[1610]),  .coef_in(coef[586]), .rdup_out(a1_wr[586]), .rdlo_out(a1_wr[1610]));
			radix2 #(.width(width)) rd_st0_587  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[587]), .rdlo_in(a0_wr[1611]),  .coef_in(coef[587]), .rdup_out(a1_wr[587]), .rdlo_out(a1_wr[1611]));
			radix2 #(.width(width)) rd_st0_588  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[588]), .rdlo_in(a0_wr[1612]),  .coef_in(coef[588]), .rdup_out(a1_wr[588]), .rdlo_out(a1_wr[1612]));
			radix2 #(.width(width)) rd_st0_589  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[589]), .rdlo_in(a0_wr[1613]),  .coef_in(coef[589]), .rdup_out(a1_wr[589]), .rdlo_out(a1_wr[1613]));
			radix2 #(.width(width)) rd_st0_590  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[590]), .rdlo_in(a0_wr[1614]),  .coef_in(coef[590]), .rdup_out(a1_wr[590]), .rdlo_out(a1_wr[1614]));
			radix2 #(.width(width)) rd_st0_591  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[591]), .rdlo_in(a0_wr[1615]),  .coef_in(coef[591]), .rdup_out(a1_wr[591]), .rdlo_out(a1_wr[1615]));
			radix2 #(.width(width)) rd_st0_592  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[592]), .rdlo_in(a0_wr[1616]),  .coef_in(coef[592]), .rdup_out(a1_wr[592]), .rdlo_out(a1_wr[1616]));
			radix2 #(.width(width)) rd_st0_593  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[593]), .rdlo_in(a0_wr[1617]),  .coef_in(coef[593]), .rdup_out(a1_wr[593]), .rdlo_out(a1_wr[1617]));
			radix2 #(.width(width)) rd_st0_594  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[594]), .rdlo_in(a0_wr[1618]),  .coef_in(coef[594]), .rdup_out(a1_wr[594]), .rdlo_out(a1_wr[1618]));
			radix2 #(.width(width)) rd_st0_595  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[595]), .rdlo_in(a0_wr[1619]),  .coef_in(coef[595]), .rdup_out(a1_wr[595]), .rdlo_out(a1_wr[1619]));
			radix2 #(.width(width)) rd_st0_596  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[596]), .rdlo_in(a0_wr[1620]),  .coef_in(coef[596]), .rdup_out(a1_wr[596]), .rdlo_out(a1_wr[1620]));
			radix2 #(.width(width)) rd_st0_597  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[597]), .rdlo_in(a0_wr[1621]),  .coef_in(coef[597]), .rdup_out(a1_wr[597]), .rdlo_out(a1_wr[1621]));
			radix2 #(.width(width)) rd_st0_598  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[598]), .rdlo_in(a0_wr[1622]),  .coef_in(coef[598]), .rdup_out(a1_wr[598]), .rdlo_out(a1_wr[1622]));
			radix2 #(.width(width)) rd_st0_599  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[599]), .rdlo_in(a0_wr[1623]),  .coef_in(coef[599]), .rdup_out(a1_wr[599]), .rdlo_out(a1_wr[1623]));
			radix2 #(.width(width)) rd_st0_600  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[600]), .rdlo_in(a0_wr[1624]),  .coef_in(coef[600]), .rdup_out(a1_wr[600]), .rdlo_out(a1_wr[1624]));
			radix2 #(.width(width)) rd_st0_601  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[601]), .rdlo_in(a0_wr[1625]),  .coef_in(coef[601]), .rdup_out(a1_wr[601]), .rdlo_out(a1_wr[1625]));
			radix2 #(.width(width)) rd_st0_602  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[602]), .rdlo_in(a0_wr[1626]),  .coef_in(coef[602]), .rdup_out(a1_wr[602]), .rdlo_out(a1_wr[1626]));
			radix2 #(.width(width)) rd_st0_603  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[603]), .rdlo_in(a0_wr[1627]),  .coef_in(coef[603]), .rdup_out(a1_wr[603]), .rdlo_out(a1_wr[1627]));
			radix2 #(.width(width)) rd_st0_604  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[604]), .rdlo_in(a0_wr[1628]),  .coef_in(coef[604]), .rdup_out(a1_wr[604]), .rdlo_out(a1_wr[1628]));
			radix2 #(.width(width)) rd_st0_605  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[605]), .rdlo_in(a0_wr[1629]),  .coef_in(coef[605]), .rdup_out(a1_wr[605]), .rdlo_out(a1_wr[1629]));
			radix2 #(.width(width)) rd_st0_606  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[606]), .rdlo_in(a0_wr[1630]),  .coef_in(coef[606]), .rdup_out(a1_wr[606]), .rdlo_out(a1_wr[1630]));
			radix2 #(.width(width)) rd_st0_607  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[607]), .rdlo_in(a0_wr[1631]),  .coef_in(coef[607]), .rdup_out(a1_wr[607]), .rdlo_out(a1_wr[1631]));
			radix2 #(.width(width)) rd_st0_608  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[608]), .rdlo_in(a0_wr[1632]),  .coef_in(coef[608]), .rdup_out(a1_wr[608]), .rdlo_out(a1_wr[1632]));
			radix2 #(.width(width)) rd_st0_609  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[609]), .rdlo_in(a0_wr[1633]),  .coef_in(coef[609]), .rdup_out(a1_wr[609]), .rdlo_out(a1_wr[1633]));
			radix2 #(.width(width)) rd_st0_610  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[610]), .rdlo_in(a0_wr[1634]),  .coef_in(coef[610]), .rdup_out(a1_wr[610]), .rdlo_out(a1_wr[1634]));
			radix2 #(.width(width)) rd_st0_611  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[611]), .rdlo_in(a0_wr[1635]),  .coef_in(coef[611]), .rdup_out(a1_wr[611]), .rdlo_out(a1_wr[1635]));
			radix2 #(.width(width)) rd_st0_612  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[612]), .rdlo_in(a0_wr[1636]),  .coef_in(coef[612]), .rdup_out(a1_wr[612]), .rdlo_out(a1_wr[1636]));
			radix2 #(.width(width)) rd_st0_613  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[613]), .rdlo_in(a0_wr[1637]),  .coef_in(coef[613]), .rdup_out(a1_wr[613]), .rdlo_out(a1_wr[1637]));
			radix2 #(.width(width)) rd_st0_614  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[614]), .rdlo_in(a0_wr[1638]),  .coef_in(coef[614]), .rdup_out(a1_wr[614]), .rdlo_out(a1_wr[1638]));
			radix2 #(.width(width)) rd_st0_615  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[615]), .rdlo_in(a0_wr[1639]),  .coef_in(coef[615]), .rdup_out(a1_wr[615]), .rdlo_out(a1_wr[1639]));
			radix2 #(.width(width)) rd_st0_616  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[616]), .rdlo_in(a0_wr[1640]),  .coef_in(coef[616]), .rdup_out(a1_wr[616]), .rdlo_out(a1_wr[1640]));
			radix2 #(.width(width)) rd_st0_617  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[617]), .rdlo_in(a0_wr[1641]),  .coef_in(coef[617]), .rdup_out(a1_wr[617]), .rdlo_out(a1_wr[1641]));
			radix2 #(.width(width)) rd_st0_618  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[618]), .rdlo_in(a0_wr[1642]),  .coef_in(coef[618]), .rdup_out(a1_wr[618]), .rdlo_out(a1_wr[1642]));
			radix2 #(.width(width)) rd_st0_619  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[619]), .rdlo_in(a0_wr[1643]),  .coef_in(coef[619]), .rdup_out(a1_wr[619]), .rdlo_out(a1_wr[1643]));
			radix2 #(.width(width)) rd_st0_620  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[620]), .rdlo_in(a0_wr[1644]),  .coef_in(coef[620]), .rdup_out(a1_wr[620]), .rdlo_out(a1_wr[1644]));
			radix2 #(.width(width)) rd_st0_621  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[621]), .rdlo_in(a0_wr[1645]),  .coef_in(coef[621]), .rdup_out(a1_wr[621]), .rdlo_out(a1_wr[1645]));
			radix2 #(.width(width)) rd_st0_622  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[622]), .rdlo_in(a0_wr[1646]),  .coef_in(coef[622]), .rdup_out(a1_wr[622]), .rdlo_out(a1_wr[1646]));
			radix2 #(.width(width)) rd_st0_623  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[623]), .rdlo_in(a0_wr[1647]),  .coef_in(coef[623]), .rdup_out(a1_wr[623]), .rdlo_out(a1_wr[1647]));
			radix2 #(.width(width)) rd_st0_624  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[624]), .rdlo_in(a0_wr[1648]),  .coef_in(coef[624]), .rdup_out(a1_wr[624]), .rdlo_out(a1_wr[1648]));
			radix2 #(.width(width)) rd_st0_625  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[625]), .rdlo_in(a0_wr[1649]),  .coef_in(coef[625]), .rdup_out(a1_wr[625]), .rdlo_out(a1_wr[1649]));
			radix2 #(.width(width)) rd_st0_626  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[626]), .rdlo_in(a0_wr[1650]),  .coef_in(coef[626]), .rdup_out(a1_wr[626]), .rdlo_out(a1_wr[1650]));
			radix2 #(.width(width)) rd_st0_627  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[627]), .rdlo_in(a0_wr[1651]),  .coef_in(coef[627]), .rdup_out(a1_wr[627]), .rdlo_out(a1_wr[1651]));
			radix2 #(.width(width)) rd_st0_628  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[628]), .rdlo_in(a0_wr[1652]),  .coef_in(coef[628]), .rdup_out(a1_wr[628]), .rdlo_out(a1_wr[1652]));
			radix2 #(.width(width)) rd_st0_629  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[629]), .rdlo_in(a0_wr[1653]),  .coef_in(coef[629]), .rdup_out(a1_wr[629]), .rdlo_out(a1_wr[1653]));
			radix2 #(.width(width)) rd_st0_630  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[630]), .rdlo_in(a0_wr[1654]),  .coef_in(coef[630]), .rdup_out(a1_wr[630]), .rdlo_out(a1_wr[1654]));
			radix2 #(.width(width)) rd_st0_631  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[631]), .rdlo_in(a0_wr[1655]),  .coef_in(coef[631]), .rdup_out(a1_wr[631]), .rdlo_out(a1_wr[1655]));
			radix2 #(.width(width)) rd_st0_632  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[632]), .rdlo_in(a0_wr[1656]),  .coef_in(coef[632]), .rdup_out(a1_wr[632]), .rdlo_out(a1_wr[1656]));
			radix2 #(.width(width)) rd_st0_633  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[633]), .rdlo_in(a0_wr[1657]),  .coef_in(coef[633]), .rdup_out(a1_wr[633]), .rdlo_out(a1_wr[1657]));
			radix2 #(.width(width)) rd_st0_634  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[634]), .rdlo_in(a0_wr[1658]),  .coef_in(coef[634]), .rdup_out(a1_wr[634]), .rdlo_out(a1_wr[1658]));
			radix2 #(.width(width)) rd_st0_635  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[635]), .rdlo_in(a0_wr[1659]),  .coef_in(coef[635]), .rdup_out(a1_wr[635]), .rdlo_out(a1_wr[1659]));
			radix2 #(.width(width)) rd_st0_636  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[636]), .rdlo_in(a0_wr[1660]),  .coef_in(coef[636]), .rdup_out(a1_wr[636]), .rdlo_out(a1_wr[1660]));
			radix2 #(.width(width)) rd_st0_637  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[637]), .rdlo_in(a0_wr[1661]),  .coef_in(coef[637]), .rdup_out(a1_wr[637]), .rdlo_out(a1_wr[1661]));
			radix2 #(.width(width)) rd_st0_638  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[638]), .rdlo_in(a0_wr[1662]),  .coef_in(coef[638]), .rdup_out(a1_wr[638]), .rdlo_out(a1_wr[1662]));
			radix2 #(.width(width)) rd_st0_639  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[639]), .rdlo_in(a0_wr[1663]),  .coef_in(coef[639]), .rdup_out(a1_wr[639]), .rdlo_out(a1_wr[1663]));
			radix2 #(.width(width)) rd_st0_640  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[640]), .rdlo_in(a0_wr[1664]),  .coef_in(coef[640]), .rdup_out(a1_wr[640]), .rdlo_out(a1_wr[1664]));
			radix2 #(.width(width)) rd_st0_641  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[641]), .rdlo_in(a0_wr[1665]),  .coef_in(coef[641]), .rdup_out(a1_wr[641]), .rdlo_out(a1_wr[1665]));
			radix2 #(.width(width)) rd_st0_642  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[642]), .rdlo_in(a0_wr[1666]),  .coef_in(coef[642]), .rdup_out(a1_wr[642]), .rdlo_out(a1_wr[1666]));
			radix2 #(.width(width)) rd_st0_643  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[643]), .rdlo_in(a0_wr[1667]),  .coef_in(coef[643]), .rdup_out(a1_wr[643]), .rdlo_out(a1_wr[1667]));
			radix2 #(.width(width)) rd_st0_644  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[644]), .rdlo_in(a0_wr[1668]),  .coef_in(coef[644]), .rdup_out(a1_wr[644]), .rdlo_out(a1_wr[1668]));
			radix2 #(.width(width)) rd_st0_645  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[645]), .rdlo_in(a0_wr[1669]),  .coef_in(coef[645]), .rdup_out(a1_wr[645]), .rdlo_out(a1_wr[1669]));
			radix2 #(.width(width)) rd_st0_646  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[646]), .rdlo_in(a0_wr[1670]),  .coef_in(coef[646]), .rdup_out(a1_wr[646]), .rdlo_out(a1_wr[1670]));
			radix2 #(.width(width)) rd_st0_647  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[647]), .rdlo_in(a0_wr[1671]),  .coef_in(coef[647]), .rdup_out(a1_wr[647]), .rdlo_out(a1_wr[1671]));
			radix2 #(.width(width)) rd_st0_648  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[648]), .rdlo_in(a0_wr[1672]),  .coef_in(coef[648]), .rdup_out(a1_wr[648]), .rdlo_out(a1_wr[1672]));
			radix2 #(.width(width)) rd_st0_649  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[649]), .rdlo_in(a0_wr[1673]),  .coef_in(coef[649]), .rdup_out(a1_wr[649]), .rdlo_out(a1_wr[1673]));
			radix2 #(.width(width)) rd_st0_650  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[650]), .rdlo_in(a0_wr[1674]),  .coef_in(coef[650]), .rdup_out(a1_wr[650]), .rdlo_out(a1_wr[1674]));
			radix2 #(.width(width)) rd_st0_651  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[651]), .rdlo_in(a0_wr[1675]),  .coef_in(coef[651]), .rdup_out(a1_wr[651]), .rdlo_out(a1_wr[1675]));
			radix2 #(.width(width)) rd_st0_652  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[652]), .rdlo_in(a0_wr[1676]),  .coef_in(coef[652]), .rdup_out(a1_wr[652]), .rdlo_out(a1_wr[1676]));
			radix2 #(.width(width)) rd_st0_653  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[653]), .rdlo_in(a0_wr[1677]),  .coef_in(coef[653]), .rdup_out(a1_wr[653]), .rdlo_out(a1_wr[1677]));
			radix2 #(.width(width)) rd_st0_654  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[654]), .rdlo_in(a0_wr[1678]),  .coef_in(coef[654]), .rdup_out(a1_wr[654]), .rdlo_out(a1_wr[1678]));
			radix2 #(.width(width)) rd_st0_655  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[655]), .rdlo_in(a0_wr[1679]),  .coef_in(coef[655]), .rdup_out(a1_wr[655]), .rdlo_out(a1_wr[1679]));
			radix2 #(.width(width)) rd_st0_656  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[656]), .rdlo_in(a0_wr[1680]),  .coef_in(coef[656]), .rdup_out(a1_wr[656]), .rdlo_out(a1_wr[1680]));
			radix2 #(.width(width)) rd_st0_657  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[657]), .rdlo_in(a0_wr[1681]),  .coef_in(coef[657]), .rdup_out(a1_wr[657]), .rdlo_out(a1_wr[1681]));
			radix2 #(.width(width)) rd_st0_658  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[658]), .rdlo_in(a0_wr[1682]),  .coef_in(coef[658]), .rdup_out(a1_wr[658]), .rdlo_out(a1_wr[1682]));
			radix2 #(.width(width)) rd_st0_659  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[659]), .rdlo_in(a0_wr[1683]),  .coef_in(coef[659]), .rdup_out(a1_wr[659]), .rdlo_out(a1_wr[1683]));
			radix2 #(.width(width)) rd_st0_660  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[660]), .rdlo_in(a0_wr[1684]),  .coef_in(coef[660]), .rdup_out(a1_wr[660]), .rdlo_out(a1_wr[1684]));
			radix2 #(.width(width)) rd_st0_661  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[661]), .rdlo_in(a0_wr[1685]),  .coef_in(coef[661]), .rdup_out(a1_wr[661]), .rdlo_out(a1_wr[1685]));
			radix2 #(.width(width)) rd_st0_662  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[662]), .rdlo_in(a0_wr[1686]),  .coef_in(coef[662]), .rdup_out(a1_wr[662]), .rdlo_out(a1_wr[1686]));
			radix2 #(.width(width)) rd_st0_663  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[663]), .rdlo_in(a0_wr[1687]),  .coef_in(coef[663]), .rdup_out(a1_wr[663]), .rdlo_out(a1_wr[1687]));
			radix2 #(.width(width)) rd_st0_664  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[664]), .rdlo_in(a0_wr[1688]),  .coef_in(coef[664]), .rdup_out(a1_wr[664]), .rdlo_out(a1_wr[1688]));
			radix2 #(.width(width)) rd_st0_665  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[665]), .rdlo_in(a0_wr[1689]),  .coef_in(coef[665]), .rdup_out(a1_wr[665]), .rdlo_out(a1_wr[1689]));
			radix2 #(.width(width)) rd_st0_666  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[666]), .rdlo_in(a0_wr[1690]),  .coef_in(coef[666]), .rdup_out(a1_wr[666]), .rdlo_out(a1_wr[1690]));
			radix2 #(.width(width)) rd_st0_667  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[667]), .rdlo_in(a0_wr[1691]),  .coef_in(coef[667]), .rdup_out(a1_wr[667]), .rdlo_out(a1_wr[1691]));
			radix2 #(.width(width)) rd_st0_668  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[668]), .rdlo_in(a0_wr[1692]),  .coef_in(coef[668]), .rdup_out(a1_wr[668]), .rdlo_out(a1_wr[1692]));
			radix2 #(.width(width)) rd_st0_669  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[669]), .rdlo_in(a0_wr[1693]),  .coef_in(coef[669]), .rdup_out(a1_wr[669]), .rdlo_out(a1_wr[1693]));
			radix2 #(.width(width)) rd_st0_670  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[670]), .rdlo_in(a0_wr[1694]),  .coef_in(coef[670]), .rdup_out(a1_wr[670]), .rdlo_out(a1_wr[1694]));
			radix2 #(.width(width)) rd_st0_671  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[671]), .rdlo_in(a0_wr[1695]),  .coef_in(coef[671]), .rdup_out(a1_wr[671]), .rdlo_out(a1_wr[1695]));
			radix2 #(.width(width)) rd_st0_672  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[672]), .rdlo_in(a0_wr[1696]),  .coef_in(coef[672]), .rdup_out(a1_wr[672]), .rdlo_out(a1_wr[1696]));
			radix2 #(.width(width)) rd_st0_673  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[673]), .rdlo_in(a0_wr[1697]),  .coef_in(coef[673]), .rdup_out(a1_wr[673]), .rdlo_out(a1_wr[1697]));
			radix2 #(.width(width)) rd_st0_674  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[674]), .rdlo_in(a0_wr[1698]),  .coef_in(coef[674]), .rdup_out(a1_wr[674]), .rdlo_out(a1_wr[1698]));
			radix2 #(.width(width)) rd_st0_675  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[675]), .rdlo_in(a0_wr[1699]),  .coef_in(coef[675]), .rdup_out(a1_wr[675]), .rdlo_out(a1_wr[1699]));
			radix2 #(.width(width)) rd_st0_676  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[676]), .rdlo_in(a0_wr[1700]),  .coef_in(coef[676]), .rdup_out(a1_wr[676]), .rdlo_out(a1_wr[1700]));
			radix2 #(.width(width)) rd_st0_677  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[677]), .rdlo_in(a0_wr[1701]),  .coef_in(coef[677]), .rdup_out(a1_wr[677]), .rdlo_out(a1_wr[1701]));
			radix2 #(.width(width)) rd_st0_678  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[678]), .rdlo_in(a0_wr[1702]),  .coef_in(coef[678]), .rdup_out(a1_wr[678]), .rdlo_out(a1_wr[1702]));
			radix2 #(.width(width)) rd_st0_679  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[679]), .rdlo_in(a0_wr[1703]),  .coef_in(coef[679]), .rdup_out(a1_wr[679]), .rdlo_out(a1_wr[1703]));
			radix2 #(.width(width)) rd_st0_680  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[680]), .rdlo_in(a0_wr[1704]),  .coef_in(coef[680]), .rdup_out(a1_wr[680]), .rdlo_out(a1_wr[1704]));
			radix2 #(.width(width)) rd_st0_681  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[681]), .rdlo_in(a0_wr[1705]),  .coef_in(coef[681]), .rdup_out(a1_wr[681]), .rdlo_out(a1_wr[1705]));
			radix2 #(.width(width)) rd_st0_682  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[682]), .rdlo_in(a0_wr[1706]),  .coef_in(coef[682]), .rdup_out(a1_wr[682]), .rdlo_out(a1_wr[1706]));
			radix2 #(.width(width)) rd_st0_683  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[683]), .rdlo_in(a0_wr[1707]),  .coef_in(coef[683]), .rdup_out(a1_wr[683]), .rdlo_out(a1_wr[1707]));
			radix2 #(.width(width)) rd_st0_684  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[684]), .rdlo_in(a0_wr[1708]),  .coef_in(coef[684]), .rdup_out(a1_wr[684]), .rdlo_out(a1_wr[1708]));
			radix2 #(.width(width)) rd_st0_685  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[685]), .rdlo_in(a0_wr[1709]),  .coef_in(coef[685]), .rdup_out(a1_wr[685]), .rdlo_out(a1_wr[1709]));
			radix2 #(.width(width)) rd_st0_686  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[686]), .rdlo_in(a0_wr[1710]),  .coef_in(coef[686]), .rdup_out(a1_wr[686]), .rdlo_out(a1_wr[1710]));
			radix2 #(.width(width)) rd_st0_687  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[687]), .rdlo_in(a0_wr[1711]),  .coef_in(coef[687]), .rdup_out(a1_wr[687]), .rdlo_out(a1_wr[1711]));
			radix2 #(.width(width)) rd_st0_688  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[688]), .rdlo_in(a0_wr[1712]),  .coef_in(coef[688]), .rdup_out(a1_wr[688]), .rdlo_out(a1_wr[1712]));
			radix2 #(.width(width)) rd_st0_689  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[689]), .rdlo_in(a0_wr[1713]),  .coef_in(coef[689]), .rdup_out(a1_wr[689]), .rdlo_out(a1_wr[1713]));
			radix2 #(.width(width)) rd_st0_690  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[690]), .rdlo_in(a0_wr[1714]),  .coef_in(coef[690]), .rdup_out(a1_wr[690]), .rdlo_out(a1_wr[1714]));
			radix2 #(.width(width)) rd_st0_691  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[691]), .rdlo_in(a0_wr[1715]),  .coef_in(coef[691]), .rdup_out(a1_wr[691]), .rdlo_out(a1_wr[1715]));
			radix2 #(.width(width)) rd_st0_692  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[692]), .rdlo_in(a0_wr[1716]),  .coef_in(coef[692]), .rdup_out(a1_wr[692]), .rdlo_out(a1_wr[1716]));
			radix2 #(.width(width)) rd_st0_693  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[693]), .rdlo_in(a0_wr[1717]),  .coef_in(coef[693]), .rdup_out(a1_wr[693]), .rdlo_out(a1_wr[1717]));
			radix2 #(.width(width)) rd_st0_694  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[694]), .rdlo_in(a0_wr[1718]),  .coef_in(coef[694]), .rdup_out(a1_wr[694]), .rdlo_out(a1_wr[1718]));
			radix2 #(.width(width)) rd_st0_695  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[695]), .rdlo_in(a0_wr[1719]),  .coef_in(coef[695]), .rdup_out(a1_wr[695]), .rdlo_out(a1_wr[1719]));
			radix2 #(.width(width)) rd_st0_696  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[696]), .rdlo_in(a0_wr[1720]),  .coef_in(coef[696]), .rdup_out(a1_wr[696]), .rdlo_out(a1_wr[1720]));
			radix2 #(.width(width)) rd_st0_697  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[697]), .rdlo_in(a0_wr[1721]),  .coef_in(coef[697]), .rdup_out(a1_wr[697]), .rdlo_out(a1_wr[1721]));
			radix2 #(.width(width)) rd_st0_698  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[698]), .rdlo_in(a0_wr[1722]),  .coef_in(coef[698]), .rdup_out(a1_wr[698]), .rdlo_out(a1_wr[1722]));
			radix2 #(.width(width)) rd_st0_699  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[699]), .rdlo_in(a0_wr[1723]),  .coef_in(coef[699]), .rdup_out(a1_wr[699]), .rdlo_out(a1_wr[1723]));
			radix2 #(.width(width)) rd_st0_700  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[700]), .rdlo_in(a0_wr[1724]),  .coef_in(coef[700]), .rdup_out(a1_wr[700]), .rdlo_out(a1_wr[1724]));
			radix2 #(.width(width)) rd_st0_701  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[701]), .rdlo_in(a0_wr[1725]),  .coef_in(coef[701]), .rdup_out(a1_wr[701]), .rdlo_out(a1_wr[1725]));
			radix2 #(.width(width)) rd_st0_702  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[702]), .rdlo_in(a0_wr[1726]),  .coef_in(coef[702]), .rdup_out(a1_wr[702]), .rdlo_out(a1_wr[1726]));
			radix2 #(.width(width)) rd_st0_703  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[703]), .rdlo_in(a0_wr[1727]),  .coef_in(coef[703]), .rdup_out(a1_wr[703]), .rdlo_out(a1_wr[1727]));
			radix2 #(.width(width)) rd_st0_704  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[704]), .rdlo_in(a0_wr[1728]),  .coef_in(coef[704]), .rdup_out(a1_wr[704]), .rdlo_out(a1_wr[1728]));
			radix2 #(.width(width)) rd_st0_705  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[705]), .rdlo_in(a0_wr[1729]),  .coef_in(coef[705]), .rdup_out(a1_wr[705]), .rdlo_out(a1_wr[1729]));
			radix2 #(.width(width)) rd_st0_706  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[706]), .rdlo_in(a0_wr[1730]),  .coef_in(coef[706]), .rdup_out(a1_wr[706]), .rdlo_out(a1_wr[1730]));
			radix2 #(.width(width)) rd_st0_707  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[707]), .rdlo_in(a0_wr[1731]),  .coef_in(coef[707]), .rdup_out(a1_wr[707]), .rdlo_out(a1_wr[1731]));
			radix2 #(.width(width)) rd_st0_708  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[708]), .rdlo_in(a0_wr[1732]),  .coef_in(coef[708]), .rdup_out(a1_wr[708]), .rdlo_out(a1_wr[1732]));
			radix2 #(.width(width)) rd_st0_709  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[709]), .rdlo_in(a0_wr[1733]),  .coef_in(coef[709]), .rdup_out(a1_wr[709]), .rdlo_out(a1_wr[1733]));
			radix2 #(.width(width)) rd_st0_710  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[710]), .rdlo_in(a0_wr[1734]),  .coef_in(coef[710]), .rdup_out(a1_wr[710]), .rdlo_out(a1_wr[1734]));
			radix2 #(.width(width)) rd_st0_711  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[711]), .rdlo_in(a0_wr[1735]),  .coef_in(coef[711]), .rdup_out(a1_wr[711]), .rdlo_out(a1_wr[1735]));
			radix2 #(.width(width)) rd_st0_712  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[712]), .rdlo_in(a0_wr[1736]),  .coef_in(coef[712]), .rdup_out(a1_wr[712]), .rdlo_out(a1_wr[1736]));
			radix2 #(.width(width)) rd_st0_713  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[713]), .rdlo_in(a0_wr[1737]),  .coef_in(coef[713]), .rdup_out(a1_wr[713]), .rdlo_out(a1_wr[1737]));
			radix2 #(.width(width)) rd_st0_714  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[714]), .rdlo_in(a0_wr[1738]),  .coef_in(coef[714]), .rdup_out(a1_wr[714]), .rdlo_out(a1_wr[1738]));
			radix2 #(.width(width)) rd_st0_715  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[715]), .rdlo_in(a0_wr[1739]),  .coef_in(coef[715]), .rdup_out(a1_wr[715]), .rdlo_out(a1_wr[1739]));
			radix2 #(.width(width)) rd_st0_716  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[716]), .rdlo_in(a0_wr[1740]),  .coef_in(coef[716]), .rdup_out(a1_wr[716]), .rdlo_out(a1_wr[1740]));
			radix2 #(.width(width)) rd_st0_717  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[717]), .rdlo_in(a0_wr[1741]),  .coef_in(coef[717]), .rdup_out(a1_wr[717]), .rdlo_out(a1_wr[1741]));
			radix2 #(.width(width)) rd_st0_718  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[718]), .rdlo_in(a0_wr[1742]),  .coef_in(coef[718]), .rdup_out(a1_wr[718]), .rdlo_out(a1_wr[1742]));
			radix2 #(.width(width)) rd_st0_719  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[719]), .rdlo_in(a0_wr[1743]),  .coef_in(coef[719]), .rdup_out(a1_wr[719]), .rdlo_out(a1_wr[1743]));
			radix2 #(.width(width)) rd_st0_720  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[720]), .rdlo_in(a0_wr[1744]),  .coef_in(coef[720]), .rdup_out(a1_wr[720]), .rdlo_out(a1_wr[1744]));
			radix2 #(.width(width)) rd_st0_721  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[721]), .rdlo_in(a0_wr[1745]),  .coef_in(coef[721]), .rdup_out(a1_wr[721]), .rdlo_out(a1_wr[1745]));
			radix2 #(.width(width)) rd_st0_722  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[722]), .rdlo_in(a0_wr[1746]),  .coef_in(coef[722]), .rdup_out(a1_wr[722]), .rdlo_out(a1_wr[1746]));
			radix2 #(.width(width)) rd_st0_723  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[723]), .rdlo_in(a0_wr[1747]),  .coef_in(coef[723]), .rdup_out(a1_wr[723]), .rdlo_out(a1_wr[1747]));
			radix2 #(.width(width)) rd_st0_724  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[724]), .rdlo_in(a0_wr[1748]),  .coef_in(coef[724]), .rdup_out(a1_wr[724]), .rdlo_out(a1_wr[1748]));
			radix2 #(.width(width)) rd_st0_725  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[725]), .rdlo_in(a0_wr[1749]),  .coef_in(coef[725]), .rdup_out(a1_wr[725]), .rdlo_out(a1_wr[1749]));
			radix2 #(.width(width)) rd_st0_726  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[726]), .rdlo_in(a0_wr[1750]),  .coef_in(coef[726]), .rdup_out(a1_wr[726]), .rdlo_out(a1_wr[1750]));
			radix2 #(.width(width)) rd_st0_727  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[727]), .rdlo_in(a0_wr[1751]),  .coef_in(coef[727]), .rdup_out(a1_wr[727]), .rdlo_out(a1_wr[1751]));
			radix2 #(.width(width)) rd_st0_728  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[728]), .rdlo_in(a0_wr[1752]),  .coef_in(coef[728]), .rdup_out(a1_wr[728]), .rdlo_out(a1_wr[1752]));
			radix2 #(.width(width)) rd_st0_729  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[729]), .rdlo_in(a0_wr[1753]),  .coef_in(coef[729]), .rdup_out(a1_wr[729]), .rdlo_out(a1_wr[1753]));
			radix2 #(.width(width)) rd_st0_730  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[730]), .rdlo_in(a0_wr[1754]),  .coef_in(coef[730]), .rdup_out(a1_wr[730]), .rdlo_out(a1_wr[1754]));
			radix2 #(.width(width)) rd_st0_731  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[731]), .rdlo_in(a0_wr[1755]),  .coef_in(coef[731]), .rdup_out(a1_wr[731]), .rdlo_out(a1_wr[1755]));
			radix2 #(.width(width)) rd_st0_732  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[732]), .rdlo_in(a0_wr[1756]),  .coef_in(coef[732]), .rdup_out(a1_wr[732]), .rdlo_out(a1_wr[1756]));
			radix2 #(.width(width)) rd_st0_733  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[733]), .rdlo_in(a0_wr[1757]),  .coef_in(coef[733]), .rdup_out(a1_wr[733]), .rdlo_out(a1_wr[1757]));
			radix2 #(.width(width)) rd_st0_734  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[734]), .rdlo_in(a0_wr[1758]),  .coef_in(coef[734]), .rdup_out(a1_wr[734]), .rdlo_out(a1_wr[1758]));
			radix2 #(.width(width)) rd_st0_735  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[735]), .rdlo_in(a0_wr[1759]),  .coef_in(coef[735]), .rdup_out(a1_wr[735]), .rdlo_out(a1_wr[1759]));
			radix2 #(.width(width)) rd_st0_736  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[736]), .rdlo_in(a0_wr[1760]),  .coef_in(coef[736]), .rdup_out(a1_wr[736]), .rdlo_out(a1_wr[1760]));
			radix2 #(.width(width)) rd_st0_737  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[737]), .rdlo_in(a0_wr[1761]),  .coef_in(coef[737]), .rdup_out(a1_wr[737]), .rdlo_out(a1_wr[1761]));
			radix2 #(.width(width)) rd_st0_738  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[738]), .rdlo_in(a0_wr[1762]),  .coef_in(coef[738]), .rdup_out(a1_wr[738]), .rdlo_out(a1_wr[1762]));
			radix2 #(.width(width)) rd_st0_739  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[739]), .rdlo_in(a0_wr[1763]),  .coef_in(coef[739]), .rdup_out(a1_wr[739]), .rdlo_out(a1_wr[1763]));
			radix2 #(.width(width)) rd_st0_740  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[740]), .rdlo_in(a0_wr[1764]),  .coef_in(coef[740]), .rdup_out(a1_wr[740]), .rdlo_out(a1_wr[1764]));
			radix2 #(.width(width)) rd_st0_741  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[741]), .rdlo_in(a0_wr[1765]),  .coef_in(coef[741]), .rdup_out(a1_wr[741]), .rdlo_out(a1_wr[1765]));
			radix2 #(.width(width)) rd_st0_742  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[742]), .rdlo_in(a0_wr[1766]),  .coef_in(coef[742]), .rdup_out(a1_wr[742]), .rdlo_out(a1_wr[1766]));
			radix2 #(.width(width)) rd_st0_743  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[743]), .rdlo_in(a0_wr[1767]),  .coef_in(coef[743]), .rdup_out(a1_wr[743]), .rdlo_out(a1_wr[1767]));
			radix2 #(.width(width)) rd_st0_744  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[744]), .rdlo_in(a0_wr[1768]),  .coef_in(coef[744]), .rdup_out(a1_wr[744]), .rdlo_out(a1_wr[1768]));
			radix2 #(.width(width)) rd_st0_745  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[745]), .rdlo_in(a0_wr[1769]),  .coef_in(coef[745]), .rdup_out(a1_wr[745]), .rdlo_out(a1_wr[1769]));
			radix2 #(.width(width)) rd_st0_746  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[746]), .rdlo_in(a0_wr[1770]),  .coef_in(coef[746]), .rdup_out(a1_wr[746]), .rdlo_out(a1_wr[1770]));
			radix2 #(.width(width)) rd_st0_747  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[747]), .rdlo_in(a0_wr[1771]),  .coef_in(coef[747]), .rdup_out(a1_wr[747]), .rdlo_out(a1_wr[1771]));
			radix2 #(.width(width)) rd_st0_748  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[748]), .rdlo_in(a0_wr[1772]),  .coef_in(coef[748]), .rdup_out(a1_wr[748]), .rdlo_out(a1_wr[1772]));
			radix2 #(.width(width)) rd_st0_749  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[749]), .rdlo_in(a0_wr[1773]),  .coef_in(coef[749]), .rdup_out(a1_wr[749]), .rdlo_out(a1_wr[1773]));
			radix2 #(.width(width)) rd_st0_750  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[750]), .rdlo_in(a0_wr[1774]),  .coef_in(coef[750]), .rdup_out(a1_wr[750]), .rdlo_out(a1_wr[1774]));
			radix2 #(.width(width)) rd_st0_751  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[751]), .rdlo_in(a0_wr[1775]),  .coef_in(coef[751]), .rdup_out(a1_wr[751]), .rdlo_out(a1_wr[1775]));
			radix2 #(.width(width)) rd_st0_752  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[752]), .rdlo_in(a0_wr[1776]),  .coef_in(coef[752]), .rdup_out(a1_wr[752]), .rdlo_out(a1_wr[1776]));
			radix2 #(.width(width)) rd_st0_753  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[753]), .rdlo_in(a0_wr[1777]),  .coef_in(coef[753]), .rdup_out(a1_wr[753]), .rdlo_out(a1_wr[1777]));
			radix2 #(.width(width)) rd_st0_754  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[754]), .rdlo_in(a0_wr[1778]),  .coef_in(coef[754]), .rdup_out(a1_wr[754]), .rdlo_out(a1_wr[1778]));
			radix2 #(.width(width)) rd_st0_755  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[755]), .rdlo_in(a0_wr[1779]),  .coef_in(coef[755]), .rdup_out(a1_wr[755]), .rdlo_out(a1_wr[1779]));
			radix2 #(.width(width)) rd_st0_756  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[756]), .rdlo_in(a0_wr[1780]),  .coef_in(coef[756]), .rdup_out(a1_wr[756]), .rdlo_out(a1_wr[1780]));
			radix2 #(.width(width)) rd_st0_757  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[757]), .rdlo_in(a0_wr[1781]),  .coef_in(coef[757]), .rdup_out(a1_wr[757]), .rdlo_out(a1_wr[1781]));
			radix2 #(.width(width)) rd_st0_758  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[758]), .rdlo_in(a0_wr[1782]),  .coef_in(coef[758]), .rdup_out(a1_wr[758]), .rdlo_out(a1_wr[1782]));
			radix2 #(.width(width)) rd_st0_759  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[759]), .rdlo_in(a0_wr[1783]),  .coef_in(coef[759]), .rdup_out(a1_wr[759]), .rdlo_out(a1_wr[1783]));
			radix2 #(.width(width)) rd_st0_760  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[760]), .rdlo_in(a0_wr[1784]),  .coef_in(coef[760]), .rdup_out(a1_wr[760]), .rdlo_out(a1_wr[1784]));
			radix2 #(.width(width)) rd_st0_761  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[761]), .rdlo_in(a0_wr[1785]),  .coef_in(coef[761]), .rdup_out(a1_wr[761]), .rdlo_out(a1_wr[1785]));
			radix2 #(.width(width)) rd_st0_762  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[762]), .rdlo_in(a0_wr[1786]),  .coef_in(coef[762]), .rdup_out(a1_wr[762]), .rdlo_out(a1_wr[1786]));
			radix2 #(.width(width)) rd_st0_763  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[763]), .rdlo_in(a0_wr[1787]),  .coef_in(coef[763]), .rdup_out(a1_wr[763]), .rdlo_out(a1_wr[1787]));
			radix2 #(.width(width)) rd_st0_764  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[764]), .rdlo_in(a0_wr[1788]),  .coef_in(coef[764]), .rdup_out(a1_wr[764]), .rdlo_out(a1_wr[1788]));
			radix2 #(.width(width)) rd_st0_765  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[765]), .rdlo_in(a0_wr[1789]),  .coef_in(coef[765]), .rdup_out(a1_wr[765]), .rdlo_out(a1_wr[1789]));
			radix2 #(.width(width)) rd_st0_766  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[766]), .rdlo_in(a0_wr[1790]),  .coef_in(coef[766]), .rdup_out(a1_wr[766]), .rdlo_out(a1_wr[1790]));
			radix2 #(.width(width)) rd_st0_767  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[767]), .rdlo_in(a0_wr[1791]),  .coef_in(coef[767]), .rdup_out(a1_wr[767]), .rdlo_out(a1_wr[1791]));
			radix2 #(.width(width)) rd_st0_768  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[768]), .rdlo_in(a0_wr[1792]),  .coef_in(coef[768]), .rdup_out(a1_wr[768]), .rdlo_out(a1_wr[1792]));
			radix2 #(.width(width)) rd_st0_769  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[769]), .rdlo_in(a0_wr[1793]),  .coef_in(coef[769]), .rdup_out(a1_wr[769]), .rdlo_out(a1_wr[1793]));
			radix2 #(.width(width)) rd_st0_770  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[770]), .rdlo_in(a0_wr[1794]),  .coef_in(coef[770]), .rdup_out(a1_wr[770]), .rdlo_out(a1_wr[1794]));
			radix2 #(.width(width)) rd_st0_771  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[771]), .rdlo_in(a0_wr[1795]),  .coef_in(coef[771]), .rdup_out(a1_wr[771]), .rdlo_out(a1_wr[1795]));
			radix2 #(.width(width)) rd_st0_772  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[772]), .rdlo_in(a0_wr[1796]),  .coef_in(coef[772]), .rdup_out(a1_wr[772]), .rdlo_out(a1_wr[1796]));
			radix2 #(.width(width)) rd_st0_773  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[773]), .rdlo_in(a0_wr[1797]),  .coef_in(coef[773]), .rdup_out(a1_wr[773]), .rdlo_out(a1_wr[1797]));
			radix2 #(.width(width)) rd_st0_774  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[774]), .rdlo_in(a0_wr[1798]),  .coef_in(coef[774]), .rdup_out(a1_wr[774]), .rdlo_out(a1_wr[1798]));
			radix2 #(.width(width)) rd_st0_775  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[775]), .rdlo_in(a0_wr[1799]),  .coef_in(coef[775]), .rdup_out(a1_wr[775]), .rdlo_out(a1_wr[1799]));
			radix2 #(.width(width)) rd_st0_776  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[776]), .rdlo_in(a0_wr[1800]),  .coef_in(coef[776]), .rdup_out(a1_wr[776]), .rdlo_out(a1_wr[1800]));
			radix2 #(.width(width)) rd_st0_777  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[777]), .rdlo_in(a0_wr[1801]),  .coef_in(coef[777]), .rdup_out(a1_wr[777]), .rdlo_out(a1_wr[1801]));
			radix2 #(.width(width)) rd_st0_778  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[778]), .rdlo_in(a0_wr[1802]),  .coef_in(coef[778]), .rdup_out(a1_wr[778]), .rdlo_out(a1_wr[1802]));
			radix2 #(.width(width)) rd_st0_779  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[779]), .rdlo_in(a0_wr[1803]),  .coef_in(coef[779]), .rdup_out(a1_wr[779]), .rdlo_out(a1_wr[1803]));
			radix2 #(.width(width)) rd_st0_780  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[780]), .rdlo_in(a0_wr[1804]),  .coef_in(coef[780]), .rdup_out(a1_wr[780]), .rdlo_out(a1_wr[1804]));
			radix2 #(.width(width)) rd_st0_781  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[781]), .rdlo_in(a0_wr[1805]),  .coef_in(coef[781]), .rdup_out(a1_wr[781]), .rdlo_out(a1_wr[1805]));
			radix2 #(.width(width)) rd_st0_782  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[782]), .rdlo_in(a0_wr[1806]),  .coef_in(coef[782]), .rdup_out(a1_wr[782]), .rdlo_out(a1_wr[1806]));
			radix2 #(.width(width)) rd_st0_783  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[783]), .rdlo_in(a0_wr[1807]),  .coef_in(coef[783]), .rdup_out(a1_wr[783]), .rdlo_out(a1_wr[1807]));
			radix2 #(.width(width)) rd_st0_784  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[784]), .rdlo_in(a0_wr[1808]),  .coef_in(coef[784]), .rdup_out(a1_wr[784]), .rdlo_out(a1_wr[1808]));
			radix2 #(.width(width)) rd_st0_785  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[785]), .rdlo_in(a0_wr[1809]),  .coef_in(coef[785]), .rdup_out(a1_wr[785]), .rdlo_out(a1_wr[1809]));
			radix2 #(.width(width)) rd_st0_786  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[786]), .rdlo_in(a0_wr[1810]),  .coef_in(coef[786]), .rdup_out(a1_wr[786]), .rdlo_out(a1_wr[1810]));
			radix2 #(.width(width)) rd_st0_787  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[787]), .rdlo_in(a0_wr[1811]),  .coef_in(coef[787]), .rdup_out(a1_wr[787]), .rdlo_out(a1_wr[1811]));
			radix2 #(.width(width)) rd_st0_788  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[788]), .rdlo_in(a0_wr[1812]),  .coef_in(coef[788]), .rdup_out(a1_wr[788]), .rdlo_out(a1_wr[1812]));
			radix2 #(.width(width)) rd_st0_789  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[789]), .rdlo_in(a0_wr[1813]),  .coef_in(coef[789]), .rdup_out(a1_wr[789]), .rdlo_out(a1_wr[1813]));
			radix2 #(.width(width)) rd_st0_790  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[790]), .rdlo_in(a0_wr[1814]),  .coef_in(coef[790]), .rdup_out(a1_wr[790]), .rdlo_out(a1_wr[1814]));
			radix2 #(.width(width)) rd_st0_791  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[791]), .rdlo_in(a0_wr[1815]),  .coef_in(coef[791]), .rdup_out(a1_wr[791]), .rdlo_out(a1_wr[1815]));
			radix2 #(.width(width)) rd_st0_792  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[792]), .rdlo_in(a0_wr[1816]),  .coef_in(coef[792]), .rdup_out(a1_wr[792]), .rdlo_out(a1_wr[1816]));
			radix2 #(.width(width)) rd_st0_793  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[793]), .rdlo_in(a0_wr[1817]),  .coef_in(coef[793]), .rdup_out(a1_wr[793]), .rdlo_out(a1_wr[1817]));
			radix2 #(.width(width)) rd_st0_794  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[794]), .rdlo_in(a0_wr[1818]),  .coef_in(coef[794]), .rdup_out(a1_wr[794]), .rdlo_out(a1_wr[1818]));
			radix2 #(.width(width)) rd_st0_795  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[795]), .rdlo_in(a0_wr[1819]),  .coef_in(coef[795]), .rdup_out(a1_wr[795]), .rdlo_out(a1_wr[1819]));
			radix2 #(.width(width)) rd_st0_796  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[796]), .rdlo_in(a0_wr[1820]),  .coef_in(coef[796]), .rdup_out(a1_wr[796]), .rdlo_out(a1_wr[1820]));
			radix2 #(.width(width)) rd_st0_797  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[797]), .rdlo_in(a0_wr[1821]),  .coef_in(coef[797]), .rdup_out(a1_wr[797]), .rdlo_out(a1_wr[1821]));
			radix2 #(.width(width)) rd_st0_798  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[798]), .rdlo_in(a0_wr[1822]),  .coef_in(coef[798]), .rdup_out(a1_wr[798]), .rdlo_out(a1_wr[1822]));
			radix2 #(.width(width)) rd_st0_799  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[799]), .rdlo_in(a0_wr[1823]),  .coef_in(coef[799]), .rdup_out(a1_wr[799]), .rdlo_out(a1_wr[1823]));
			radix2 #(.width(width)) rd_st0_800  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[800]), .rdlo_in(a0_wr[1824]),  .coef_in(coef[800]), .rdup_out(a1_wr[800]), .rdlo_out(a1_wr[1824]));
			radix2 #(.width(width)) rd_st0_801  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[801]), .rdlo_in(a0_wr[1825]),  .coef_in(coef[801]), .rdup_out(a1_wr[801]), .rdlo_out(a1_wr[1825]));
			radix2 #(.width(width)) rd_st0_802  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[802]), .rdlo_in(a0_wr[1826]),  .coef_in(coef[802]), .rdup_out(a1_wr[802]), .rdlo_out(a1_wr[1826]));
			radix2 #(.width(width)) rd_st0_803  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[803]), .rdlo_in(a0_wr[1827]),  .coef_in(coef[803]), .rdup_out(a1_wr[803]), .rdlo_out(a1_wr[1827]));
			radix2 #(.width(width)) rd_st0_804  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[804]), .rdlo_in(a0_wr[1828]),  .coef_in(coef[804]), .rdup_out(a1_wr[804]), .rdlo_out(a1_wr[1828]));
			radix2 #(.width(width)) rd_st0_805  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[805]), .rdlo_in(a0_wr[1829]),  .coef_in(coef[805]), .rdup_out(a1_wr[805]), .rdlo_out(a1_wr[1829]));
			radix2 #(.width(width)) rd_st0_806  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[806]), .rdlo_in(a0_wr[1830]),  .coef_in(coef[806]), .rdup_out(a1_wr[806]), .rdlo_out(a1_wr[1830]));
			radix2 #(.width(width)) rd_st0_807  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[807]), .rdlo_in(a0_wr[1831]),  .coef_in(coef[807]), .rdup_out(a1_wr[807]), .rdlo_out(a1_wr[1831]));
			radix2 #(.width(width)) rd_st0_808  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[808]), .rdlo_in(a0_wr[1832]),  .coef_in(coef[808]), .rdup_out(a1_wr[808]), .rdlo_out(a1_wr[1832]));
			radix2 #(.width(width)) rd_st0_809  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[809]), .rdlo_in(a0_wr[1833]),  .coef_in(coef[809]), .rdup_out(a1_wr[809]), .rdlo_out(a1_wr[1833]));
			radix2 #(.width(width)) rd_st0_810  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[810]), .rdlo_in(a0_wr[1834]),  .coef_in(coef[810]), .rdup_out(a1_wr[810]), .rdlo_out(a1_wr[1834]));
			radix2 #(.width(width)) rd_st0_811  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[811]), .rdlo_in(a0_wr[1835]),  .coef_in(coef[811]), .rdup_out(a1_wr[811]), .rdlo_out(a1_wr[1835]));
			radix2 #(.width(width)) rd_st0_812  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[812]), .rdlo_in(a0_wr[1836]),  .coef_in(coef[812]), .rdup_out(a1_wr[812]), .rdlo_out(a1_wr[1836]));
			radix2 #(.width(width)) rd_st0_813  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[813]), .rdlo_in(a0_wr[1837]),  .coef_in(coef[813]), .rdup_out(a1_wr[813]), .rdlo_out(a1_wr[1837]));
			radix2 #(.width(width)) rd_st0_814  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[814]), .rdlo_in(a0_wr[1838]),  .coef_in(coef[814]), .rdup_out(a1_wr[814]), .rdlo_out(a1_wr[1838]));
			radix2 #(.width(width)) rd_st0_815  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[815]), .rdlo_in(a0_wr[1839]),  .coef_in(coef[815]), .rdup_out(a1_wr[815]), .rdlo_out(a1_wr[1839]));
			radix2 #(.width(width)) rd_st0_816  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[816]), .rdlo_in(a0_wr[1840]),  .coef_in(coef[816]), .rdup_out(a1_wr[816]), .rdlo_out(a1_wr[1840]));
			radix2 #(.width(width)) rd_st0_817  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[817]), .rdlo_in(a0_wr[1841]),  .coef_in(coef[817]), .rdup_out(a1_wr[817]), .rdlo_out(a1_wr[1841]));
			radix2 #(.width(width)) rd_st0_818  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[818]), .rdlo_in(a0_wr[1842]),  .coef_in(coef[818]), .rdup_out(a1_wr[818]), .rdlo_out(a1_wr[1842]));
			radix2 #(.width(width)) rd_st0_819  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[819]), .rdlo_in(a0_wr[1843]),  .coef_in(coef[819]), .rdup_out(a1_wr[819]), .rdlo_out(a1_wr[1843]));
			radix2 #(.width(width)) rd_st0_820  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[820]), .rdlo_in(a0_wr[1844]),  .coef_in(coef[820]), .rdup_out(a1_wr[820]), .rdlo_out(a1_wr[1844]));
			radix2 #(.width(width)) rd_st0_821  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[821]), .rdlo_in(a0_wr[1845]),  .coef_in(coef[821]), .rdup_out(a1_wr[821]), .rdlo_out(a1_wr[1845]));
			radix2 #(.width(width)) rd_st0_822  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[822]), .rdlo_in(a0_wr[1846]),  .coef_in(coef[822]), .rdup_out(a1_wr[822]), .rdlo_out(a1_wr[1846]));
			radix2 #(.width(width)) rd_st0_823  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[823]), .rdlo_in(a0_wr[1847]),  .coef_in(coef[823]), .rdup_out(a1_wr[823]), .rdlo_out(a1_wr[1847]));
			radix2 #(.width(width)) rd_st0_824  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[824]), .rdlo_in(a0_wr[1848]),  .coef_in(coef[824]), .rdup_out(a1_wr[824]), .rdlo_out(a1_wr[1848]));
			radix2 #(.width(width)) rd_st0_825  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[825]), .rdlo_in(a0_wr[1849]),  .coef_in(coef[825]), .rdup_out(a1_wr[825]), .rdlo_out(a1_wr[1849]));
			radix2 #(.width(width)) rd_st0_826  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[826]), .rdlo_in(a0_wr[1850]),  .coef_in(coef[826]), .rdup_out(a1_wr[826]), .rdlo_out(a1_wr[1850]));
			radix2 #(.width(width)) rd_st0_827  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[827]), .rdlo_in(a0_wr[1851]),  .coef_in(coef[827]), .rdup_out(a1_wr[827]), .rdlo_out(a1_wr[1851]));
			radix2 #(.width(width)) rd_st0_828  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[828]), .rdlo_in(a0_wr[1852]),  .coef_in(coef[828]), .rdup_out(a1_wr[828]), .rdlo_out(a1_wr[1852]));
			radix2 #(.width(width)) rd_st0_829  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[829]), .rdlo_in(a0_wr[1853]),  .coef_in(coef[829]), .rdup_out(a1_wr[829]), .rdlo_out(a1_wr[1853]));
			radix2 #(.width(width)) rd_st0_830  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[830]), .rdlo_in(a0_wr[1854]),  .coef_in(coef[830]), .rdup_out(a1_wr[830]), .rdlo_out(a1_wr[1854]));
			radix2 #(.width(width)) rd_st0_831  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[831]), .rdlo_in(a0_wr[1855]),  .coef_in(coef[831]), .rdup_out(a1_wr[831]), .rdlo_out(a1_wr[1855]));
			radix2 #(.width(width)) rd_st0_832  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[832]), .rdlo_in(a0_wr[1856]),  .coef_in(coef[832]), .rdup_out(a1_wr[832]), .rdlo_out(a1_wr[1856]));
			radix2 #(.width(width)) rd_st0_833  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[833]), .rdlo_in(a0_wr[1857]),  .coef_in(coef[833]), .rdup_out(a1_wr[833]), .rdlo_out(a1_wr[1857]));
			radix2 #(.width(width)) rd_st0_834  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[834]), .rdlo_in(a0_wr[1858]),  .coef_in(coef[834]), .rdup_out(a1_wr[834]), .rdlo_out(a1_wr[1858]));
			radix2 #(.width(width)) rd_st0_835  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[835]), .rdlo_in(a0_wr[1859]),  .coef_in(coef[835]), .rdup_out(a1_wr[835]), .rdlo_out(a1_wr[1859]));
			radix2 #(.width(width)) rd_st0_836  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[836]), .rdlo_in(a0_wr[1860]),  .coef_in(coef[836]), .rdup_out(a1_wr[836]), .rdlo_out(a1_wr[1860]));
			radix2 #(.width(width)) rd_st0_837  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[837]), .rdlo_in(a0_wr[1861]),  .coef_in(coef[837]), .rdup_out(a1_wr[837]), .rdlo_out(a1_wr[1861]));
			radix2 #(.width(width)) rd_st0_838  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[838]), .rdlo_in(a0_wr[1862]),  .coef_in(coef[838]), .rdup_out(a1_wr[838]), .rdlo_out(a1_wr[1862]));
			radix2 #(.width(width)) rd_st0_839  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[839]), .rdlo_in(a0_wr[1863]),  .coef_in(coef[839]), .rdup_out(a1_wr[839]), .rdlo_out(a1_wr[1863]));
			radix2 #(.width(width)) rd_st0_840  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[840]), .rdlo_in(a0_wr[1864]),  .coef_in(coef[840]), .rdup_out(a1_wr[840]), .rdlo_out(a1_wr[1864]));
			radix2 #(.width(width)) rd_st0_841  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[841]), .rdlo_in(a0_wr[1865]),  .coef_in(coef[841]), .rdup_out(a1_wr[841]), .rdlo_out(a1_wr[1865]));
			radix2 #(.width(width)) rd_st0_842  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[842]), .rdlo_in(a0_wr[1866]),  .coef_in(coef[842]), .rdup_out(a1_wr[842]), .rdlo_out(a1_wr[1866]));
			radix2 #(.width(width)) rd_st0_843  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[843]), .rdlo_in(a0_wr[1867]),  .coef_in(coef[843]), .rdup_out(a1_wr[843]), .rdlo_out(a1_wr[1867]));
			radix2 #(.width(width)) rd_st0_844  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[844]), .rdlo_in(a0_wr[1868]),  .coef_in(coef[844]), .rdup_out(a1_wr[844]), .rdlo_out(a1_wr[1868]));
			radix2 #(.width(width)) rd_st0_845  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[845]), .rdlo_in(a0_wr[1869]),  .coef_in(coef[845]), .rdup_out(a1_wr[845]), .rdlo_out(a1_wr[1869]));
			radix2 #(.width(width)) rd_st0_846  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[846]), .rdlo_in(a0_wr[1870]),  .coef_in(coef[846]), .rdup_out(a1_wr[846]), .rdlo_out(a1_wr[1870]));
			radix2 #(.width(width)) rd_st0_847  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[847]), .rdlo_in(a0_wr[1871]),  .coef_in(coef[847]), .rdup_out(a1_wr[847]), .rdlo_out(a1_wr[1871]));
			radix2 #(.width(width)) rd_st0_848  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[848]), .rdlo_in(a0_wr[1872]),  .coef_in(coef[848]), .rdup_out(a1_wr[848]), .rdlo_out(a1_wr[1872]));
			radix2 #(.width(width)) rd_st0_849  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[849]), .rdlo_in(a0_wr[1873]),  .coef_in(coef[849]), .rdup_out(a1_wr[849]), .rdlo_out(a1_wr[1873]));
			radix2 #(.width(width)) rd_st0_850  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[850]), .rdlo_in(a0_wr[1874]),  .coef_in(coef[850]), .rdup_out(a1_wr[850]), .rdlo_out(a1_wr[1874]));
			radix2 #(.width(width)) rd_st0_851  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[851]), .rdlo_in(a0_wr[1875]),  .coef_in(coef[851]), .rdup_out(a1_wr[851]), .rdlo_out(a1_wr[1875]));
			radix2 #(.width(width)) rd_st0_852  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[852]), .rdlo_in(a0_wr[1876]),  .coef_in(coef[852]), .rdup_out(a1_wr[852]), .rdlo_out(a1_wr[1876]));
			radix2 #(.width(width)) rd_st0_853  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[853]), .rdlo_in(a0_wr[1877]),  .coef_in(coef[853]), .rdup_out(a1_wr[853]), .rdlo_out(a1_wr[1877]));
			radix2 #(.width(width)) rd_st0_854  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[854]), .rdlo_in(a0_wr[1878]),  .coef_in(coef[854]), .rdup_out(a1_wr[854]), .rdlo_out(a1_wr[1878]));
			radix2 #(.width(width)) rd_st0_855  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[855]), .rdlo_in(a0_wr[1879]),  .coef_in(coef[855]), .rdup_out(a1_wr[855]), .rdlo_out(a1_wr[1879]));
			radix2 #(.width(width)) rd_st0_856  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[856]), .rdlo_in(a0_wr[1880]),  .coef_in(coef[856]), .rdup_out(a1_wr[856]), .rdlo_out(a1_wr[1880]));
			radix2 #(.width(width)) rd_st0_857  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[857]), .rdlo_in(a0_wr[1881]),  .coef_in(coef[857]), .rdup_out(a1_wr[857]), .rdlo_out(a1_wr[1881]));
			radix2 #(.width(width)) rd_st0_858  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[858]), .rdlo_in(a0_wr[1882]),  .coef_in(coef[858]), .rdup_out(a1_wr[858]), .rdlo_out(a1_wr[1882]));
			radix2 #(.width(width)) rd_st0_859  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[859]), .rdlo_in(a0_wr[1883]),  .coef_in(coef[859]), .rdup_out(a1_wr[859]), .rdlo_out(a1_wr[1883]));
			radix2 #(.width(width)) rd_st0_860  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[860]), .rdlo_in(a0_wr[1884]),  .coef_in(coef[860]), .rdup_out(a1_wr[860]), .rdlo_out(a1_wr[1884]));
			radix2 #(.width(width)) rd_st0_861  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[861]), .rdlo_in(a0_wr[1885]),  .coef_in(coef[861]), .rdup_out(a1_wr[861]), .rdlo_out(a1_wr[1885]));
			radix2 #(.width(width)) rd_st0_862  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[862]), .rdlo_in(a0_wr[1886]),  .coef_in(coef[862]), .rdup_out(a1_wr[862]), .rdlo_out(a1_wr[1886]));
			radix2 #(.width(width)) rd_st0_863  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[863]), .rdlo_in(a0_wr[1887]),  .coef_in(coef[863]), .rdup_out(a1_wr[863]), .rdlo_out(a1_wr[1887]));
			radix2 #(.width(width)) rd_st0_864  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[864]), .rdlo_in(a0_wr[1888]),  .coef_in(coef[864]), .rdup_out(a1_wr[864]), .rdlo_out(a1_wr[1888]));
			radix2 #(.width(width)) rd_st0_865  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[865]), .rdlo_in(a0_wr[1889]),  .coef_in(coef[865]), .rdup_out(a1_wr[865]), .rdlo_out(a1_wr[1889]));
			radix2 #(.width(width)) rd_st0_866  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[866]), .rdlo_in(a0_wr[1890]),  .coef_in(coef[866]), .rdup_out(a1_wr[866]), .rdlo_out(a1_wr[1890]));
			radix2 #(.width(width)) rd_st0_867  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[867]), .rdlo_in(a0_wr[1891]),  .coef_in(coef[867]), .rdup_out(a1_wr[867]), .rdlo_out(a1_wr[1891]));
			radix2 #(.width(width)) rd_st0_868  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[868]), .rdlo_in(a0_wr[1892]),  .coef_in(coef[868]), .rdup_out(a1_wr[868]), .rdlo_out(a1_wr[1892]));
			radix2 #(.width(width)) rd_st0_869  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[869]), .rdlo_in(a0_wr[1893]),  .coef_in(coef[869]), .rdup_out(a1_wr[869]), .rdlo_out(a1_wr[1893]));
			radix2 #(.width(width)) rd_st0_870  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[870]), .rdlo_in(a0_wr[1894]),  .coef_in(coef[870]), .rdup_out(a1_wr[870]), .rdlo_out(a1_wr[1894]));
			radix2 #(.width(width)) rd_st0_871  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[871]), .rdlo_in(a0_wr[1895]),  .coef_in(coef[871]), .rdup_out(a1_wr[871]), .rdlo_out(a1_wr[1895]));
			radix2 #(.width(width)) rd_st0_872  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[872]), .rdlo_in(a0_wr[1896]),  .coef_in(coef[872]), .rdup_out(a1_wr[872]), .rdlo_out(a1_wr[1896]));
			radix2 #(.width(width)) rd_st0_873  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[873]), .rdlo_in(a0_wr[1897]),  .coef_in(coef[873]), .rdup_out(a1_wr[873]), .rdlo_out(a1_wr[1897]));
			radix2 #(.width(width)) rd_st0_874  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[874]), .rdlo_in(a0_wr[1898]),  .coef_in(coef[874]), .rdup_out(a1_wr[874]), .rdlo_out(a1_wr[1898]));
			radix2 #(.width(width)) rd_st0_875  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[875]), .rdlo_in(a0_wr[1899]),  .coef_in(coef[875]), .rdup_out(a1_wr[875]), .rdlo_out(a1_wr[1899]));
			radix2 #(.width(width)) rd_st0_876  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[876]), .rdlo_in(a0_wr[1900]),  .coef_in(coef[876]), .rdup_out(a1_wr[876]), .rdlo_out(a1_wr[1900]));
			radix2 #(.width(width)) rd_st0_877  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[877]), .rdlo_in(a0_wr[1901]),  .coef_in(coef[877]), .rdup_out(a1_wr[877]), .rdlo_out(a1_wr[1901]));
			radix2 #(.width(width)) rd_st0_878  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[878]), .rdlo_in(a0_wr[1902]),  .coef_in(coef[878]), .rdup_out(a1_wr[878]), .rdlo_out(a1_wr[1902]));
			radix2 #(.width(width)) rd_st0_879  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[879]), .rdlo_in(a0_wr[1903]),  .coef_in(coef[879]), .rdup_out(a1_wr[879]), .rdlo_out(a1_wr[1903]));
			radix2 #(.width(width)) rd_st0_880  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[880]), .rdlo_in(a0_wr[1904]),  .coef_in(coef[880]), .rdup_out(a1_wr[880]), .rdlo_out(a1_wr[1904]));
			radix2 #(.width(width)) rd_st0_881  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[881]), .rdlo_in(a0_wr[1905]),  .coef_in(coef[881]), .rdup_out(a1_wr[881]), .rdlo_out(a1_wr[1905]));
			radix2 #(.width(width)) rd_st0_882  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[882]), .rdlo_in(a0_wr[1906]),  .coef_in(coef[882]), .rdup_out(a1_wr[882]), .rdlo_out(a1_wr[1906]));
			radix2 #(.width(width)) rd_st0_883  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[883]), .rdlo_in(a0_wr[1907]),  .coef_in(coef[883]), .rdup_out(a1_wr[883]), .rdlo_out(a1_wr[1907]));
			radix2 #(.width(width)) rd_st0_884  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[884]), .rdlo_in(a0_wr[1908]),  .coef_in(coef[884]), .rdup_out(a1_wr[884]), .rdlo_out(a1_wr[1908]));
			radix2 #(.width(width)) rd_st0_885  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[885]), .rdlo_in(a0_wr[1909]),  .coef_in(coef[885]), .rdup_out(a1_wr[885]), .rdlo_out(a1_wr[1909]));
			radix2 #(.width(width)) rd_st0_886  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[886]), .rdlo_in(a0_wr[1910]),  .coef_in(coef[886]), .rdup_out(a1_wr[886]), .rdlo_out(a1_wr[1910]));
			radix2 #(.width(width)) rd_st0_887  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[887]), .rdlo_in(a0_wr[1911]),  .coef_in(coef[887]), .rdup_out(a1_wr[887]), .rdlo_out(a1_wr[1911]));
			radix2 #(.width(width)) rd_st0_888  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[888]), .rdlo_in(a0_wr[1912]),  .coef_in(coef[888]), .rdup_out(a1_wr[888]), .rdlo_out(a1_wr[1912]));
			radix2 #(.width(width)) rd_st0_889  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[889]), .rdlo_in(a0_wr[1913]),  .coef_in(coef[889]), .rdup_out(a1_wr[889]), .rdlo_out(a1_wr[1913]));
			radix2 #(.width(width)) rd_st0_890  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[890]), .rdlo_in(a0_wr[1914]),  .coef_in(coef[890]), .rdup_out(a1_wr[890]), .rdlo_out(a1_wr[1914]));
			radix2 #(.width(width)) rd_st0_891  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[891]), .rdlo_in(a0_wr[1915]),  .coef_in(coef[891]), .rdup_out(a1_wr[891]), .rdlo_out(a1_wr[1915]));
			radix2 #(.width(width)) rd_st0_892  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[892]), .rdlo_in(a0_wr[1916]),  .coef_in(coef[892]), .rdup_out(a1_wr[892]), .rdlo_out(a1_wr[1916]));
			radix2 #(.width(width)) rd_st0_893  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[893]), .rdlo_in(a0_wr[1917]),  .coef_in(coef[893]), .rdup_out(a1_wr[893]), .rdlo_out(a1_wr[1917]));
			radix2 #(.width(width)) rd_st0_894  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[894]), .rdlo_in(a0_wr[1918]),  .coef_in(coef[894]), .rdup_out(a1_wr[894]), .rdlo_out(a1_wr[1918]));
			radix2 #(.width(width)) rd_st0_895  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[895]), .rdlo_in(a0_wr[1919]),  .coef_in(coef[895]), .rdup_out(a1_wr[895]), .rdlo_out(a1_wr[1919]));
			radix2 #(.width(width)) rd_st0_896  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[896]), .rdlo_in(a0_wr[1920]),  .coef_in(coef[896]), .rdup_out(a1_wr[896]), .rdlo_out(a1_wr[1920]));
			radix2 #(.width(width)) rd_st0_897  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[897]), .rdlo_in(a0_wr[1921]),  .coef_in(coef[897]), .rdup_out(a1_wr[897]), .rdlo_out(a1_wr[1921]));
			radix2 #(.width(width)) rd_st0_898  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[898]), .rdlo_in(a0_wr[1922]),  .coef_in(coef[898]), .rdup_out(a1_wr[898]), .rdlo_out(a1_wr[1922]));
			radix2 #(.width(width)) rd_st0_899  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[899]), .rdlo_in(a0_wr[1923]),  .coef_in(coef[899]), .rdup_out(a1_wr[899]), .rdlo_out(a1_wr[1923]));
			radix2 #(.width(width)) rd_st0_900  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[900]), .rdlo_in(a0_wr[1924]),  .coef_in(coef[900]), .rdup_out(a1_wr[900]), .rdlo_out(a1_wr[1924]));
			radix2 #(.width(width)) rd_st0_901  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[901]), .rdlo_in(a0_wr[1925]),  .coef_in(coef[901]), .rdup_out(a1_wr[901]), .rdlo_out(a1_wr[1925]));
			radix2 #(.width(width)) rd_st0_902  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[902]), .rdlo_in(a0_wr[1926]),  .coef_in(coef[902]), .rdup_out(a1_wr[902]), .rdlo_out(a1_wr[1926]));
			radix2 #(.width(width)) rd_st0_903  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[903]), .rdlo_in(a0_wr[1927]),  .coef_in(coef[903]), .rdup_out(a1_wr[903]), .rdlo_out(a1_wr[1927]));
			radix2 #(.width(width)) rd_st0_904  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[904]), .rdlo_in(a0_wr[1928]),  .coef_in(coef[904]), .rdup_out(a1_wr[904]), .rdlo_out(a1_wr[1928]));
			radix2 #(.width(width)) rd_st0_905  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[905]), .rdlo_in(a0_wr[1929]),  .coef_in(coef[905]), .rdup_out(a1_wr[905]), .rdlo_out(a1_wr[1929]));
			radix2 #(.width(width)) rd_st0_906  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[906]), .rdlo_in(a0_wr[1930]),  .coef_in(coef[906]), .rdup_out(a1_wr[906]), .rdlo_out(a1_wr[1930]));
			radix2 #(.width(width)) rd_st0_907  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[907]), .rdlo_in(a0_wr[1931]),  .coef_in(coef[907]), .rdup_out(a1_wr[907]), .rdlo_out(a1_wr[1931]));
			radix2 #(.width(width)) rd_st0_908  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[908]), .rdlo_in(a0_wr[1932]),  .coef_in(coef[908]), .rdup_out(a1_wr[908]), .rdlo_out(a1_wr[1932]));
			radix2 #(.width(width)) rd_st0_909  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[909]), .rdlo_in(a0_wr[1933]),  .coef_in(coef[909]), .rdup_out(a1_wr[909]), .rdlo_out(a1_wr[1933]));
			radix2 #(.width(width)) rd_st0_910  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[910]), .rdlo_in(a0_wr[1934]),  .coef_in(coef[910]), .rdup_out(a1_wr[910]), .rdlo_out(a1_wr[1934]));
			radix2 #(.width(width)) rd_st0_911  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[911]), .rdlo_in(a0_wr[1935]),  .coef_in(coef[911]), .rdup_out(a1_wr[911]), .rdlo_out(a1_wr[1935]));
			radix2 #(.width(width)) rd_st0_912  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[912]), .rdlo_in(a0_wr[1936]),  .coef_in(coef[912]), .rdup_out(a1_wr[912]), .rdlo_out(a1_wr[1936]));
			radix2 #(.width(width)) rd_st0_913  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[913]), .rdlo_in(a0_wr[1937]),  .coef_in(coef[913]), .rdup_out(a1_wr[913]), .rdlo_out(a1_wr[1937]));
			radix2 #(.width(width)) rd_st0_914  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[914]), .rdlo_in(a0_wr[1938]),  .coef_in(coef[914]), .rdup_out(a1_wr[914]), .rdlo_out(a1_wr[1938]));
			radix2 #(.width(width)) rd_st0_915  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[915]), .rdlo_in(a0_wr[1939]),  .coef_in(coef[915]), .rdup_out(a1_wr[915]), .rdlo_out(a1_wr[1939]));
			radix2 #(.width(width)) rd_st0_916  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[916]), .rdlo_in(a0_wr[1940]),  .coef_in(coef[916]), .rdup_out(a1_wr[916]), .rdlo_out(a1_wr[1940]));
			radix2 #(.width(width)) rd_st0_917  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[917]), .rdlo_in(a0_wr[1941]),  .coef_in(coef[917]), .rdup_out(a1_wr[917]), .rdlo_out(a1_wr[1941]));
			radix2 #(.width(width)) rd_st0_918  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[918]), .rdlo_in(a0_wr[1942]),  .coef_in(coef[918]), .rdup_out(a1_wr[918]), .rdlo_out(a1_wr[1942]));
			radix2 #(.width(width)) rd_st0_919  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[919]), .rdlo_in(a0_wr[1943]),  .coef_in(coef[919]), .rdup_out(a1_wr[919]), .rdlo_out(a1_wr[1943]));
			radix2 #(.width(width)) rd_st0_920  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[920]), .rdlo_in(a0_wr[1944]),  .coef_in(coef[920]), .rdup_out(a1_wr[920]), .rdlo_out(a1_wr[1944]));
			radix2 #(.width(width)) rd_st0_921  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[921]), .rdlo_in(a0_wr[1945]),  .coef_in(coef[921]), .rdup_out(a1_wr[921]), .rdlo_out(a1_wr[1945]));
			radix2 #(.width(width)) rd_st0_922  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[922]), .rdlo_in(a0_wr[1946]),  .coef_in(coef[922]), .rdup_out(a1_wr[922]), .rdlo_out(a1_wr[1946]));
			radix2 #(.width(width)) rd_st0_923  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[923]), .rdlo_in(a0_wr[1947]),  .coef_in(coef[923]), .rdup_out(a1_wr[923]), .rdlo_out(a1_wr[1947]));
			radix2 #(.width(width)) rd_st0_924  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[924]), .rdlo_in(a0_wr[1948]),  .coef_in(coef[924]), .rdup_out(a1_wr[924]), .rdlo_out(a1_wr[1948]));
			radix2 #(.width(width)) rd_st0_925  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[925]), .rdlo_in(a0_wr[1949]),  .coef_in(coef[925]), .rdup_out(a1_wr[925]), .rdlo_out(a1_wr[1949]));
			radix2 #(.width(width)) rd_st0_926  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[926]), .rdlo_in(a0_wr[1950]),  .coef_in(coef[926]), .rdup_out(a1_wr[926]), .rdlo_out(a1_wr[1950]));
			radix2 #(.width(width)) rd_st0_927  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[927]), .rdlo_in(a0_wr[1951]),  .coef_in(coef[927]), .rdup_out(a1_wr[927]), .rdlo_out(a1_wr[1951]));
			radix2 #(.width(width)) rd_st0_928  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[928]), .rdlo_in(a0_wr[1952]),  .coef_in(coef[928]), .rdup_out(a1_wr[928]), .rdlo_out(a1_wr[1952]));
			radix2 #(.width(width)) rd_st0_929  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[929]), .rdlo_in(a0_wr[1953]),  .coef_in(coef[929]), .rdup_out(a1_wr[929]), .rdlo_out(a1_wr[1953]));
			radix2 #(.width(width)) rd_st0_930  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[930]), .rdlo_in(a0_wr[1954]),  .coef_in(coef[930]), .rdup_out(a1_wr[930]), .rdlo_out(a1_wr[1954]));
			radix2 #(.width(width)) rd_st0_931  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[931]), .rdlo_in(a0_wr[1955]),  .coef_in(coef[931]), .rdup_out(a1_wr[931]), .rdlo_out(a1_wr[1955]));
			radix2 #(.width(width)) rd_st0_932  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[932]), .rdlo_in(a0_wr[1956]),  .coef_in(coef[932]), .rdup_out(a1_wr[932]), .rdlo_out(a1_wr[1956]));
			radix2 #(.width(width)) rd_st0_933  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[933]), .rdlo_in(a0_wr[1957]),  .coef_in(coef[933]), .rdup_out(a1_wr[933]), .rdlo_out(a1_wr[1957]));
			radix2 #(.width(width)) rd_st0_934  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[934]), .rdlo_in(a0_wr[1958]),  .coef_in(coef[934]), .rdup_out(a1_wr[934]), .rdlo_out(a1_wr[1958]));
			radix2 #(.width(width)) rd_st0_935  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[935]), .rdlo_in(a0_wr[1959]),  .coef_in(coef[935]), .rdup_out(a1_wr[935]), .rdlo_out(a1_wr[1959]));
			radix2 #(.width(width)) rd_st0_936  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[936]), .rdlo_in(a0_wr[1960]),  .coef_in(coef[936]), .rdup_out(a1_wr[936]), .rdlo_out(a1_wr[1960]));
			radix2 #(.width(width)) rd_st0_937  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[937]), .rdlo_in(a0_wr[1961]),  .coef_in(coef[937]), .rdup_out(a1_wr[937]), .rdlo_out(a1_wr[1961]));
			radix2 #(.width(width)) rd_st0_938  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[938]), .rdlo_in(a0_wr[1962]),  .coef_in(coef[938]), .rdup_out(a1_wr[938]), .rdlo_out(a1_wr[1962]));
			radix2 #(.width(width)) rd_st0_939  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[939]), .rdlo_in(a0_wr[1963]),  .coef_in(coef[939]), .rdup_out(a1_wr[939]), .rdlo_out(a1_wr[1963]));
			radix2 #(.width(width)) rd_st0_940  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[940]), .rdlo_in(a0_wr[1964]),  .coef_in(coef[940]), .rdup_out(a1_wr[940]), .rdlo_out(a1_wr[1964]));
			radix2 #(.width(width)) rd_st0_941  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[941]), .rdlo_in(a0_wr[1965]),  .coef_in(coef[941]), .rdup_out(a1_wr[941]), .rdlo_out(a1_wr[1965]));
			radix2 #(.width(width)) rd_st0_942  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[942]), .rdlo_in(a0_wr[1966]),  .coef_in(coef[942]), .rdup_out(a1_wr[942]), .rdlo_out(a1_wr[1966]));
			radix2 #(.width(width)) rd_st0_943  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[943]), .rdlo_in(a0_wr[1967]),  .coef_in(coef[943]), .rdup_out(a1_wr[943]), .rdlo_out(a1_wr[1967]));
			radix2 #(.width(width)) rd_st0_944  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[944]), .rdlo_in(a0_wr[1968]),  .coef_in(coef[944]), .rdup_out(a1_wr[944]), .rdlo_out(a1_wr[1968]));
			radix2 #(.width(width)) rd_st0_945  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[945]), .rdlo_in(a0_wr[1969]),  .coef_in(coef[945]), .rdup_out(a1_wr[945]), .rdlo_out(a1_wr[1969]));
			radix2 #(.width(width)) rd_st0_946  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[946]), .rdlo_in(a0_wr[1970]),  .coef_in(coef[946]), .rdup_out(a1_wr[946]), .rdlo_out(a1_wr[1970]));
			radix2 #(.width(width)) rd_st0_947  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[947]), .rdlo_in(a0_wr[1971]),  .coef_in(coef[947]), .rdup_out(a1_wr[947]), .rdlo_out(a1_wr[1971]));
			radix2 #(.width(width)) rd_st0_948  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[948]), .rdlo_in(a0_wr[1972]),  .coef_in(coef[948]), .rdup_out(a1_wr[948]), .rdlo_out(a1_wr[1972]));
			radix2 #(.width(width)) rd_st0_949  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[949]), .rdlo_in(a0_wr[1973]),  .coef_in(coef[949]), .rdup_out(a1_wr[949]), .rdlo_out(a1_wr[1973]));
			radix2 #(.width(width)) rd_st0_950  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[950]), .rdlo_in(a0_wr[1974]),  .coef_in(coef[950]), .rdup_out(a1_wr[950]), .rdlo_out(a1_wr[1974]));
			radix2 #(.width(width)) rd_st0_951  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[951]), .rdlo_in(a0_wr[1975]),  .coef_in(coef[951]), .rdup_out(a1_wr[951]), .rdlo_out(a1_wr[1975]));
			radix2 #(.width(width)) rd_st0_952  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[952]), .rdlo_in(a0_wr[1976]),  .coef_in(coef[952]), .rdup_out(a1_wr[952]), .rdlo_out(a1_wr[1976]));
			radix2 #(.width(width)) rd_st0_953  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[953]), .rdlo_in(a0_wr[1977]),  .coef_in(coef[953]), .rdup_out(a1_wr[953]), .rdlo_out(a1_wr[1977]));
			radix2 #(.width(width)) rd_st0_954  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[954]), .rdlo_in(a0_wr[1978]),  .coef_in(coef[954]), .rdup_out(a1_wr[954]), .rdlo_out(a1_wr[1978]));
			radix2 #(.width(width)) rd_st0_955  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[955]), .rdlo_in(a0_wr[1979]),  .coef_in(coef[955]), .rdup_out(a1_wr[955]), .rdlo_out(a1_wr[1979]));
			radix2 #(.width(width)) rd_st0_956  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[956]), .rdlo_in(a0_wr[1980]),  .coef_in(coef[956]), .rdup_out(a1_wr[956]), .rdlo_out(a1_wr[1980]));
			radix2 #(.width(width)) rd_st0_957  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[957]), .rdlo_in(a0_wr[1981]),  .coef_in(coef[957]), .rdup_out(a1_wr[957]), .rdlo_out(a1_wr[1981]));
			radix2 #(.width(width)) rd_st0_958  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[958]), .rdlo_in(a0_wr[1982]),  .coef_in(coef[958]), .rdup_out(a1_wr[958]), .rdlo_out(a1_wr[1982]));
			radix2 #(.width(width)) rd_st0_959  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[959]), .rdlo_in(a0_wr[1983]),  .coef_in(coef[959]), .rdup_out(a1_wr[959]), .rdlo_out(a1_wr[1983]));
			radix2 #(.width(width)) rd_st0_960  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[960]), .rdlo_in(a0_wr[1984]),  .coef_in(coef[960]), .rdup_out(a1_wr[960]), .rdlo_out(a1_wr[1984]));
			radix2 #(.width(width)) rd_st0_961  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[961]), .rdlo_in(a0_wr[1985]),  .coef_in(coef[961]), .rdup_out(a1_wr[961]), .rdlo_out(a1_wr[1985]));
			radix2 #(.width(width)) rd_st0_962  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[962]), .rdlo_in(a0_wr[1986]),  .coef_in(coef[962]), .rdup_out(a1_wr[962]), .rdlo_out(a1_wr[1986]));
			radix2 #(.width(width)) rd_st0_963  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[963]), .rdlo_in(a0_wr[1987]),  .coef_in(coef[963]), .rdup_out(a1_wr[963]), .rdlo_out(a1_wr[1987]));
			radix2 #(.width(width)) rd_st0_964  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[964]), .rdlo_in(a0_wr[1988]),  .coef_in(coef[964]), .rdup_out(a1_wr[964]), .rdlo_out(a1_wr[1988]));
			radix2 #(.width(width)) rd_st0_965  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[965]), .rdlo_in(a0_wr[1989]),  .coef_in(coef[965]), .rdup_out(a1_wr[965]), .rdlo_out(a1_wr[1989]));
			radix2 #(.width(width)) rd_st0_966  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[966]), .rdlo_in(a0_wr[1990]),  .coef_in(coef[966]), .rdup_out(a1_wr[966]), .rdlo_out(a1_wr[1990]));
			radix2 #(.width(width)) rd_st0_967  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[967]), .rdlo_in(a0_wr[1991]),  .coef_in(coef[967]), .rdup_out(a1_wr[967]), .rdlo_out(a1_wr[1991]));
			radix2 #(.width(width)) rd_st0_968  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[968]), .rdlo_in(a0_wr[1992]),  .coef_in(coef[968]), .rdup_out(a1_wr[968]), .rdlo_out(a1_wr[1992]));
			radix2 #(.width(width)) rd_st0_969  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[969]), .rdlo_in(a0_wr[1993]),  .coef_in(coef[969]), .rdup_out(a1_wr[969]), .rdlo_out(a1_wr[1993]));
			radix2 #(.width(width)) rd_st0_970  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[970]), .rdlo_in(a0_wr[1994]),  .coef_in(coef[970]), .rdup_out(a1_wr[970]), .rdlo_out(a1_wr[1994]));
			radix2 #(.width(width)) rd_st0_971  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[971]), .rdlo_in(a0_wr[1995]),  .coef_in(coef[971]), .rdup_out(a1_wr[971]), .rdlo_out(a1_wr[1995]));
			radix2 #(.width(width)) rd_st0_972  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[972]), .rdlo_in(a0_wr[1996]),  .coef_in(coef[972]), .rdup_out(a1_wr[972]), .rdlo_out(a1_wr[1996]));
			radix2 #(.width(width)) rd_st0_973  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[973]), .rdlo_in(a0_wr[1997]),  .coef_in(coef[973]), .rdup_out(a1_wr[973]), .rdlo_out(a1_wr[1997]));
			radix2 #(.width(width)) rd_st0_974  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[974]), .rdlo_in(a0_wr[1998]),  .coef_in(coef[974]), .rdup_out(a1_wr[974]), .rdlo_out(a1_wr[1998]));
			radix2 #(.width(width)) rd_st0_975  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[975]), .rdlo_in(a0_wr[1999]),  .coef_in(coef[975]), .rdup_out(a1_wr[975]), .rdlo_out(a1_wr[1999]));
			radix2 #(.width(width)) rd_st0_976  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[976]), .rdlo_in(a0_wr[2000]),  .coef_in(coef[976]), .rdup_out(a1_wr[976]), .rdlo_out(a1_wr[2000]));
			radix2 #(.width(width)) rd_st0_977  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[977]), .rdlo_in(a0_wr[2001]),  .coef_in(coef[977]), .rdup_out(a1_wr[977]), .rdlo_out(a1_wr[2001]));
			radix2 #(.width(width)) rd_st0_978  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[978]), .rdlo_in(a0_wr[2002]),  .coef_in(coef[978]), .rdup_out(a1_wr[978]), .rdlo_out(a1_wr[2002]));
			radix2 #(.width(width)) rd_st0_979  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[979]), .rdlo_in(a0_wr[2003]),  .coef_in(coef[979]), .rdup_out(a1_wr[979]), .rdlo_out(a1_wr[2003]));
			radix2 #(.width(width)) rd_st0_980  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[980]), .rdlo_in(a0_wr[2004]),  .coef_in(coef[980]), .rdup_out(a1_wr[980]), .rdlo_out(a1_wr[2004]));
			radix2 #(.width(width)) rd_st0_981  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[981]), .rdlo_in(a0_wr[2005]),  .coef_in(coef[981]), .rdup_out(a1_wr[981]), .rdlo_out(a1_wr[2005]));
			radix2 #(.width(width)) rd_st0_982  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[982]), .rdlo_in(a0_wr[2006]),  .coef_in(coef[982]), .rdup_out(a1_wr[982]), .rdlo_out(a1_wr[2006]));
			radix2 #(.width(width)) rd_st0_983  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[983]), .rdlo_in(a0_wr[2007]),  .coef_in(coef[983]), .rdup_out(a1_wr[983]), .rdlo_out(a1_wr[2007]));
			radix2 #(.width(width)) rd_st0_984  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[984]), .rdlo_in(a0_wr[2008]),  .coef_in(coef[984]), .rdup_out(a1_wr[984]), .rdlo_out(a1_wr[2008]));
			radix2 #(.width(width)) rd_st0_985  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[985]), .rdlo_in(a0_wr[2009]),  .coef_in(coef[985]), .rdup_out(a1_wr[985]), .rdlo_out(a1_wr[2009]));
			radix2 #(.width(width)) rd_st0_986  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[986]), .rdlo_in(a0_wr[2010]),  .coef_in(coef[986]), .rdup_out(a1_wr[986]), .rdlo_out(a1_wr[2010]));
			radix2 #(.width(width)) rd_st0_987  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[987]), .rdlo_in(a0_wr[2011]),  .coef_in(coef[987]), .rdup_out(a1_wr[987]), .rdlo_out(a1_wr[2011]));
			radix2 #(.width(width)) rd_st0_988  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[988]), .rdlo_in(a0_wr[2012]),  .coef_in(coef[988]), .rdup_out(a1_wr[988]), .rdlo_out(a1_wr[2012]));
			radix2 #(.width(width)) rd_st0_989  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[989]), .rdlo_in(a0_wr[2013]),  .coef_in(coef[989]), .rdup_out(a1_wr[989]), .rdlo_out(a1_wr[2013]));
			radix2 #(.width(width)) rd_st0_990  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[990]), .rdlo_in(a0_wr[2014]),  .coef_in(coef[990]), .rdup_out(a1_wr[990]), .rdlo_out(a1_wr[2014]));
			radix2 #(.width(width)) rd_st0_991  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[991]), .rdlo_in(a0_wr[2015]),  .coef_in(coef[991]), .rdup_out(a1_wr[991]), .rdlo_out(a1_wr[2015]));
			radix2 #(.width(width)) rd_st0_992  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[992]), .rdlo_in(a0_wr[2016]),  .coef_in(coef[992]), .rdup_out(a1_wr[992]), .rdlo_out(a1_wr[2016]));
			radix2 #(.width(width)) rd_st0_993  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[993]), .rdlo_in(a0_wr[2017]),  .coef_in(coef[993]), .rdup_out(a1_wr[993]), .rdlo_out(a1_wr[2017]));
			radix2 #(.width(width)) rd_st0_994  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[994]), .rdlo_in(a0_wr[2018]),  .coef_in(coef[994]), .rdup_out(a1_wr[994]), .rdlo_out(a1_wr[2018]));
			radix2 #(.width(width)) rd_st0_995  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[995]), .rdlo_in(a0_wr[2019]),  .coef_in(coef[995]), .rdup_out(a1_wr[995]), .rdlo_out(a1_wr[2019]));
			radix2 #(.width(width)) rd_st0_996  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[996]), .rdlo_in(a0_wr[2020]),  .coef_in(coef[996]), .rdup_out(a1_wr[996]), .rdlo_out(a1_wr[2020]));
			radix2 #(.width(width)) rd_st0_997  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[997]), .rdlo_in(a0_wr[2021]),  .coef_in(coef[997]), .rdup_out(a1_wr[997]), .rdlo_out(a1_wr[2021]));
			radix2 #(.width(width)) rd_st0_998  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[998]), .rdlo_in(a0_wr[2022]),  .coef_in(coef[998]), .rdup_out(a1_wr[998]), .rdlo_out(a1_wr[2022]));
			radix2 #(.width(width)) rd_st0_999  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[999]), .rdlo_in(a0_wr[2023]),  .coef_in(coef[999]), .rdup_out(a1_wr[999]), .rdlo_out(a1_wr[2023]));
			radix2 #(.width(width)) rd_st0_1000  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[1000]), .rdlo_in(a0_wr[2024]),  .coef_in(coef[1000]), .rdup_out(a1_wr[1000]), .rdlo_out(a1_wr[2024]));
			radix2 #(.width(width)) rd_st0_1001  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[1001]), .rdlo_in(a0_wr[2025]),  .coef_in(coef[1001]), .rdup_out(a1_wr[1001]), .rdlo_out(a1_wr[2025]));
			radix2 #(.width(width)) rd_st0_1002  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[1002]), .rdlo_in(a0_wr[2026]),  .coef_in(coef[1002]), .rdup_out(a1_wr[1002]), .rdlo_out(a1_wr[2026]));
			radix2 #(.width(width)) rd_st0_1003  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[1003]), .rdlo_in(a0_wr[2027]),  .coef_in(coef[1003]), .rdup_out(a1_wr[1003]), .rdlo_out(a1_wr[2027]));
			radix2 #(.width(width)) rd_st0_1004  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[1004]), .rdlo_in(a0_wr[2028]),  .coef_in(coef[1004]), .rdup_out(a1_wr[1004]), .rdlo_out(a1_wr[2028]));
			radix2 #(.width(width)) rd_st0_1005  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[1005]), .rdlo_in(a0_wr[2029]),  .coef_in(coef[1005]), .rdup_out(a1_wr[1005]), .rdlo_out(a1_wr[2029]));
			radix2 #(.width(width)) rd_st0_1006  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[1006]), .rdlo_in(a0_wr[2030]),  .coef_in(coef[1006]), .rdup_out(a1_wr[1006]), .rdlo_out(a1_wr[2030]));
			radix2 #(.width(width)) rd_st0_1007  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[1007]), .rdlo_in(a0_wr[2031]),  .coef_in(coef[1007]), .rdup_out(a1_wr[1007]), .rdlo_out(a1_wr[2031]));
			radix2 #(.width(width)) rd_st0_1008  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[1008]), .rdlo_in(a0_wr[2032]),  .coef_in(coef[1008]), .rdup_out(a1_wr[1008]), .rdlo_out(a1_wr[2032]));
			radix2 #(.width(width)) rd_st0_1009  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[1009]), .rdlo_in(a0_wr[2033]),  .coef_in(coef[1009]), .rdup_out(a1_wr[1009]), .rdlo_out(a1_wr[2033]));
			radix2 #(.width(width)) rd_st0_1010  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[1010]), .rdlo_in(a0_wr[2034]),  .coef_in(coef[1010]), .rdup_out(a1_wr[1010]), .rdlo_out(a1_wr[2034]));
			radix2 #(.width(width)) rd_st0_1011  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[1011]), .rdlo_in(a0_wr[2035]),  .coef_in(coef[1011]), .rdup_out(a1_wr[1011]), .rdlo_out(a1_wr[2035]));
			radix2 #(.width(width)) rd_st0_1012  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[1012]), .rdlo_in(a0_wr[2036]),  .coef_in(coef[1012]), .rdup_out(a1_wr[1012]), .rdlo_out(a1_wr[2036]));
			radix2 #(.width(width)) rd_st0_1013  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[1013]), .rdlo_in(a0_wr[2037]),  .coef_in(coef[1013]), .rdup_out(a1_wr[1013]), .rdlo_out(a1_wr[2037]));
			radix2 #(.width(width)) rd_st0_1014  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[1014]), .rdlo_in(a0_wr[2038]),  .coef_in(coef[1014]), .rdup_out(a1_wr[1014]), .rdlo_out(a1_wr[2038]));
			radix2 #(.width(width)) rd_st0_1015  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[1015]), .rdlo_in(a0_wr[2039]),  .coef_in(coef[1015]), .rdup_out(a1_wr[1015]), .rdlo_out(a1_wr[2039]));
			radix2 #(.width(width)) rd_st0_1016  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[1016]), .rdlo_in(a0_wr[2040]),  .coef_in(coef[1016]), .rdup_out(a1_wr[1016]), .rdlo_out(a1_wr[2040]));
			radix2 #(.width(width)) rd_st0_1017  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[1017]), .rdlo_in(a0_wr[2041]),  .coef_in(coef[1017]), .rdup_out(a1_wr[1017]), .rdlo_out(a1_wr[2041]));
			radix2 #(.width(width)) rd_st0_1018  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[1018]), .rdlo_in(a0_wr[2042]),  .coef_in(coef[1018]), .rdup_out(a1_wr[1018]), .rdlo_out(a1_wr[2042]));
			radix2 #(.width(width)) rd_st0_1019  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[1019]), .rdlo_in(a0_wr[2043]),  .coef_in(coef[1019]), .rdup_out(a1_wr[1019]), .rdlo_out(a1_wr[2043]));
			radix2 #(.width(width)) rd_st0_1020  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[1020]), .rdlo_in(a0_wr[2044]),  .coef_in(coef[1020]), .rdup_out(a1_wr[1020]), .rdlo_out(a1_wr[2044]));
			radix2 #(.width(width)) rd_st0_1021  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[1021]), .rdlo_in(a0_wr[2045]),  .coef_in(coef[1021]), .rdup_out(a1_wr[1021]), .rdlo_out(a1_wr[2045]));
			radix2 #(.width(width)) rd_st0_1022  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[1022]), .rdlo_in(a0_wr[2046]),  .coef_in(coef[1022]), .rdup_out(a1_wr[1022]), .rdlo_out(a1_wr[2046]));
			radix2 #(.width(width)) rd_st0_1023  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a0_wr[1023]), .rdlo_in(a0_wr[2047]),  .coef_in(coef[1023]), .rdup_out(a1_wr[1023]), .rdlo_out(a1_wr[2047]));

		//--- radix stage 1
			radix2 #(.width(width)) rd_st1_0   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[0]), .rdlo_in(a1_wr[512]),  .coef_in(coef[0]), .rdup_out(a2_wr[0]), .rdlo_out(a2_wr[512]));
			radix2 #(.width(width)) rd_st1_1   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1]), .rdlo_in(a1_wr[513]),  .coef_in(coef[2]), .rdup_out(a2_wr[1]), .rdlo_out(a2_wr[513]));
			radix2 #(.width(width)) rd_st1_2   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[2]), .rdlo_in(a1_wr[514]),  .coef_in(coef[4]), .rdup_out(a2_wr[2]), .rdlo_out(a2_wr[514]));
			radix2 #(.width(width)) rd_st1_3   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[3]), .rdlo_in(a1_wr[515]),  .coef_in(coef[6]), .rdup_out(a2_wr[3]), .rdlo_out(a2_wr[515]));
			radix2 #(.width(width)) rd_st1_4   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[4]), .rdlo_in(a1_wr[516]),  .coef_in(coef[8]), .rdup_out(a2_wr[4]), .rdlo_out(a2_wr[516]));
			radix2 #(.width(width)) rd_st1_5   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[5]), .rdlo_in(a1_wr[517]),  .coef_in(coef[10]), .rdup_out(a2_wr[5]), .rdlo_out(a2_wr[517]));
			radix2 #(.width(width)) rd_st1_6   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[6]), .rdlo_in(a1_wr[518]),  .coef_in(coef[12]), .rdup_out(a2_wr[6]), .rdlo_out(a2_wr[518]));
			radix2 #(.width(width)) rd_st1_7   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[7]), .rdlo_in(a1_wr[519]),  .coef_in(coef[14]), .rdup_out(a2_wr[7]), .rdlo_out(a2_wr[519]));
			radix2 #(.width(width)) rd_st1_8   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[8]), .rdlo_in(a1_wr[520]),  .coef_in(coef[16]), .rdup_out(a2_wr[8]), .rdlo_out(a2_wr[520]));
			radix2 #(.width(width)) rd_st1_9   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[9]), .rdlo_in(a1_wr[521]),  .coef_in(coef[18]), .rdup_out(a2_wr[9]), .rdlo_out(a2_wr[521]));
			radix2 #(.width(width)) rd_st1_10  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[10]), .rdlo_in(a1_wr[522]),  .coef_in(coef[20]), .rdup_out(a2_wr[10]), .rdlo_out(a2_wr[522]));
			radix2 #(.width(width)) rd_st1_11  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[11]), .rdlo_in(a1_wr[523]),  .coef_in(coef[22]), .rdup_out(a2_wr[11]), .rdlo_out(a2_wr[523]));
			radix2 #(.width(width)) rd_st1_12  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[12]), .rdlo_in(a1_wr[524]),  .coef_in(coef[24]), .rdup_out(a2_wr[12]), .rdlo_out(a2_wr[524]));
			radix2 #(.width(width)) rd_st1_13  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[13]), .rdlo_in(a1_wr[525]),  .coef_in(coef[26]), .rdup_out(a2_wr[13]), .rdlo_out(a2_wr[525]));
			radix2 #(.width(width)) rd_st1_14  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[14]), .rdlo_in(a1_wr[526]),  .coef_in(coef[28]), .rdup_out(a2_wr[14]), .rdlo_out(a2_wr[526]));
			radix2 #(.width(width)) rd_st1_15  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[15]), .rdlo_in(a1_wr[527]),  .coef_in(coef[30]), .rdup_out(a2_wr[15]), .rdlo_out(a2_wr[527]));
			radix2 #(.width(width)) rd_st1_16  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[16]), .rdlo_in(a1_wr[528]),  .coef_in(coef[32]), .rdup_out(a2_wr[16]), .rdlo_out(a2_wr[528]));
			radix2 #(.width(width)) rd_st1_17  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[17]), .rdlo_in(a1_wr[529]),  .coef_in(coef[34]), .rdup_out(a2_wr[17]), .rdlo_out(a2_wr[529]));
			radix2 #(.width(width)) rd_st1_18  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[18]), .rdlo_in(a1_wr[530]),  .coef_in(coef[36]), .rdup_out(a2_wr[18]), .rdlo_out(a2_wr[530]));
			radix2 #(.width(width)) rd_st1_19  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[19]), .rdlo_in(a1_wr[531]),  .coef_in(coef[38]), .rdup_out(a2_wr[19]), .rdlo_out(a2_wr[531]));
			radix2 #(.width(width)) rd_st1_20  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[20]), .rdlo_in(a1_wr[532]),  .coef_in(coef[40]), .rdup_out(a2_wr[20]), .rdlo_out(a2_wr[532]));
			radix2 #(.width(width)) rd_st1_21  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[21]), .rdlo_in(a1_wr[533]),  .coef_in(coef[42]), .rdup_out(a2_wr[21]), .rdlo_out(a2_wr[533]));
			radix2 #(.width(width)) rd_st1_22  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[22]), .rdlo_in(a1_wr[534]),  .coef_in(coef[44]), .rdup_out(a2_wr[22]), .rdlo_out(a2_wr[534]));
			radix2 #(.width(width)) rd_st1_23  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[23]), .rdlo_in(a1_wr[535]),  .coef_in(coef[46]), .rdup_out(a2_wr[23]), .rdlo_out(a2_wr[535]));
			radix2 #(.width(width)) rd_st1_24  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[24]), .rdlo_in(a1_wr[536]),  .coef_in(coef[48]), .rdup_out(a2_wr[24]), .rdlo_out(a2_wr[536]));
			radix2 #(.width(width)) rd_st1_25  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[25]), .rdlo_in(a1_wr[537]),  .coef_in(coef[50]), .rdup_out(a2_wr[25]), .rdlo_out(a2_wr[537]));
			radix2 #(.width(width)) rd_st1_26  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[26]), .rdlo_in(a1_wr[538]),  .coef_in(coef[52]), .rdup_out(a2_wr[26]), .rdlo_out(a2_wr[538]));
			radix2 #(.width(width)) rd_st1_27  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[27]), .rdlo_in(a1_wr[539]),  .coef_in(coef[54]), .rdup_out(a2_wr[27]), .rdlo_out(a2_wr[539]));
			radix2 #(.width(width)) rd_st1_28  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[28]), .rdlo_in(a1_wr[540]),  .coef_in(coef[56]), .rdup_out(a2_wr[28]), .rdlo_out(a2_wr[540]));
			radix2 #(.width(width)) rd_st1_29  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[29]), .rdlo_in(a1_wr[541]),  .coef_in(coef[58]), .rdup_out(a2_wr[29]), .rdlo_out(a2_wr[541]));
			radix2 #(.width(width)) rd_st1_30  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[30]), .rdlo_in(a1_wr[542]),  .coef_in(coef[60]), .rdup_out(a2_wr[30]), .rdlo_out(a2_wr[542]));
			radix2 #(.width(width)) rd_st1_31  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[31]), .rdlo_in(a1_wr[543]),  .coef_in(coef[62]), .rdup_out(a2_wr[31]), .rdlo_out(a2_wr[543]));
			radix2 #(.width(width)) rd_st1_32  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[32]), .rdlo_in(a1_wr[544]),  .coef_in(coef[64]), .rdup_out(a2_wr[32]), .rdlo_out(a2_wr[544]));
			radix2 #(.width(width)) rd_st1_33  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[33]), .rdlo_in(a1_wr[545]),  .coef_in(coef[66]), .rdup_out(a2_wr[33]), .rdlo_out(a2_wr[545]));
			radix2 #(.width(width)) rd_st1_34  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[34]), .rdlo_in(a1_wr[546]),  .coef_in(coef[68]), .rdup_out(a2_wr[34]), .rdlo_out(a2_wr[546]));
			radix2 #(.width(width)) rd_st1_35  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[35]), .rdlo_in(a1_wr[547]),  .coef_in(coef[70]), .rdup_out(a2_wr[35]), .rdlo_out(a2_wr[547]));
			radix2 #(.width(width)) rd_st1_36  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[36]), .rdlo_in(a1_wr[548]),  .coef_in(coef[72]), .rdup_out(a2_wr[36]), .rdlo_out(a2_wr[548]));
			radix2 #(.width(width)) rd_st1_37  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[37]), .rdlo_in(a1_wr[549]),  .coef_in(coef[74]), .rdup_out(a2_wr[37]), .rdlo_out(a2_wr[549]));
			radix2 #(.width(width)) rd_st1_38  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[38]), .rdlo_in(a1_wr[550]),  .coef_in(coef[76]), .rdup_out(a2_wr[38]), .rdlo_out(a2_wr[550]));
			radix2 #(.width(width)) rd_st1_39  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[39]), .rdlo_in(a1_wr[551]),  .coef_in(coef[78]), .rdup_out(a2_wr[39]), .rdlo_out(a2_wr[551]));
			radix2 #(.width(width)) rd_st1_40  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[40]), .rdlo_in(a1_wr[552]),  .coef_in(coef[80]), .rdup_out(a2_wr[40]), .rdlo_out(a2_wr[552]));
			radix2 #(.width(width)) rd_st1_41  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[41]), .rdlo_in(a1_wr[553]),  .coef_in(coef[82]), .rdup_out(a2_wr[41]), .rdlo_out(a2_wr[553]));
			radix2 #(.width(width)) rd_st1_42  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[42]), .rdlo_in(a1_wr[554]),  .coef_in(coef[84]), .rdup_out(a2_wr[42]), .rdlo_out(a2_wr[554]));
			radix2 #(.width(width)) rd_st1_43  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[43]), .rdlo_in(a1_wr[555]),  .coef_in(coef[86]), .rdup_out(a2_wr[43]), .rdlo_out(a2_wr[555]));
			radix2 #(.width(width)) rd_st1_44  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[44]), .rdlo_in(a1_wr[556]),  .coef_in(coef[88]), .rdup_out(a2_wr[44]), .rdlo_out(a2_wr[556]));
			radix2 #(.width(width)) rd_st1_45  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[45]), .rdlo_in(a1_wr[557]),  .coef_in(coef[90]), .rdup_out(a2_wr[45]), .rdlo_out(a2_wr[557]));
			radix2 #(.width(width)) rd_st1_46  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[46]), .rdlo_in(a1_wr[558]),  .coef_in(coef[92]), .rdup_out(a2_wr[46]), .rdlo_out(a2_wr[558]));
			radix2 #(.width(width)) rd_st1_47  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[47]), .rdlo_in(a1_wr[559]),  .coef_in(coef[94]), .rdup_out(a2_wr[47]), .rdlo_out(a2_wr[559]));
			radix2 #(.width(width)) rd_st1_48  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[48]), .rdlo_in(a1_wr[560]),  .coef_in(coef[96]), .rdup_out(a2_wr[48]), .rdlo_out(a2_wr[560]));
			radix2 #(.width(width)) rd_st1_49  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[49]), .rdlo_in(a1_wr[561]),  .coef_in(coef[98]), .rdup_out(a2_wr[49]), .rdlo_out(a2_wr[561]));
			radix2 #(.width(width)) rd_st1_50  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[50]), .rdlo_in(a1_wr[562]),  .coef_in(coef[100]), .rdup_out(a2_wr[50]), .rdlo_out(a2_wr[562]));
			radix2 #(.width(width)) rd_st1_51  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[51]), .rdlo_in(a1_wr[563]),  .coef_in(coef[102]), .rdup_out(a2_wr[51]), .rdlo_out(a2_wr[563]));
			radix2 #(.width(width)) rd_st1_52  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[52]), .rdlo_in(a1_wr[564]),  .coef_in(coef[104]), .rdup_out(a2_wr[52]), .rdlo_out(a2_wr[564]));
			radix2 #(.width(width)) rd_st1_53  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[53]), .rdlo_in(a1_wr[565]),  .coef_in(coef[106]), .rdup_out(a2_wr[53]), .rdlo_out(a2_wr[565]));
			radix2 #(.width(width)) rd_st1_54  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[54]), .rdlo_in(a1_wr[566]),  .coef_in(coef[108]), .rdup_out(a2_wr[54]), .rdlo_out(a2_wr[566]));
			radix2 #(.width(width)) rd_st1_55  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[55]), .rdlo_in(a1_wr[567]),  .coef_in(coef[110]), .rdup_out(a2_wr[55]), .rdlo_out(a2_wr[567]));
			radix2 #(.width(width)) rd_st1_56  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[56]), .rdlo_in(a1_wr[568]),  .coef_in(coef[112]), .rdup_out(a2_wr[56]), .rdlo_out(a2_wr[568]));
			radix2 #(.width(width)) rd_st1_57  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[57]), .rdlo_in(a1_wr[569]),  .coef_in(coef[114]), .rdup_out(a2_wr[57]), .rdlo_out(a2_wr[569]));
			radix2 #(.width(width)) rd_st1_58  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[58]), .rdlo_in(a1_wr[570]),  .coef_in(coef[116]), .rdup_out(a2_wr[58]), .rdlo_out(a2_wr[570]));
			radix2 #(.width(width)) rd_st1_59  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[59]), .rdlo_in(a1_wr[571]),  .coef_in(coef[118]), .rdup_out(a2_wr[59]), .rdlo_out(a2_wr[571]));
			radix2 #(.width(width)) rd_st1_60  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[60]), .rdlo_in(a1_wr[572]),  .coef_in(coef[120]), .rdup_out(a2_wr[60]), .rdlo_out(a2_wr[572]));
			radix2 #(.width(width)) rd_st1_61  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[61]), .rdlo_in(a1_wr[573]),  .coef_in(coef[122]), .rdup_out(a2_wr[61]), .rdlo_out(a2_wr[573]));
			radix2 #(.width(width)) rd_st1_62  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[62]), .rdlo_in(a1_wr[574]),  .coef_in(coef[124]), .rdup_out(a2_wr[62]), .rdlo_out(a2_wr[574]));
			radix2 #(.width(width)) rd_st1_63  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[63]), .rdlo_in(a1_wr[575]),  .coef_in(coef[126]), .rdup_out(a2_wr[63]), .rdlo_out(a2_wr[575]));
			radix2 #(.width(width)) rd_st1_64  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[64]), .rdlo_in(a1_wr[576]),  .coef_in(coef[128]), .rdup_out(a2_wr[64]), .rdlo_out(a2_wr[576]));
			radix2 #(.width(width)) rd_st1_65  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[65]), .rdlo_in(a1_wr[577]),  .coef_in(coef[130]), .rdup_out(a2_wr[65]), .rdlo_out(a2_wr[577]));
			radix2 #(.width(width)) rd_st1_66  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[66]), .rdlo_in(a1_wr[578]),  .coef_in(coef[132]), .rdup_out(a2_wr[66]), .rdlo_out(a2_wr[578]));
			radix2 #(.width(width)) rd_st1_67  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[67]), .rdlo_in(a1_wr[579]),  .coef_in(coef[134]), .rdup_out(a2_wr[67]), .rdlo_out(a2_wr[579]));
			radix2 #(.width(width)) rd_st1_68  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[68]), .rdlo_in(a1_wr[580]),  .coef_in(coef[136]), .rdup_out(a2_wr[68]), .rdlo_out(a2_wr[580]));
			radix2 #(.width(width)) rd_st1_69  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[69]), .rdlo_in(a1_wr[581]),  .coef_in(coef[138]), .rdup_out(a2_wr[69]), .rdlo_out(a2_wr[581]));
			radix2 #(.width(width)) rd_st1_70  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[70]), .rdlo_in(a1_wr[582]),  .coef_in(coef[140]), .rdup_out(a2_wr[70]), .rdlo_out(a2_wr[582]));
			radix2 #(.width(width)) rd_st1_71  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[71]), .rdlo_in(a1_wr[583]),  .coef_in(coef[142]), .rdup_out(a2_wr[71]), .rdlo_out(a2_wr[583]));
			radix2 #(.width(width)) rd_st1_72  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[72]), .rdlo_in(a1_wr[584]),  .coef_in(coef[144]), .rdup_out(a2_wr[72]), .rdlo_out(a2_wr[584]));
			radix2 #(.width(width)) rd_st1_73  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[73]), .rdlo_in(a1_wr[585]),  .coef_in(coef[146]), .rdup_out(a2_wr[73]), .rdlo_out(a2_wr[585]));
			radix2 #(.width(width)) rd_st1_74  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[74]), .rdlo_in(a1_wr[586]),  .coef_in(coef[148]), .rdup_out(a2_wr[74]), .rdlo_out(a2_wr[586]));
			radix2 #(.width(width)) rd_st1_75  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[75]), .rdlo_in(a1_wr[587]),  .coef_in(coef[150]), .rdup_out(a2_wr[75]), .rdlo_out(a2_wr[587]));
			radix2 #(.width(width)) rd_st1_76  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[76]), .rdlo_in(a1_wr[588]),  .coef_in(coef[152]), .rdup_out(a2_wr[76]), .rdlo_out(a2_wr[588]));
			radix2 #(.width(width)) rd_st1_77  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[77]), .rdlo_in(a1_wr[589]),  .coef_in(coef[154]), .rdup_out(a2_wr[77]), .rdlo_out(a2_wr[589]));
			radix2 #(.width(width)) rd_st1_78  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[78]), .rdlo_in(a1_wr[590]),  .coef_in(coef[156]), .rdup_out(a2_wr[78]), .rdlo_out(a2_wr[590]));
			radix2 #(.width(width)) rd_st1_79  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[79]), .rdlo_in(a1_wr[591]),  .coef_in(coef[158]), .rdup_out(a2_wr[79]), .rdlo_out(a2_wr[591]));
			radix2 #(.width(width)) rd_st1_80  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[80]), .rdlo_in(a1_wr[592]),  .coef_in(coef[160]), .rdup_out(a2_wr[80]), .rdlo_out(a2_wr[592]));
			radix2 #(.width(width)) rd_st1_81  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[81]), .rdlo_in(a1_wr[593]),  .coef_in(coef[162]), .rdup_out(a2_wr[81]), .rdlo_out(a2_wr[593]));
			radix2 #(.width(width)) rd_st1_82  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[82]), .rdlo_in(a1_wr[594]),  .coef_in(coef[164]), .rdup_out(a2_wr[82]), .rdlo_out(a2_wr[594]));
			radix2 #(.width(width)) rd_st1_83  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[83]), .rdlo_in(a1_wr[595]),  .coef_in(coef[166]), .rdup_out(a2_wr[83]), .rdlo_out(a2_wr[595]));
			radix2 #(.width(width)) rd_st1_84  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[84]), .rdlo_in(a1_wr[596]),  .coef_in(coef[168]), .rdup_out(a2_wr[84]), .rdlo_out(a2_wr[596]));
			radix2 #(.width(width)) rd_st1_85  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[85]), .rdlo_in(a1_wr[597]),  .coef_in(coef[170]), .rdup_out(a2_wr[85]), .rdlo_out(a2_wr[597]));
			radix2 #(.width(width)) rd_st1_86  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[86]), .rdlo_in(a1_wr[598]),  .coef_in(coef[172]), .rdup_out(a2_wr[86]), .rdlo_out(a2_wr[598]));
			radix2 #(.width(width)) rd_st1_87  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[87]), .rdlo_in(a1_wr[599]),  .coef_in(coef[174]), .rdup_out(a2_wr[87]), .rdlo_out(a2_wr[599]));
			radix2 #(.width(width)) rd_st1_88  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[88]), .rdlo_in(a1_wr[600]),  .coef_in(coef[176]), .rdup_out(a2_wr[88]), .rdlo_out(a2_wr[600]));
			radix2 #(.width(width)) rd_st1_89  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[89]), .rdlo_in(a1_wr[601]),  .coef_in(coef[178]), .rdup_out(a2_wr[89]), .rdlo_out(a2_wr[601]));
			radix2 #(.width(width)) rd_st1_90  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[90]), .rdlo_in(a1_wr[602]),  .coef_in(coef[180]), .rdup_out(a2_wr[90]), .rdlo_out(a2_wr[602]));
			radix2 #(.width(width)) rd_st1_91  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[91]), .rdlo_in(a1_wr[603]),  .coef_in(coef[182]), .rdup_out(a2_wr[91]), .rdlo_out(a2_wr[603]));
			radix2 #(.width(width)) rd_st1_92  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[92]), .rdlo_in(a1_wr[604]),  .coef_in(coef[184]), .rdup_out(a2_wr[92]), .rdlo_out(a2_wr[604]));
			radix2 #(.width(width)) rd_st1_93  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[93]), .rdlo_in(a1_wr[605]),  .coef_in(coef[186]), .rdup_out(a2_wr[93]), .rdlo_out(a2_wr[605]));
			radix2 #(.width(width)) rd_st1_94  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[94]), .rdlo_in(a1_wr[606]),  .coef_in(coef[188]), .rdup_out(a2_wr[94]), .rdlo_out(a2_wr[606]));
			radix2 #(.width(width)) rd_st1_95  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[95]), .rdlo_in(a1_wr[607]),  .coef_in(coef[190]), .rdup_out(a2_wr[95]), .rdlo_out(a2_wr[607]));
			radix2 #(.width(width)) rd_st1_96  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[96]), .rdlo_in(a1_wr[608]),  .coef_in(coef[192]), .rdup_out(a2_wr[96]), .rdlo_out(a2_wr[608]));
			radix2 #(.width(width)) rd_st1_97  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[97]), .rdlo_in(a1_wr[609]),  .coef_in(coef[194]), .rdup_out(a2_wr[97]), .rdlo_out(a2_wr[609]));
			radix2 #(.width(width)) rd_st1_98  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[98]), .rdlo_in(a1_wr[610]),  .coef_in(coef[196]), .rdup_out(a2_wr[98]), .rdlo_out(a2_wr[610]));
			radix2 #(.width(width)) rd_st1_99  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[99]), .rdlo_in(a1_wr[611]),  .coef_in(coef[198]), .rdup_out(a2_wr[99]), .rdlo_out(a2_wr[611]));
			radix2 #(.width(width)) rd_st1_100  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[100]), .rdlo_in(a1_wr[612]),  .coef_in(coef[200]), .rdup_out(a2_wr[100]), .rdlo_out(a2_wr[612]));
			radix2 #(.width(width)) rd_st1_101  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[101]), .rdlo_in(a1_wr[613]),  .coef_in(coef[202]), .rdup_out(a2_wr[101]), .rdlo_out(a2_wr[613]));
			radix2 #(.width(width)) rd_st1_102  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[102]), .rdlo_in(a1_wr[614]),  .coef_in(coef[204]), .rdup_out(a2_wr[102]), .rdlo_out(a2_wr[614]));
			radix2 #(.width(width)) rd_st1_103  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[103]), .rdlo_in(a1_wr[615]),  .coef_in(coef[206]), .rdup_out(a2_wr[103]), .rdlo_out(a2_wr[615]));
			radix2 #(.width(width)) rd_st1_104  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[104]), .rdlo_in(a1_wr[616]),  .coef_in(coef[208]), .rdup_out(a2_wr[104]), .rdlo_out(a2_wr[616]));
			radix2 #(.width(width)) rd_st1_105  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[105]), .rdlo_in(a1_wr[617]),  .coef_in(coef[210]), .rdup_out(a2_wr[105]), .rdlo_out(a2_wr[617]));
			radix2 #(.width(width)) rd_st1_106  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[106]), .rdlo_in(a1_wr[618]),  .coef_in(coef[212]), .rdup_out(a2_wr[106]), .rdlo_out(a2_wr[618]));
			radix2 #(.width(width)) rd_st1_107  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[107]), .rdlo_in(a1_wr[619]),  .coef_in(coef[214]), .rdup_out(a2_wr[107]), .rdlo_out(a2_wr[619]));
			radix2 #(.width(width)) rd_st1_108  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[108]), .rdlo_in(a1_wr[620]),  .coef_in(coef[216]), .rdup_out(a2_wr[108]), .rdlo_out(a2_wr[620]));
			radix2 #(.width(width)) rd_st1_109  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[109]), .rdlo_in(a1_wr[621]),  .coef_in(coef[218]), .rdup_out(a2_wr[109]), .rdlo_out(a2_wr[621]));
			radix2 #(.width(width)) rd_st1_110  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[110]), .rdlo_in(a1_wr[622]),  .coef_in(coef[220]), .rdup_out(a2_wr[110]), .rdlo_out(a2_wr[622]));
			radix2 #(.width(width)) rd_st1_111  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[111]), .rdlo_in(a1_wr[623]),  .coef_in(coef[222]), .rdup_out(a2_wr[111]), .rdlo_out(a2_wr[623]));
			radix2 #(.width(width)) rd_st1_112  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[112]), .rdlo_in(a1_wr[624]),  .coef_in(coef[224]), .rdup_out(a2_wr[112]), .rdlo_out(a2_wr[624]));
			radix2 #(.width(width)) rd_st1_113  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[113]), .rdlo_in(a1_wr[625]),  .coef_in(coef[226]), .rdup_out(a2_wr[113]), .rdlo_out(a2_wr[625]));
			radix2 #(.width(width)) rd_st1_114  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[114]), .rdlo_in(a1_wr[626]),  .coef_in(coef[228]), .rdup_out(a2_wr[114]), .rdlo_out(a2_wr[626]));
			radix2 #(.width(width)) rd_st1_115  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[115]), .rdlo_in(a1_wr[627]),  .coef_in(coef[230]), .rdup_out(a2_wr[115]), .rdlo_out(a2_wr[627]));
			radix2 #(.width(width)) rd_st1_116  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[116]), .rdlo_in(a1_wr[628]),  .coef_in(coef[232]), .rdup_out(a2_wr[116]), .rdlo_out(a2_wr[628]));
			radix2 #(.width(width)) rd_st1_117  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[117]), .rdlo_in(a1_wr[629]),  .coef_in(coef[234]), .rdup_out(a2_wr[117]), .rdlo_out(a2_wr[629]));
			radix2 #(.width(width)) rd_st1_118  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[118]), .rdlo_in(a1_wr[630]),  .coef_in(coef[236]), .rdup_out(a2_wr[118]), .rdlo_out(a2_wr[630]));
			radix2 #(.width(width)) rd_st1_119  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[119]), .rdlo_in(a1_wr[631]),  .coef_in(coef[238]), .rdup_out(a2_wr[119]), .rdlo_out(a2_wr[631]));
			radix2 #(.width(width)) rd_st1_120  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[120]), .rdlo_in(a1_wr[632]),  .coef_in(coef[240]), .rdup_out(a2_wr[120]), .rdlo_out(a2_wr[632]));
			radix2 #(.width(width)) rd_st1_121  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[121]), .rdlo_in(a1_wr[633]),  .coef_in(coef[242]), .rdup_out(a2_wr[121]), .rdlo_out(a2_wr[633]));
			radix2 #(.width(width)) rd_st1_122  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[122]), .rdlo_in(a1_wr[634]),  .coef_in(coef[244]), .rdup_out(a2_wr[122]), .rdlo_out(a2_wr[634]));
			radix2 #(.width(width)) rd_st1_123  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[123]), .rdlo_in(a1_wr[635]),  .coef_in(coef[246]), .rdup_out(a2_wr[123]), .rdlo_out(a2_wr[635]));
			radix2 #(.width(width)) rd_st1_124  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[124]), .rdlo_in(a1_wr[636]),  .coef_in(coef[248]), .rdup_out(a2_wr[124]), .rdlo_out(a2_wr[636]));
			radix2 #(.width(width)) rd_st1_125  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[125]), .rdlo_in(a1_wr[637]),  .coef_in(coef[250]), .rdup_out(a2_wr[125]), .rdlo_out(a2_wr[637]));
			radix2 #(.width(width)) rd_st1_126  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[126]), .rdlo_in(a1_wr[638]),  .coef_in(coef[252]), .rdup_out(a2_wr[126]), .rdlo_out(a2_wr[638]));
			radix2 #(.width(width)) rd_st1_127  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[127]), .rdlo_in(a1_wr[639]),  .coef_in(coef[254]), .rdup_out(a2_wr[127]), .rdlo_out(a2_wr[639]));
			radix2 #(.width(width)) rd_st1_128  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[128]), .rdlo_in(a1_wr[640]),  .coef_in(coef[256]), .rdup_out(a2_wr[128]), .rdlo_out(a2_wr[640]));
			radix2 #(.width(width)) rd_st1_129  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[129]), .rdlo_in(a1_wr[641]),  .coef_in(coef[258]), .rdup_out(a2_wr[129]), .rdlo_out(a2_wr[641]));
			radix2 #(.width(width)) rd_st1_130  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[130]), .rdlo_in(a1_wr[642]),  .coef_in(coef[260]), .rdup_out(a2_wr[130]), .rdlo_out(a2_wr[642]));
			radix2 #(.width(width)) rd_st1_131  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[131]), .rdlo_in(a1_wr[643]),  .coef_in(coef[262]), .rdup_out(a2_wr[131]), .rdlo_out(a2_wr[643]));
			radix2 #(.width(width)) rd_st1_132  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[132]), .rdlo_in(a1_wr[644]),  .coef_in(coef[264]), .rdup_out(a2_wr[132]), .rdlo_out(a2_wr[644]));
			radix2 #(.width(width)) rd_st1_133  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[133]), .rdlo_in(a1_wr[645]),  .coef_in(coef[266]), .rdup_out(a2_wr[133]), .rdlo_out(a2_wr[645]));
			radix2 #(.width(width)) rd_st1_134  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[134]), .rdlo_in(a1_wr[646]),  .coef_in(coef[268]), .rdup_out(a2_wr[134]), .rdlo_out(a2_wr[646]));
			radix2 #(.width(width)) rd_st1_135  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[135]), .rdlo_in(a1_wr[647]),  .coef_in(coef[270]), .rdup_out(a2_wr[135]), .rdlo_out(a2_wr[647]));
			radix2 #(.width(width)) rd_st1_136  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[136]), .rdlo_in(a1_wr[648]),  .coef_in(coef[272]), .rdup_out(a2_wr[136]), .rdlo_out(a2_wr[648]));
			radix2 #(.width(width)) rd_st1_137  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[137]), .rdlo_in(a1_wr[649]),  .coef_in(coef[274]), .rdup_out(a2_wr[137]), .rdlo_out(a2_wr[649]));
			radix2 #(.width(width)) rd_st1_138  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[138]), .rdlo_in(a1_wr[650]),  .coef_in(coef[276]), .rdup_out(a2_wr[138]), .rdlo_out(a2_wr[650]));
			radix2 #(.width(width)) rd_st1_139  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[139]), .rdlo_in(a1_wr[651]),  .coef_in(coef[278]), .rdup_out(a2_wr[139]), .rdlo_out(a2_wr[651]));
			radix2 #(.width(width)) rd_st1_140  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[140]), .rdlo_in(a1_wr[652]),  .coef_in(coef[280]), .rdup_out(a2_wr[140]), .rdlo_out(a2_wr[652]));
			radix2 #(.width(width)) rd_st1_141  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[141]), .rdlo_in(a1_wr[653]),  .coef_in(coef[282]), .rdup_out(a2_wr[141]), .rdlo_out(a2_wr[653]));
			radix2 #(.width(width)) rd_st1_142  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[142]), .rdlo_in(a1_wr[654]),  .coef_in(coef[284]), .rdup_out(a2_wr[142]), .rdlo_out(a2_wr[654]));
			radix2 #(.width(width)) rd_st1_143  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[143]), .rdlo_in(a1_wr[655]),  .coef_in(coef[286]), .rdup_out(a2_wr[143]), .rdlo_out(a2_wr[655]));
			radix2 #(.width(width)) rd_st1_144  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[144]), .rdlo_in(a1_wr[656]),  .coef_in(coef[288]), .rdup_out(a2_wr[144]), .rdlo_out(a2_wr[656]));
			radix2 #(.width(width)) rd_st1_145  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[145]), .rdlo_in(a1_wr[657]),  .coef_in(coef[290]), .rdup_out(a2_wr[145]), .rdlo_out(a2_wr[657]));
			radix2 #(.width(width)) rd_st1_146  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[146]), .rdlo_in(a1_wr[658]),  .coef_in(coef[292]), .rdup_out(a2_wr[146]), .rdlo_out(a2_wr[658]));
			radix2 #(.width(width)) rd_st1_147  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[147]), .rdlo_in(a1_wr[659]),  .coef_in(coef[294]), .rdup_out(a2_wr[147]), .rdlo_out(a2_wr[659]));
			radix2 #(.width(width)) rd_st1_148  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[148]), .rdlo_in(a1_wr[660]),  .coef_in(coef[296]), .rdup_out(a2_wr[148]), .rdlo_out(a2_wr[660]));
			radix2 #(.width(width)) rd_st1_149  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[149]), .rdlo_in(a1_wr[661]),  .coef_in(coef[298]), .rdup_out(a2_wr[149]), .rdlo_out(a2_wr[661]));
			radix2 #(.width(width)) rd_st1_150  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[150]), .rdlo_in(a1_wr[662]),  .coef_in(coef[300]), .rdup_out(a2_wr[150]), .rdlo_out(a2_wr[662]));
			radix2 #(.width(width)) rd_st1_151  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[151]), .rdlo_in(a1_wr[663]),  .coef_in(coef[302]), .rdup_out(a2_wr[151]), .rdlo_out(a2_wr[663]));
			radix2 #(.width(width)) rd_st1_152  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[152]), .rdlo_in(a1_wr[664]),  .coef_in(coef[304]), .rdup_out(a2_wr[152]), .rdlo_out(a2_wr[664]));
			radix2 #(.width(width)) rd_st1_153  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[153]), .rdlo_in(a1_wr[665]),  .coef_in(coef[306]), .rdup_out(a2_wr[153]), .rdlo_out(a2_wr[665]));
			radix2 #(.width(width)) rd_st1_154  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[154]), .rdlo_in(a1_wr[666]),  .coef_in(coef[308]), .rdup_out(a2_wr[154]), .rdlo_out(a2_wr[666]));
			radix2 #(.width(width)) rd_st1_155  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[155]), .rdlo_in(a1_wr[667]),  .coef_in(coef[310]), .rdup_out(a2_wr[155]), .rdlo_out(a2_wr[667]));
			radix2 #(.width(width)) rd_st1_156  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[156]), .rdlo_in(a1_wr[668]),  .coef_in(coef[312]), .rdup_out(a2_wr[156]), .rdlo_out(a2_wr[668]));
			radix2 #(.width(width)) rd_st1_157  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[157]), .rdlo_in(a1_wr[669]),  .coef_in(coef[314]), .rdup_out(a2_wr[157]), .rdlo_out(a2_wr[669]));
			radix2 #(.width(width)) rd_st1_158  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[158]), .rdlo_in(a1_wr[670]),  .coef_in(coef[316]), .rdup_out(a2_wr[158]), .rdlo_out(a2_wr[670]));
			radix2 #(.width(width)) rd_st1_159  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[159]), .rdlo_in(a1_wr[671]),  .coef_in(coef[318]), .rdup_out(a2_wr[159]), .rdlo_out(a2_wr[671]));
			radix2 #(.width(width)) rd_st1_160  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[160]), .rdlo_in(a1_wr[672]),  .coef_in(coef[320]), .rdup_out(a2_wr[160]), .rdlo_out(a2_wr[672]));
			radix2 #(.width(width)) rd_st1_161  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[161]), .rdlo_in(a1_wr[673]),  .coef_in(coef[322]), .rdup_out(a2_wr[161]), .rdlo_out(a2_wr[673]));
			radix2 #(.width(width)) rd_st1_162  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[162]), .rdlo_in(a1_wr[674]),  .coef_in(coef[324]), .rdup_out(a2_wr[162]), .rdlo_out(a2_wr[674]));
			radix2 #(.width(width)) rd_st1_163  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[163]), .rdlo_in(a1_wr[675]),  .coef_in(coef[326]), .rdup_out(a2_wr[163]), .rdlo_out(a2_wr[675]));
			radix2 #(.width(width)) rd_st1_164  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[164]), .rdlo_in(a1_wr[676]),  .coef_in(coef[328]), .rdup_out(a2_wr[164]), .rdlo_out(a2_wr[676]));
			radix2 #(.width(width)) rd_st1_165  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[165]), .rdlo_in(a1_wr[677]),  .coef_in(coef[330]), .rdup_out(a2_wr[165]), .rdlo_out(a2_wr[677]));
			radix2 #(.width(width)) rd_st1_166  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[166]), .rdlo_in(a1_wr[678]),  .coef_in(coef[332]), .rdup_out(a2_wr[166]), .rdlo_out(a2_wr[678]));
			radix2 #(.width(width)) rd_st1_167  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[167]), .rdlo_in(a1_wr[679]),  .coef_in(coef[334]), .rdup_out(a2_wr[167]), .rdlo_out(a2_wr[679]));
			radix2 #(.width(width)) rd_st1_168  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[168]), .rdlo_in(a1_wr[680]),  .coef_in(coef[336]), .rdup_out(a2_wr[168]), .rdlo_out(a2_wr[680]));
			radix2 #(.width(width)) rd_st1_169  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[169]), .rdlo_in(a1_wr[681]),  .coef_in(coef[338]), .rdup_out(a2_wr[169]), .rdlo_out(a2_wr[681]));
			radix2 #(.width(width)) rd_st1_170  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[170]), .rdlo_in(a1_wr[682]),  .coef_in(coef[340]), .rdup_out(a2_wr[170]), .rdlo_out(a2_wr[682]));
			radix2 #(.width(width)) rd_st1_171  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[171]), .rdlo_in(a1_wr[683]),  .coef_in(coef[342]), .rdup_out(a2_wr[171]), .rdlo_out(a2_wr[683]));
			radix2 #(.width(width)) rd_st1_172  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[172]), .rdlo_in(a1_wr[684]),  .coef_in(coef[344]), .rdup_out(a2_wr[172]), .rdlo_out(a2_wr[684]));
			radix2 #(.width(width)) rd_st1_173  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[173]), .rdlo_in(a1_wr[685]),  .coef_in(coef[346]), .rdup_out(a2_wr[173]), .rdlo_out(a2_wr[685]));
			radix2 #(.width(width)) rd_st1_174  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[174]), .rdlo_in(a1_wr[686]),  .coef_in(coef[348]), .rdup_out(a2_wr[174]), .rdlo_out(a2_wr[686]));
			radix2 #(.width(width)) rd_st1_175  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[175]), .rdlo_in(a1_wr[687]),  .coef_in(coef[350]), .rdup_out(a2_wr[175]), .rdlo_out(a2_wr[687]));
			radix2 #(.width(width)) rd_st1_176  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[176]), .rdlo_in(a1_wr[688]),  .coef_in(coef[352]), .rdup_out(a2_wr[176]), .rdlo_out(a2_wr[688]));
			radix2 #(.width(width)) rd_st1_177  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[177]), .rdlo_in(a1_wr[689]),  .coef_in(coef[354]), .rdup_out(a2_wr[177]), .rdlo_out(a2_wr[689]));
			radix2 #(.width(width)) rd_st1_178  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[178]), .rdlo_in(a1_wr[690]),  .coef_in(coef[356]), .rdup_out(a2_wr[178]), .rdlo_out(a2_wr[690]));
			radix2 #(.width(width)) rd_st1_179  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[179]), .rdlo_in(a1_wr[691]),  .coef_in(coef[358]), .rdup_out(a2_wr[179]), .rdlo_out(a2_wr[691]));
			radix2 #(.width(width)) rd_st1_180  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[180]), .rdlo_in(a1_wr[692]),  .coef_in(coef[360]), .rdup_out(a2_wr[180]), .rdlo_out(a2_wr[692]));
			radix2 #(.width(width)) rd_st1_181  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[181]), .rdlo_in(a1_wr[693]),  .coef_in(coef[362]), .rdup_out(a2_wr[181]), .rdlo_out(a2_wr[693]));
			radix2 #(.width(width)) rd_st1_182  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[182]), .rdlo_in(a1_wr[694]),  .coef_in(coef[364]), .rdup_out(a2_wr[182]), .rdlo_out(a2_wr[694]));
			radix2 #(.width(width)) rd_st1_183  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[183]), .rdlo_in(a1_wr[695]),  .coef_in(coef[366]), .rdup_out(a2_wr[183]), .rdlo_out(a2_wr[695]));
			radix2 #(.width(width)) rd_st1_184  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[184]), .rdlo_in(a1_wr[696]),  .coef_in(coef[368]), .rdup_out(a2_wr[184]), .rdlo_out(a2_wr[696]));
			radix2 #(.width(width)) rd_st1_185  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[185]), .rdlo_in(a1_wr[697]),  .coef_in(coef[370]), .rdup_out(a2_wr[185]), .rdlo_out(a2_wr[697]));
			radix2 #(.width(width)) rd_st1_186  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[186]), .rdlo_in(a1_wr[698]),  .coef_in(coef[372]), .rdup_out(a2_wr[186]), .rdlo_out(a2_wr[698]));
			radix2 #(.width(width)) rd_st1_187  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[187]), .rdlo_in(a1_wr[699]),  .coef_in(coef[374]), .rdup_out(a2_wr[187]), .rdlo_out(a2_wr[699]));
			radix2 #(.width(width)) rd_st1_188  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[188]), .rdlo_in(a1_wr[700]),  .coef_in(coef[376]), .rdup_out(a2_wr[188]), .rdlo_out(a2_wr[700]));
			radix2 #(.width(width)) rd_st1_189  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[189]), .rdlo_in(a1_wr[701]),  .coef_in(coef[378]), .rdup_out(a2_wr[189]), .rdlo_out(a2_wr[701]));
			radix2 #(.width(width)) rd_st1_190  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[190]), .rdlo_in(a1_wr[702]),  .coef_in(coef[380]), .rdup_out(a2_wr[190]), .rdlo_out(a2_wr[702]));
			radix2 #(.width(width)) rd_st1_191  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[191]), .rdlo_in(a1_wr[703]),  .coef_in(coef[382]), .rdup_out(a2_wr[191]), .rdlo_out(a2_wr[703]));
			radix2 #(.width(width)) rd_st1_192  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[192]), .rdlo_in(a1_wr[704]),  .coef_in(coef[384]), .rdup_out(a2_wr[192]), .rdlo_out(a2_wr[704]));
			radix2 #(.width(width)) rd_st1_193  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[193]), .rdlo_in(a1_wr[705]),  .coef_in(coef[386]), .rdup_out(a2_wr[193]), .rdlo_out(a2_wr[705]));
			radix2 #(.width(width)) rd_st1_194  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[194]), .rdlo_in(a1_wr[706]),  .coef_in(coef[388]), .rdup_out(a2_wr[194]), .rdlo_out(a2_wr[706]));
			radix2 #(.width(width)) rd_st1_195  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[195]), .rdlo_in(a1_wr[707]),  .coef_in(coef[390]), .rdup_out(a2_wr[195]), .rdlo_out(a2_wr[707]));
			radix2 #(.width(width)) rd_st1_196  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[196]), .rdlo_in(a1_wr[708]),  .coef_in(coef[392]), .rdup_out(a2_wr[196]), .rdlo_out(a2_wr[708]));
			radix2 #(.width(width)) rd_st1_197  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[197]), .rdlo_in(a1_wr[709]),  .coef_in(coef[394]), .rdup_out(a2_wr[197]), .rdlo_out(a2_wr[709]));
			radix2 #(.width(width)) rd_st1_198  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[198]), .rdlo_in(a1_wr[710]),  .coef_in(coef[396]), .rdup_out(a2_wr[198]), .rdlo_out(a2_wr[710]));
			radix2 #(.width(width)) rd_st1_199  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[199]), .rdlo_in(a1_wr[711]),  .coef_in(coef[398]), .rdup_out(a2_wr[199]), .rdlo_out(a2_wr[711]));
			radix2 #(.width(width)) rd_st1_200  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[200]), .rdlo_in(a1_wr[712]),  .coef_in(coef[400]), .rdup_out(a2_wr[200]), .rdlo_out(a2_wr[712]));
			radix2 #(.width(width)) rd_st1_201  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[201]), .rdlo_in(a1_wr[713]),  .coef_in(coef[402]), .rdup_out(a2_wr[201]), .rdlo_out(a2_wr[713]));
			radix2 #(.width(width)) rd_st1_202  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[202]), .rdlo_in(a1_wr[714]),  .coef_in(coef[404]), .rdup_out(a2_wr[202]), .rdlo_out(a2_wr[714]));
			radix2 #(.width(width)) rd_st1_203  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[203]), .rdlo_in(a1_wr[715]),  .coef_in(coef[406]), .rdup_out(a2_wr[203]), .rdlo_out(a2_wr[715]));
			radix2 #(.width(width)) rd_st1_204  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[204]), .rdlo_in(a1_wr[716]),  .coef_in(coef[408]), .rdup_out(a2_wr[204]), .rdlo_out(a2_wr[716]));
			radix2 #(.width(width)) rd_st1_205  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[205]), .rdlo_in(a1_wr[717]),  .coef_in(coef[410]), .rdup_out(a2_wr[205]), .rdlo_out(a2_wr[717]));
			radix2 #(.width(width)) rd_st1_206  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[206]), .rdlo_in(a1_wr[718]),  .coef_in(coef[412]), .rdup_out(a2_wr[206]), .rdlo_out(a2_wr[718]));
			radix2 #(.width(width)) rd_st1_207  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[207]), .rdlo_in(a1_wr[719]),  .coef_in(coef[414]), .rdup_out(a2_wr[207]), .rdlo_out(a2_wr[719]));
			radix2 #(.width(width)) rd_st1_208  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[208]), .rdlo_in(a1_wr[720]),  .coef_in(coef[416]), .rdup_out(a2_wr[208]), .rdlo_out(a2_wr[720]));
			radix2 #(.width(width)) rd_st1_209  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[209]), .rdlo_in(a1_wr[721]),  .coef_in(coef[418]), .rdup_out(a2_wr[209]), .rdlo_out(a2_wr[721]));
			radix2 #(.width(width)) rd_st1_210  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[210]), .rdlo_in(a1_wr[722]),  .coef_in(coef[420]), .rdup_out(a2_wr[210]), .rdlo_out(a2_wr[722]));
			radix2 #(.width(width)) rd_st1_211  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[211]), .rdlo_in(a1_wr[723]),  .coef_in(coef[422]), .rdup_out(a2_wr[211]), .rdlo_out(a2_wr[723]));
			radix2 #(.width(width)) rd_st1_212  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[212]), .rdlo_in(a1_wr[724]),  .coef_in(coef[424]), .rdup_out(a2_wr[212]), .rdlo_out(a2_wr[724]));
			radix2 #(.width(width)) rd_st1_213  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[213]), .rdlo_in(a1_wr[725]),  .coef_in(coef[426]), .rdup_out(a2_wr[213]), .rdlo_out(a2_wr[725]));
			radix2 #(.width(width)) rd_st1_214  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[214]), .rdlo_in(a1_wr[726]),  .coef_in(coef[428]), .rdup_out(a2_wr[214]), .rdlo_out(a2_wr[726]));
			radix2 #(.width(width)) rd_st1_215  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[215]), .rdlo_in(a1_wr[727]),  .coef_in(coef[430]), .rdup_out(a2_wr[215]), .rdlo_out(a2_wr[727]));
			radix2 #(.width(width)) rd_st1_216  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[216]), .rdlo_in(a1_wr[728]),  .coef_in(coef[432]), .rdup_out(a2_wr[216]), .rdlo_out(a2_wr[728]));
			radix2 #(.width(width)) rd_st1_217  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[217]), .rdlo_in(a1_wr[729]),  .coef_in(coef[434]), .rdup_out(a2_wr[217]), .rdlo_out(a2_wr[729]));
			radix2 #(.width(width)) rd_st1_218  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[218]), .rdlo_in(a1_wr[730]),  .coef_in(coef[436]), .rdup_out(a2_wr[218]), .rdlo_out(a2_wr[730]));
			radix2 #(.width(width)) rd_st1_219  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[219]), .rdlo_in(a1_wr[731]),  .coef_in(coef[438]), .rdup_out(a2_wr[219]), .rdlo_out(a2_wr[731]));
			radix2 #(.width(width)) rd_st1_220  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[220]), .rdlo_in(a1_wr[732]),  .coef_in(coef[440]), .rdup_out(a2_wr[220]), .rdlo_out(a2_wr[732]));
			radix2 #(.width(width)) rd_st1_221  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[221]), .rdlo_in(a1_wr[733]),  .coef_in(coef[442]), .rdup_out(a2_wr[221]), .rdlo_out(a2_wr[733]));
			radix2 #(.width(width)) rd_st1_222  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[222]), .rdlo_in(a1_wr[734]),  .coef_in(coef[444]), .rdup_out(a2_wr[222]), .rdlo_out(a2_wr[734]));
			radix2 #(.width(width)) rd_st1_223  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[223]), .rdlo_in(a1_wr[735]),  .coef_in(coef[446]), .rdup_out(a2_wr[223]), .rdlo_out(a2_wr[735]));
			radix2 #(.width(width)) rd_st1_224  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[224]), .rdlo_in(a1_wr[736]),  .coef_in(coef[448]), .rdup_out(a2_wr[224]), .rdlo_out(a2_wr[736]));
			radix2 #(.width(width)) rd_st1_225  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[225]), .rdlo_in(a1_wr[737]),  .coef_in(coef[450]), .rdup_out(a2_wr[225]), .rdlo_out(a2_wr[737]));
			radix2 #(.width(width)) rd_st1_226  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[226]), .rdlo_in(a1_wr[738]),  .coef_in(coef[452]), .rdup_out(a2_wr[226]), .rdlo_out(a2_wr[738]));
			radix2 #(.width(width)) rd_st1_227  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[227]), .rdlo_in(a1_wr[739]),  .coef_in(coef[454]), .rdup_out(a2_wr[227]), .rdlo_out(a2_wr[739]));
			radix2 #(.width(width)) rd_st1_228  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[228]), .rdlo_in(a1_wr[740]),  .coef_in(coef[456]), .rdup_out(a2_wr[228]), .rdlo_out(a2_wr[740]));
			radix2 #(.width(width)) rd_st1_229  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[229]), .rdlo_in(a1_wr[741]),  .coef_in(coef[458]), .rdup_out(a2_wr[229]), .rdlo_out(a2_wr[741]));
			radix2 #(.width(width)) rd_st1_230  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[230]), .rdlo_in(a1_wr[742]),  .coef_in(coef[460]), .rdup_out(a2_wr[230]), .rdlo_out(a2_wr[742]));
			radix2 #(.width(width)) rd_st1_231  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[231]), .rdlo_in(a1_wr[743]),  .coef_in(coef[462]), .rdup_out(a2_wr[231]), .rdlo_out(a2_wr[743]));
			radix2 #(.width(width)) rd_st1_232  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[232]), .rdlo_in(a1_wr[744]),  .coef_in(coef[464]), .rdup_out(a2_wr[232]), .rdlo_out(a2_wr[744]));
			radix2 #(.width(width)) rd_st1_233  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[233]), .rdlo_in(a1_wr[745]),  .coef_in(coef[466]), .rdup_out(a2_wr[233]), .rdlo_out(a2_wr[745]));
			radix2 #(.width(width)) rd_st1_234  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[234]), .rdlo_in(a1_wr[746]),  .coef_in(coef[468]), .rdup_out(a2_wr[234]), .rdlo_out(a2_wr[746]));
			radix2 #(.width(width)) rd_st1_235  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[235]), .rdlo_in(a1_wr[747]),  .coef_in(coef[470]), .rdup_out(a2_wr[235]), .rdlo_out(a2_wr[747]));
			radix2 #(.width(width)) rd_st1_236  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[236]), .rdlo_in(a1_wr[748]),  .coef_in(coef[472]), .rdup_out(a2_wr[236]), .rdlo_out(a2_wr[748]));
			radix2 #(.width(width)) rd_st1_237  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[237]), .rdlo_in(a1_wr[749]),  .coef_in(coef[474]), .rdup_out(a2_wr[237]), .rdlo_out(a2_wr[749]));
			radix2 #(.width(width)) rd_st1_238  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[238]), .rdlo_in(a1_wr[750]),  .coef_in(coef[476]), .rdup_out(a2_wr[238]), .rdlo_out(a2_wr[750]));
			radix2 #(.width(width)) rd_st1_239  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[239]), .rdlo_in(a1_wr[751]),  .coef_in(coef[478]), .rdup_out(a2_wr[239]), .rdlo_out(a2_wr[751]));
			radix2 #(.width(width)) rd_st1_240  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[240]), .rdlo_in(a1_wr[752]),  .coef_in(coef[480]), .rdup_out(a2_wr[240]), .rdlo_out(a2_wr[752]));
			radix2 #(.width(width)) rd_st1_241  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[241]), .rdlo_in(a1_wr[753]),  .coef_in(coef[482]), .rdup_out(a2_wr[241]), .rdlo_out(a2_wr[753]));
			radix2 #(.width(width)) rd_st1_242  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[242]), .rdlo_in(a1_wr[754]),  .coef_in(coef[484]), .rdup_out(a2_wr[242]), .rdlo_out(a2_wr[754]));
			radix2 #(.width(width)) rd_st1_243  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[243]), .rdlo_in(a1_wr[755]),  .coef_in(coef[486]), .rdup_out(a2_wr[243]), .rdlo_out(a2_wr[755]));
			radix2 #(.width(width)) rd_st1_244  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[244]), .rdlo_in(a1_wr[756]),  .coef_in(coef[488]), .rdup_out(a2_wr[244]), .rdlo_out(a2_wr[756]));
			radix2 #(.width(width)) rd_st1_245  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[245]), .rdlo_in(a1_wr[757]),  .coef_in(coef[490]), .rdup_out(a2_wr[245]), .rdlo_out(a2_wr[757]));
			radix2 #(.width(width)) rd_st1_246  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[246]), .rdlo_in(a1_wr[758]),  .coef_in(coef[492]), .rdup_out(a2_wr[246]), .rdlo_out(a2_wr[758]));
			radix2 #(.width(width)) rd_st1_247  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[247]), .rdlo_in(a1_wr[759]),  .coef_in(coef[494]), .rdup_out(a2_wr[247]), .rdlo_out(a2_wr[759]));
			radix2 #(.width(width)) rd_st1_248  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[248]), .rdlo_in(a1_wr[760]),  .coef_in(coef[496]), .rdup_out(a2_wr[248]), .rdlo_out(a2_wr[760]));
			radix2 #(.width(width)) rd_st1_249  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[249]), .rdlo_in(a1_wr[761]),  .coef_in(coef[498]), .rdup_out(a2_wr[249]), .rdlo_out(a2_wr[761]));
			radix2 #(.width(width)) rd_st1_250  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[250]), .rdlo_in(a1_wr[762]),  .coef_in(coef[500]), .rdup_out(a2_wr[250]), .rdlo_out(a2_wr[762]));
			radix2 #(.width(width)) rd_st1_251  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[251]), .rdlo_in(a1_wr[763]),  .coef_in(coef[502]), .rdup_out(a2_wr[251]), .rdlo_out(a2_wr[763]));
			radix2 #(.width(width)) rd_st1_252  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[252]), .rdlo_in(a1_wr[764]),  .coef_in(coef[504]), .rdup_out(a2_wr[252]), .rdlo_out(a2_wr[764]));
			radix2 #(.width(width)) rd_st1_253  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[253]), .rdlo_in(a1_wr[765]),  .coef_in(coef[506]), .rdup_out(a2_wr[253]), .rdlo_out(a2_wr[765]));
			radix2 #(.width(width)) rd_st1_254  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[254]), .rdlo_in(a1_wr[766]),  .coef_in(coef[508]), .rdup_out(a2_wr[254]), .rdlo_out(a2_wr[766]));
			radix2 #(.width(width)) rd_st1_255  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[255]), .rdlo_in(a1_wr[767]),  .coef_in(coef[510]), .rdup_out(a2_wr[255]), .rdlo_out(a2_wr[767]));
			radix2 #(.width(width)) rd_st1_256  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[256]), .rdlo_in(a1_wr[768]),  .coef_in(coef[512]), .rdup_out(a2_wr[256]), .rdlo_out(a2_wr[768]));
			radix2 #(.width(width)) rd_st1_257  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[257]), .rdlo_in(a1_wr[769]),  .coef_in(coef[514]), .rdup_out(a2_wr[257]), .rdlo_out(a2_wr[769]));
			radix2 #(.width(width)) rd_st1_258  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[258]), .rdlo_in(a1_wr[770]),  .coef_in(coef[516]), .rdup_out(a2_wr[258]), .rdlo_out(a2_wr[770]));
			radix2 #(.width(width)) rd_st1_259  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[259]), .rdlo_in(a1_wr[771]),  .coef_in(coef[518]), .rdup_out(a2_wr[259]), .rdlo_out(a2_wr[771]));
			radix2 #(.width(width)) rd_st1_260  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[260]), .rdlo_in(a1_wr[772]),  .coef_in(coef[520]), .rdup_out(a2_wr[260]), .rdlo_out(a2_wr[772]));
			radix2 #(.width(width)) rd_st1_261  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[261]), .rdlo_in(a1_wr[773]),  .coef_in(coef[522]), .rdup_out(a2_wr[261]), .rdlo_out(a2_wr[773]));
			radix2 #(.width(width)) rd_st1_262  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[262]), .rdlo_in(a1_wr[774]),  .coef_in(coef[524]), .rdup_out(a2_wr[262]), .rdlo_out(a2_wr[774]));
			radix2 #(.width(width)) rd_st1_263  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[263]), .rdlo_in(a1_wr[775]),  .coef_in(coef[526]), .rdup_out(a2_wr[263]), .rdlo_out(a2_wr[775]));
			radix2 #(.width(width)) rd_st1_264  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[264]), .rdlo_in(a1_wr[776]),  .coef_in(coef[528]), .rdup_out(a2_wr[264]), .rdlo_out(a2_wr[776]));
			radix2 #(.width(width)) rd_st1_265  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[265]), .rdlo_in(a1_wr[777]),  .coef_in(coef[530]), .rdup_out(a2_wr[265]), .rdlo_out(a2_wr[777]));
			radix2 #(.width(width)) rd_st1_266  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[266]), .rdlo_in(a1_wr[778]),  .coef_in(coef[532]), .rdup_out(a2_wr[266]), .rdlo_out(a2_wr[778]));
			radix2 #(.width(width)) rd_st1_267  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[267]), .rdlo_in(a1_wr[779]),  .coef_in(coef[534]), .rdup_out(a2_wr[267]), .rdlo_out(a2_wr[779]));
			radix2 #(.width(width)) rd_st1_268  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[268]), .rdlo_in(a1_wr[780]),  .coef_in(coef[536]), .rdup_out(a2_wr[268]), .rdlo_out(a2_wr[780]));
			radix2 #(.width(width)) rd_st1_269  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[269]), .rdlo_in(a1_wr[781]),  .coef_in(coef[538]), .rdup_out(a2_wr[269]), .rdlo_out(a2_wr[781]));
			radix2 #(.width(width)) rd_st1_270  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[270]), .rdlo_in(a1_wr[782]),  .coef_in(coef[540]), .rdup_out(a2_wr[270]), .rdlo_out(a2_wr[782]));
			radix2 #(.width(width)) rd_st1_271  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[271]), .rdlo_in(a1_wr[783]),  .coef_in(coef[542]), .rdup_out(a2_wr[271]), .rdlo_out(a2_wr[783]));
			radix2 #(.width(width)) rd_st1_272  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[272]), .rdlo_in(a1_wr[784]),  .coef_in(coef[544]), .rdup_out(a2_wr[272]), .rdlo_out(a2_wr[784]));
			radix2 #(.width(width)) rd_st1_273  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[273]), .rdlo_in(a1_wr[785]),  .coef_in(coef[546]), .rdup_out(a2_wr[273]), .rdlo_out(a2_wr[785]));
			radix2 #(.width(width)) rd_st1_274  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[274]), .rdlo_in(a1_wr[786]),  .coef_in(coef[548]), .rdup_out(a2_wr[274]), .rdlo_out(a2_wr[786]));
			radix2 #(.width(width)) rd_st1_275  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[275]), .rdlo_in(a1_wr[787]),  .coef_in(coef[550]), .rdup_out(a2_wr[275]), .rdlo_out(a2_wr[787]));
			radix2 #(.width(width)) rd_st1_276  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[276]), .rdlo_in(a1_wr[788]),  .coef_in(coef[552]), .rdup_out(a2_wr[276]), .rdlo_out(a2_wr[788]));
			radix2 #(.width(width)) rd_st1_277  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[277]), .rdlo_in(a1_wr[789]),  .coef_in(coef[554]), .rdup_out(a2_wr[277]), .rdlo_out(a2_wr[789]));
			radix2 #(.width(width)) rd_st1_278  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[278]), .rdlo_in(a1_wr[790]),  .coef_in(coef[556]), .rdup_out(a2_wr[278]), .rdlo_out(a2_wr[790]));
			radix2 #(.width(width)) rd_st1_279  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[279]), .rdlo_in(a1_wr[791]),  .coef_in(coef[558]), .rdup_out(a2_wr[279]), .rdlo_out(a2_wr[791]));
			radix2 #(.width(width)) rd_st1_280  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[280]), .rdlo_in(a1_wr[792]),  .coef_in(coef[560]), .rdup_out(a2_wr[280]), .rdlo_out(a2_wr[792]));
			radix2 #(.width(width)) rd_st1_281  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[281]), .rdlo_in(a1_wr[793]),  .coef_in(coef[562]), .rdup_out(a2_wr[281]), .rdlo_out(a2_wr[793]));
			radix2 #(.width(width)) rd_st1_282  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[282]), .rdlo_in(a1_wr[794]),  .coef_in(coef[564]), .rdup_out(a2_wr[282]), .rdlo_out(a2_wr[794]));
			radix2 #(.width(width)) rd_st1_283  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[283]), .rdlo_in(a1_wr[795]),  .coef_in(coef[566]), .rdup_out(a2_wr[283]), .rdlo_out(a2_wr[795]));
			radix2 #(.width(width)) rd_st1_284  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[284]), .rdlo_in(a1_wr[796]),  .coef_in(coef[568]), .rdup_out(a2_wr[284]), .rdlo_out(a2_wr[796]));
			radix2 #(.width(width)) rd_st1_285  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[285]), .rdlo_in(a1_wr[797]),  .coef_in(coef[570]), .rdup_out(a2_wr[285]), .rdlo_out(a2_wr[797]));
			radix2 #(.width(width)) rd_st1_286  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[286]), .rdlo_in(a1_wr[798]),  .coef_in(coef[572]), .rdup_out(a2_wr[286]), .rdlo_out(a2_wr[798]));
			radix2 #(.width(width)) rd_st1_287  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[287]), .rdlo_in(a1_wr[799]),  .coef_in(coef[574]), .rdup_out(a2_wr[287]), .rdlo_out(a2_wr[799]));
			radix2 #(.width(width)) rd_st1_288  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[288]), .rdlo_in(a1_wr[800]),  .coef_in(coef[576]), .rdup_out(a2_wr[288]), .rdlo_out(a2_wr[800]));
			radix2 #(.width(width)) rd_st1_289  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[289]), .rdlo_in(a1_wr[801]),  .coef_in(coef[578]), .rdup_out(a2_wr[289]), .rdlo_out(a2_wr[801]));
			radix2 #(.width(width)) rd_st1_290  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[290]), .rdlo_in(a1_wr[802]),  .coef_in(coef[580]), .rdup_out(a2_wr[290]), .rdlo_out(a2_wr[802]));
			radix2 #(.width(width)) rd_st1_291  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[291]), .rdlo_in(a1_wr[803]),  .coef_in(coef[582]), .rdup_out(a2_wr[291]), .rdlo_out(a2_wr[803]));
			radix2 #(.width(width)) rd_st1_292  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[292]), .rdlo_in(a1_wr[804]),  .coef_in(coef[584]), .rdup_out(a2_wr[292]), .rdlo_out(a2_wr[804]));
			radix2 #(.width(width)) rd_st1_293  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[293]), .rdlo_in(a1_wr[805]),  .coef_in(coef[586]), .rdup_out(a2_wr[293]), .rdlo_out(a2_wr[805]));
			radix2 #(.width(width)) rd_st1_294  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[294]), .rdlo_in(a1_wr[806]),  .coef_in(coef[588]), .rdup_out(a2_wr[294]), .rdlo_out(a2_wr[806]));
			radix2 #(.width(width)) rd_st1_295  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[295]), .rdlo_in(a1_wr[807]),  .coef_in(coef[590]), .rdup_out(a2_wr[295]), .rdlo_out(a2_wr[807]));
			radix2 #(.width(width)) rd_st1_296  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[296]), .rdlo_in(a1_wr[808]),  .coef_in(coef[592]), .rdup_out(a2_wr[296]), .rdlo_out(a2_wr[808]));
			radix2 #(.width(width)) rd_st1_297  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[297]), .rdlo_in(a1_wr[809]),  .coef_in(coef[594]), .rdup_out(a2_wr[297]), .rdlo_out(a2_wr[809]));
			radix2 #(.width(width)) rd_st1_298  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[298]), .rdlo_in(a1_wr[810]),  .coef_in(coef[596]), .rdup_out(a2_wr[298]), .rdlo_out(a2_wr[810]));
			radix2 #(.width(width)) rd_st1_299  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[299]), .rdlo_in(a1_wr[811]),  .coef_in(coef[598]), .rdup_out(a2_wr[299]), .rdlo_out(a2_wr[811]));
			radix2 #(.width(width)) rd_st1_300  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[300]), .rdlo_in(a1_wr[812]),  .coef_in(coef[600]), .rdup_out(a2_wr[300]), .rdlo_out(a2_wr[812]));
			radix2 #(.width(width)) rd_st1_301  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[301]), .rdlo_in(a1_wr[813]),  .coef_in(coef[602]), .rdup_out(a2_wr[301]), .rdlo_out(a2_wr[813]));
			radix2 #(.width(width)) rd_st1_302  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[302]), .rdlo_in(a1_wr[814]),  .coef_in(coef[604]), .rdup_out(a2_wr[302]), .rdlo_out(a2_wr[814]));
			radix2 #(.width(width)) rd_st1_303  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[303]), .rdlo_in(a1_wr[815]),  .coef_in(coef[606]), .rdup_out(a2_wr[303]), .rdlo_out(a2_wr[815]));
			radix2 #(.width(width)) rd_st1_304  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[304]), .rdlo_in(a1_wr[816]),  .coef_in(coef[608]), .rdup_out(a2_wr[304]), .rdlo_out(a2_wr[816]));
			radix2 #(.width(width)) rd_st1_305  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[305]), .rdlo_in(a1_wr[817]),  .coef_in(coef[610]), .rdup_out(a2_wr[305]), .rdlo_out(a2_wr[817]));
			radix2 #(.width(width)) rd_st1_306  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[306]), .rdlo_in(a1_wr[818]),  .coef_in(coef[612]), .rdup_out(a2_wr[306]), .rdlo_out(a2_wr[818]));
			radix2 #(.width(width)) rd_st1_307  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[307]), .rdlo_in(a1_wr[819]),  .coef_in(coef[614]), .rdup_out(a2_wr[307]), .rdlo_out(a2_wr[819]));
			radix2 #(.width(width)) rd_st1_308  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[308]), .rdlo_in(a1_wr[820]),  .coef_in(coef[616]), .rdup_out(a2_wr[308]), .rdlo_out(a2_wr[820]));
			radix2 #(.width(width)) rd_st1_309  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[309]), .rdlo_in(a1_wr[821]),  .coef_in(coef[618]), .rdup_out(a2_wr[309]), .rdlo_out(a2_wr[821]));
			radix2 #(.width(width)) rd_st1_310  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[310]), .rdlo_in(a1_wr[822]),  .coef_in(coef[620]), .rdup_out(a2_wr[310]), .rdlo_out(a2_wr[822]));
			radix2 #(.width(width)) rd_st1_311  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[311]), .rdlo_in(a1_wr[823]),  .coef_in(coef[622]), .rdup_out(a2_wr[311]), .rdlo_out(a2_wr[823]));
			radix2 #(.width(width)) rd_st1_312  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[312]), .rdlo_in(a1_wr[824]),  .coef_in(coef[624]), .rdup_out(a2_wr[312]), .rdlo_out(a2_wr[824]));
			radix2 #(.width(width)) rd_st1_313  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[313]), .rdlo_in(a1_wr[825]),  .coef_in(coef[626]), .rdup_out(a2_wr[313]), .rdlo_out(a2_wr[825]));
			radix2 #(.width(width)) rd_st1_314  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[314]), .rdlo_in(a1_wr[826]),  .coef_in(coef[628]), .rdup_out(a2_wr[314]), .rdlo_out(a2_wr[826]));
			radix2 #(.width(width)) rd_st1_315  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[315]), .rdlo_in(a1_wr[827]),  .coef_in(coef[630]), .rdup_out(a2_wr[315]), .rdlo_out(a2_wr[827]));
			radix2 #(.width(width)) rd_st1_316  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[316]), .rdlo_in(a1_wr[828]),  .coef_in(coef[632]), .rdup_out(a2_wr[316]), .rdlo_out(a2_wr[828]));
			radix2 #(.width(width)) rd_st1_317  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[317]), .rdlo_in(a1_wr[829]),  .coef_in(coef[634]), .rdup_out(a2_wr[317]), .rdlo_out(a2_wr[829]));
			radix2 #(.width(width)) rd_st1_318  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[318]), .rdlo_in(a1_wr[830]),  .coef_in(coef[636]), .rdup_out(a2_wr[318]), .rdlo_out(a2_wr[830]));
			radix2 #(.width(width)) rd_st1_319  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[319]), .rdlo_in(a1_wr[831]),  .coef_in(coef[638]), .rdup_out(a2_wr[319]), .rdlo_out(a2_wr[831]));
			radix2 #(.width(width)) rd_st1_320  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[320]), .rdlo_in(a1_wr[832]),  .coef_in(coef[640]), .rdup_out(a2_wr[320]), .rdlo_out(a2_wr[832]));
			radix2 #(.width(width)) rd_st1_321  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[321]), .rdlo_in(a1_wr[833]),  .coef_in(coef[642]), .rdup_out(a2_wr[321]), .rdlo_out(a2_wr[833]));
			radix2 #(.width(width)) rd_st1_322  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[322]), .rdlo_in(a1_wr[834]),  .coef_in(coef[644]), .rdup_out(a2_wr[322]), .rdlo_out(a2_wr[834]));
			radix2 #(.width(width)) rd_st1_323  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[323]), .rdlo_in(a1_wr[835]),  .coef_in(coef[646]), .rdup_out(a2_wr[323]), .rdlo_out(a2_wr[835]));
			radix2 #(.width(width)) rd_st1_324  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[324]), .rdlo_in(a1_wr[836]),  .coef_in(coef[648]), .rdup_out(a2_wr[324]), .rdlo_out(a2_wr[836]));
			radix2 #(.width(width)) rd_st1_325  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[325]), .rdlo_in(a1_wr[837]),  .coef_in(coef[650]), .rdup_out(a2_wr[325]), .rdlo_out(a2_wr[837]));
			radix2 #(.width(width)) rd_st1_326  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[326]), .rdlo_in(a1_wr[838]),  .coef_in(coef[652]), .rdup_out(a2_wr[326]), .rdlo_out(a2_wr[838]));
			radix2 #(.width(width)) rd_st1_327  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[327]), .rdlo_in(a1_wr[839]),  .coef_in(coef[654]), .rdup_out(a2_wr[327]), .rdlo_out(a2_wr[839]));
			radix2 #(.width(width)) rd_st1_328  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[328]), .rdlo_in(a1_wr[840]),  .coef_in(coef[656]), .rdup_out(a2_wr[328]), .rdlo_out(a2_wr[840]));
			radix2 #(.width(width)) rd_st1_329  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[329]), .rdlo_in(a1_wr[841]),  .coef_in(coef[658]), .rdup_out(a2_wr[329]), .rdlo_out(a2_wr[841]));
			radix2 #(.width(width)) rd_st1_330  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[330]), .rdlo_in(a1_wr[842]),  .coef_in(coef[660]), .rdup_out(a2_wr[330]), .rdlo_out(a2_wr[842]));
			radix2 #(.width(width)) rd_st1_331  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[331]), .rdlo_in(a1_wr[843]),  .coef_in(coef[662]), .rdup_out(a2_wr[331]), .rdlo_out(a2_wr[843]));
			radix2 #(.width(width)) rd_st1_332  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[332]), .rdlo_in(a1_wr[844]),  .coef_in(coef[664]), .rdup_out(a2_wr[332]), .rdlo_out(a2_wr[844]));
			radix2 #(.width(width)) rd_st1_333  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[333]), .rdlo_in(a1_wr[845]),  .coef_in(coef[666]), .rdup_out(a2_wr[333]), .rdlo_out(a2_wr[845]));
			radix2 #(.width(width)) rd_st1_334  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[334]), .rdlo_in(a1_wr[846]),  .coef_in(coef[668]), .rdup_out(a2_wr[334]), .rdlo_out(a2_wr[846]));
			radix2 #(.width(width)) rd_st1_335  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[335]), .rdlo_in(a1_wr[847]),  .coef_in(coef[670]), .rdup_out(a2_wr[335]), .rdlo_out(a2_wr[847]));
			radix2 #(.width(width)) rd_st1_336  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[336]), .rdlo_in(a1_wr[848]),  .coef_in(coef[672]), .rdup_out(a2_wr[336]), .rdlo_out(a2_wr[848]));
			radix2 #(.width(width)) rd_st1_337  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[337]), .rdlo_in(a1_wr[849]),  .coef_in(coef[674]), .rdup_out(a2_wr[337]), .rdlo_out(a2_wr[849]));
			radix2 #(.width(width)) rd_st1_338  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[338]), .rdlo_in(a1_wr[850]),  .coef_in(coef[676]), .rdup_out(a2_wr[338]), .rdlo_out(a2_wr[850]));
			radix2 #(.width(width)) rd_st1_339  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[339]), .rdlo_in(a1_wr[851]),  .coef_in(coef[678]), .rdup_out(a2_wr[339]), .rdlo_out(a2_wr[851]));
			radix2 #(.width(width)) rd_st1_340  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[340]), .rdlo_in(a1_wr[852]),  .coef_in(coef[680]), .rdup_out(a2_wr[340]), .rdlo_out(a2_wr[852]));
			radix2 #(.width(width)) rd_st1_341  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[341]), .rdlo_in(a1_wr[853]),  .coef_in(coef[682]), .rdup_out(a2_wr[341]), .rdlo_out(a2_wr[853]));
			radix2 #(.width(width)) rd_st1_342  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[342]), .rdlo_in(a1_wr[854]),  .coef_in(coef[684]), .rdup_out(a2_wr[342]), .rdlo_out(a2_wr[854]));
			radix2 #(.width(width)) rd_st1_343  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[343]), .rdlo_in(a1_wr[855]),  .coef_in(coef[686]), .rdup_out(a2_wr[343]), .rdlo_out(a2_wr[855]));
			radix2 #(.width(width)) rd_st1_344  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[344]), .rdlo_in(a1_wr[856]),  .coef_in(coef[688]), .rdup_out(a2_wr[344]), .rdlo_out(a2_wr[856]));
			radix2 #(.width(width)) rd_st1_345  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[345]), .rdlo_in(a1_wr[857]),  .coef_in(coef[690]), .rdup_out(a2_wr[345]), .rdlo_out(a2_wr[857]));
			radix2 #(.width(width)) rd_st1_346  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[346]), .rdlo_in(a1_wr[858]),  .coef_in(coef[692]), .rdup_out(a2_wr[346]), .rdlo_out(a2_wr[858]));
			radix2 #(.width(width)) rd_st1_347  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[347]), .rdlo_in(a1_wr[859]),  .coef_in(coef[694]), .rdup_out(a2_wr[347]), .rdlo_out(a2_wr[859]));
			radix2 #(.width(width)) rd_st1_348  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[348]), .rdlo_in(a1_wr[860]),  .coef_in(coef[696]), .rdup_out(a2_wr[348]), .rdlo_out(a2_wr[860]));
			radix2 #(.width(width)) rd_st1_349  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[349]), .rdlo_in(a1_wr[861]),  .coef_in(coef[698]), .rdup_out(a2_wr[349]), .rdlo_out(a2_wr[861]));
			radix2 #(.width(width)) rd_st1_350  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[350]), .rdlo_in(a1_wr[862]),  .coef_in(coef[700]), .rdup_out(a2_wr[350]), .rdlo_out(a2_wr[862]));
			radix2 #(.width(width)) rd_st1_351  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[351]), .rdlo_in(a1_wr[863]),  .coef_in(coef[702]), .rdup_out(a2_wr[351]), .rdlo_out(a2_wr[863]));
			radix2 #(.width(width)) rd_st1_352  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[352]), .rdlo_in(a1_wr[864]),  .coef_in(coef[704]), .rdup_out(a2_wr[352]), .rdlo_out(a2_wr[864]));
			radix2 #(.width(width)) rd_st1_353  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[353]), .rdlo_in(a1_wr[865]),  .coef_in(coef[706]), .rdup_out(a2_wr[353]), .rdlo_out(a2_wr[865]));
			radix2 #(.width(width)) rd_st1_354  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[354]), .rdlo_in(a1_wr[866]),  .coef_in(coef[708]), .rdup_out(a2_wr[354]), .rdlo_out(a2_wr[866]));
			radix2 #(.width(width)) rd_st1_355  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[355]), .rdlo_in(a1_wr[867]),  .coef_in(coef[710]), .rdup_out(a2_wr[355]), .rdlo_out(a2_wr[867]));
			radix2 #(.width(width)) rd_st1_356  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[356]), .rdlo_in(a1_wr[868]),  .coef_in(coef[712]), .rdup_out(a2_wr[356]), .rdlo_out(a2_wr[868]));
			radix2 #(.width(width)) rd_st1_357  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[357]), .rdlo_in(a1_wr[869]),  .coef_in(coef[714]), .rdup_out(a2_wr[357]), .rdlo_out(a2_wr[869]));
			radix2 #(.width(width)) rd_st1_358  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[358]), .rdlo_in(a1_wr[870]),  .coef_in(coef[716]), .rdup_out(a2_wr[358]), .rdlo_out(a2_wr[870]));
			radix2 #(.width(width)) rd_st1_359  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[359]), .rdlo_in(a1_wr[871]),  .coef_in(coef[718]), .rdup_out(a2_wr[359]), .rdlo_out(a2_wr[871]));
			radix2 #(.width(width)) rd_st1_360  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[360]), .rdlo_in(a1_wr[872]),  .coef_in(coef[720]), .rdup_out(a2_wr[360]), .rdlo_out(a2_wr[872]));
			radix2 #(.width(width)) rd_st1_361  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[361]), .rdlo_in(a1_wr[873]),  .coef_in(coef[722]), .rdup_out(a2_wr[361]), .rdlo_out(a2_wr[873]));
			radix2 #(.width(width)) rd_st1_362  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[362]), .rdlo_in(a1_wr[874]),  .coef_in(coef[724]), .rdup_out(a2_wr[362]), .rdlo_out(a2_wr[874]));
			radix2 #(.width(width)) rd_st1_363  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[363]), .rdlo_in(a1_wr[875]),  .coef_in(coef[726]), .rdup_out(a2_wr[363]), .rdlo_out(a2_wr[875]));
			radix2 #(.width(width)) rd_st1_364  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[364]), .rdlo_in(a1_wr[876]),  .coef_in(coef[728]), .rdup_out(a2_wr[364]), .rdlo_out(a2_wr[876]));
			radix2 #(.width(width)) rd_st1_365  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[365]), .rdlo_in(a1_wr[877]),  .coef_in(coef[730]), .rdup_out(a2_wr[365]), .rdlo_out(a2_wr[877]));
			radix2 #(.width(width)) rd_st1_366  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[366]), .rdlo_in(a1_wr[878]),  .coef_in(coef[732]), .rdup_out(a2_wr[366]), .rdlo_out(a2_wr[878]));
			radix2 #(.width(width)) rd_st1_367  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[367]), .rdlo_in(a1_wr[879]),  .coef_in(coef[734]), .rdup_out(a2_wr[367]), .rdlo_out(a2_wr[879]));
			radix2 #(.width(width)) rd_st1_368  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[368]), .rdlo_in(a1_wr[880]),  .coef_in(coef[736]), .rdup_out(a2_wr[368]), .rdlo_out(a2_wr[880]));
			radix2 #(.width(width)) rd_st1_369  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[369]), .rdlo_in(a1_wr[881]),  .coef_in(coef[738]), .rdup_out(a2_wr[369]), .rdlo_out(a2_wr[881]));
			radix2 #(.width(width)) rd_st1_370  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[370]), .rdlo_in(a1_wr[882]),  .coef_in(coef[740]), .rdup_out(a2_wr[370]), .rdlo_out(a2_wr[882]));
			radix2 #(.width(width)) rd_st1_371  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[371]), .rdlo_in(a1_wr[883]),  .coef_in(coef[742]), .rdup_out(a2_wr[371]), .rdlo_out(a2_wr[883]));
			radix2 #(.width(width)) rd_st1_372  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[372]), .rdlo_in(a1_wr[884]),  .coef_in(coef[744]), .rdup_out(a2_wr[372]), .rdlo_out(a2_wr[884]));
			radix2 #(.width(width)) rd_st1_373  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[373]), .rdlo_in(a1_wr[885]),  .coef_in(coef[746]), .rdup_out(a2_wr[373]), .rdlo_out(a2_wr[885]));
			radix2 #(.width(width)) rd_st1_374  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[374]), .rdlo_in(a1_wr[886]),  .coef_in(coef[748]), .rdup_out(a2_wr[374]), .rdlo_out(a2_wr[886]));
			radix2 #(.width(width)) rd_st1_375  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[375]), .rdlo_in(a1_wr[887]),  .coef_in(coef[750]), .rdup_out(a2_wr[375]), .rdlo_out(a2_wr[887]));
			radix2 #(.width(width)) rd_st1_376  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[376]), .rdlo_in(a1_wr[888]),  .coef_in(coef[752]), .rdup_out(a2_wr[376]), .rdlo_out(a2_wr[888]));
			radix2 #(.width(width)) rd_st1_377  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[377]), .rdlo_in(a1_wr[889]),  .coef_in(coef[754]), .rdup_out(a2_wr[377]), .rdlo_out(a2_wr[889]));
			radix2 #(.width(width)) rd_st1_378  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[378]), .rdlo_in(a1_wr[890]),  .coef_in(coef[756]), .rdup_out(a2_wr[378]), .rdlo_out(a2_wr[890]));
			radix2 #(.width(width)) rd_st1_379  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[379]), .rdlo_in(a1_wr[891]),  .coef_in(coef[758]), .rdup_out(a2_wr[379]), .rdlo_out(a2_wr[891]));
			radix2 #(.width(width)) rd_st1_380  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[380]), .rdlo_in(a1_wr[892]),  .coef_in(coef[760]), .rdup_out(a2_wr[380]), .rdlo_out(a2_wr[892]));
			radix2 #(.width(width)) rd_st1_381  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[381]), .rdlo_in(a1_wr[893]),  .coef_in(coef[762]), .rdup_out(a2_wr[381]), .rdlo_out(a2_wr[893]));
			radix2 #(.width(width)) rd_st1_382  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[382]), .rdlo_in(a1_wr[894]),  .coef_in(coef[764]), .rdup_out(a2_wr[382]), .rdlo_out(a2_wr[894]));
			radix2 #(.width(width)) rd_st1_383  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[383]), .rdlo_in(a1_wr[895]),  .coef_in(coef[766]), .rdup_out(a2_wr[383]), .rdlo_out(a2_wr[895]));
			radix2 #(.width(width)) rd_st1_384  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[384]), .rdlo_in(a1_wr[896]),  .coef_in(coef[768]), .rdup_out(a2_wr[384]), .rdlo_out(a2_wr[896]));
			radix2 #(.width(width)) rd_st1_385  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[385]), .rdlo_in(a1_wr[897]),  .coef_in(coef[770]), .rdup_out(a2_wr[385]), .rdlo_out(a2_wr[897]));
			radix2 #(.width(width)) rd_st1_386  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[386]), .rdlo_in(a1_wr[898]),  .coef_in(coef[772]), .rdup_out(a2_wr[386]), .rdlo_out(a2_wr[898]));
			radix2 #(.width(width)) rd_st1_387  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[387]), .rdlo_in(a1_wr[899]),  .coef_in(coef[774]), .rdup_out(a2_wr[387]), .rdlo_out(a2_wr[899]));
			radix2 #(.width(width)) rd_st1_388  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[388]), .rdlo_in(a1_wr[900]),  .coef_in(coef[776]), .rdup_out(a2_wr[388]), .rdlo_out(a2_wr[900]));
			radix2 #(.width(width)) rd_st1_389  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[389]), .rdlo_in(a1_wr[901]),  .coef_in(coef[778]), .rdup_out(a2_wr[389]), .rdlo_out(a2_wr[901]));
			radix2 #(.width(width)) rd_st1_390  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[390]), .rdlo_in(a1_wr[902]),  .coef_in(coef[780]), .rdup_out(a2_wr[390]), .rdlo_out(a2_wr[902]));
			radix2 #(.width(width)) rd_st1_391  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[391]), .rdlo_in(a1_wr[903]),  .coef_in(coef[782]), .rdup_out(a2_wr[391]), .rdlo_out(a2_wr[903]));
			radix2 #(.width(width)) rd_st1_392  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[392]), .rdlo_in(a1_wr[904]),  .coef_in(coef[784]), .rdup_out(a2_wr[392]), .rdlo_out(a2_wr[904]));
			radix2 #(.width(width)) rd_st1_393  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[393]), .rdlo_in(a1_wr[905]),  .coef_in(coef[786]), .rdup_out(a2_wr[393]), .rdlo_out(a2_wr[905]));
			radix2 #(.width(width)) rd_st1_394  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[394]), .rdlo_in(a1_wr[906]),  .coef_in(coef[788]), .rdup_out(a2_wr[394]), .rdlo_out(a2_wr[906]));
			radix2 #(.width(width)) rd_st1_395  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[395]), .rdlo_in(a1_wr[907]),  .coef_in(coef[790]), .rdup_out(a2_wr[395]), .rdlo_out(a2_wr[907]));
			radix2 #(.width(width)) rd_st1_396  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[396]), .rdlo_in(a1_wr[908]),  .coef_in(coef[792]), .rdup_out(a2_wr[396]), .rdlo_out(a2_wr[908]));
			radix2 #(.width(width)) rd_st1_397  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[397]), .rdlo_in(a1_wr[909]),  .coef_in(coef[794]), .rdup_out(a2_wr[397]), .rdlo_out(a2_wr[909]));
			radix2 #(.width(width)) rd_st1_398  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[398]), .rdlo_in(a1_wr[910]),  .coef_in(coef[796]), .rdup_out(a2_wr[398]), .rdlo_out(a2_wr[910]));
			radix2 #(.width(width)) rd_st1_399  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[399]), .rdlo_in(a1_wr[911]),  .coef_in(coef[798]), .rdup_out(a2_wr[399]), .rdlo_out(a2_wr[911]));
			radix2 #(.width(width)) rd_st1_400  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[400]), .rdlo_in(a1_wr[912]),  .coef_in(coef[800]), .rdup_out(a2_wr[400]), .rdlo_out(a2_wr[912]));
			radix2 #(.width(width)) rd_st1_401  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[401]), .rdlo_in(a1_wr[913]),  .coef_in(coef[802]), .rdup_out(a2_wr[401]), .rdlo_out(a2_wr[913]));
			radix2 #(.width(width)) rd_st1_402  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[402]), .rdlo_in(a1_wr[914]),  .coef_in(coef[804]), .rdup_out(a2_wr[402]), .rdlo_out(a2_wr[914]));
			radix2 #(.width(width)) rd_st1_403  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[403]), .rdlo_in(a1_wr[915]),  .coef_in(coef[806]), .rdup_out(a2_wr[403]), .rdlo_out(a2_wr[915]));
			radix2 #(.width(width)) rd_st1_404  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[404]), .rdlo_in(a1_wr[916]),  .coef_in(coef[808]), .rdup_out(a2_wr[404]), .rdlo_out(a2_wr[916]));
			radix2 #(.width(width)) rd_st1_405  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[405]), .rdlo_in(a1_wr[917]),  .coef_in(coef[810]), .rdup_out(a2_wr[405]), .rdlo_out(a2_wr[917]));
			radix2 #(.width(width)) rd_st1_406  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[406]), .rdlo_in(a1_wr[918]),  .coef_in(coef[812]), .rdup_out(a2_wr[406]), .rdlo_out(a2_wr[918]));
			radix2 #(.width(width)) rd_st1_407  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[407]), .rdlo_in(a1_wr[919]),  .coef_in(coef[814]), .rdup_out(a2_wr[407]), .rdlo_out(a2_wr[919]));
			radix2 #(.width(width)) rd_st1_408  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[408]), .rdlo_in(a1_wr[920]),  .coef_in(coef[816]), .rdup_out(a2_wr[408]), .rdlo_out(a2_wr[920]));
			radix2 #(.width(width)) rd_st1_409  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[409]), .rdlo_in(a1_wr[921]),  .coef_in(coef[818]), .rdup_out(a2_wr[409]), .rdlo_out(a2_wr[921]));
			radix2 #(.width(width)) rd_st1_410  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[410]), .rdlo_in(a1_wr[922]),  .coef_in(coef[820]), .rdup_out(a2_wr[410]), .rdlo_out(a2_wr[922]));
			radix2 #(.width(width)) rd_st1_411  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[411]), .rdlo_in(a1_wr[923]),  .coef_in(coef[822]), .rdup_out(a2_wr[411]), .rdlo_out(a2_wr[923]));
			radix2 #(.width(width)) rd_st1_412  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[412]), .rdlo_in(a1_wr[924]),  .coef_in(coef[824]), .rdup_out(a2_wr[412]), .rdlo_out(a2_wr[924]));
			radix2 #(.width(width)) rd_st1_413  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[413]), .rdlo_in(a1_wr[925]),  .coef_in(coef[826]), .rdup_out(a2_wr[413]), .rdlo_out(a2_wr[925]));
			radix2 #(.width(width)) rd_st1_414  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[414]), .rdlo_in(a1_wr[926]),  .coef_in(coef[828]), .rdup_out(a2_wr[414]), .rdlo_out(a2_wr[926]));
			radix2 #(.width(width)) rd_st1_415  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[415]), .rdlo_in(a1_wr[927]),  .coef_in(coef[830]), .rdup_out(a2_wr[415]), .rdlo_out(a2_wr[927]));
			radix2 #(.width(width)) rd_st1_416  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[416]), .rdlo_in(a1_wr[928]),  .coef_in(coef[832]), .rdup_out(a2_wr[416]), .rdlo_out(a2_wr[928]));
			radix2 #(.width(width)) rd_st1_417  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[417]), .rdlo_in(a1_wr[929]),  .coef_in(coef[834]), .rdup_out(a2_wr[417]), .rdlo_out(a2_wr[929]));
			radix2 #(.width(width)) rd_st1_418  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[418]), .rdlo_in(a1_wr[930]),  .coef_in(coef[836]), .rdup_out(a2_wr[418]), .rdlo_out(a2_wr[930]));
			radix2 #(.width(width)) rd_st1_419  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[419]), .rdlo_in(a1_wr[931]),  .coef_in(coef[838]), .rdup_out(a2_wr[419]), .rdlo_out(a2_wr[931]));
			radix2 #(.width(width)) rd_st1_420  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[420]), .rdlo_in(a1_wr[932]),  .coef_in(coef[840]), .rdup_out(a2_wr[420]), .rdlo_out(a2_wr[932]));
			radix2 #(.width(width)) rd_st1_421  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[421]), .rdlo_in(a1_wr[933]),  .coef_in(coef[842]), .rdup_out(a2_wr[421]), .rdlo_out(a2_wr[933]));
			radix2 #(.width(width)) rd_st1_422  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[422]), .rdlo_in(a1_wr[934]),  .coef_in(coef[844]), .rdup_out(a2_wr[422]), .rdlo_out(a2_wr[934]));
			radix2 #(.width(width)) rd_st1_423  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[423]), .rdlo_in(a1_wr[935]),  .coef_in(coef[846]), .rdup_out(a2_wr[423]), .rdlo_out(a2_wr[935]));
			radix2 #(.width(width)) rd_st1_424  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[424]), .rdlo_in(a1_wr[936]),  .coef_in(coef[848]), .rdup_out(a2_wr[424]), .rdlo_out(a2_wr[936]));
			radix2 #(.width(width)) rd_st1_425  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[425]), .rdlo_in(a1_wr[937]),  .coef_in(coef[850]), .rdup_out(a2_wr[425]), .rdlo_out(a2_wr[937]));
			radix2 #(.width(width)) rd_st1_426  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[426]), .rdlo_in(a1_wr[938]),  .coef_in(coef[852]), .rdup_out(a2_wr[426]), .rdlo_out(a2_wr[938]));
			radix2 #(.width(width)) rd_st1_427  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[427]), .rdlo_in(a1_wr[939]),  .coef_in(coef[854]), .rdup_out(a2_wr[427]), .rdlo_out(a2_wr[939]));
			radix2 #(.width(width)) rd_st1_428  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[428]), .rdlo_in(a1_wr[940]),  .coef_in(coef[856]), .rdup_out(a2_wr[428]), .rdlo_out(a2_wr[940]));
			radix2 #(.width(width)) rd_st1_429  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[429]), .rdlo_in(a1_wr[941]),  .coef_in(coef[858]), .rdup_out(a2_wr[429]), .rdlo_out(a2_wr[941]));
			radix2 #(.width(width)) rd_st1_430  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[430]), .rdlo_in(a1_wr[942]),  .coef_in(coef[860]), .rdup_out(a2_wr[430]), .rdlo_out(a2_wr[942]));
			radix2 #(.width(width)) rd_st1_431  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[431]), .rdlo_in(a1_wr[943]),  .coef_in(coef[862]), .rdup_out(a2_wr[431]), .rdlo_out(a2_wr[943]));
			radix2 #(.width(width)) rd_st1_432  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[432]), .rdlo_in(a1_wr[944]),  .coef_in(coef[864]), .rdup_out(a2_wr[432]), .rdlo_out(a2_wr[944]));
			radix2 #(.width(width)) rd_st1_433  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[433]), .rdlo_in(a1_wr[945]),  .coef_in(coef[866]), .rdup_out(a2_wr[433]), .rdlo_out(a2_wr[945]));
			radix2 #(.width(width)) rd_st1_434  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[434]), .rdlo_in(a1_wr[946]),  .coef_in(coef[868]), .rdup_out(a2_wr[434]), .rdlo_out(a2_wr[946]));
			radix2 #(.width(width)) rd_st1_435  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[435]), .rdlo_in(a1_wr[947]),  .coef_in(coef[870]), .rdup_out(a2_wr[435]), .rdlo_out(a2_wr[947]));
			radix2 #(.width(width)) rd_st1_436  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[436]), .rdlo_in(a1_wr[948]),  .coef_in(coef[872]), .rdup_out(a2_wr[436]), .rdlo_out(a2_wr[948]));
			radix2 #(.width(width)) rd_st1_437  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[437]), .rdlo_in(a1_wr[949]),  .coef_in(coef[874]), .rdup_out(a2_wr[437]), .rdlo_out(a2_wr[949]));
			radix2 #(.width(width)) rd_st1_438  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[438]), .rdlo_in(a1_wr[950]),  .coef_in(coef[876]), .rdup_out(a2_wr[438]), .rdlo_out(a2_wr[950]));
			radix2 #(.width(width)) rd_st1_439  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[439]), .rdlo_in(a1_wr[951]),  .coef_in(coef[878]), .rdup_out(a2_wr[439]), .rdlo_out(a2_wr[951]));
			radix2 #(.width(width)) rd_st1_440  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[440]), .rdlo_in(a1_wr[952]),  .coef_in(coef[880]), .rdup_out(a2_wr[440]), .rdlo_out(a2_wr[952]));
			radix2 #(.width(width)) rd_st1_441  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[441]), .rdlo_in(a1_wr[953]),  .coef_in(coef[882]), .rdup_out(a2_wr[441]), .rdlo_out(a2_wr[953]));
			radix2 #(.width(width)) rd_st1_442  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[442]), .rdlo_in(a1_wr[954]),  .coef_in(coef[884]), .rdup_out(a2_wr[442]), .rdlo_out(a2_wr[954]));
			radix2 #(.width(width)) rd_st1_443  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[443]), .rdlo_in(a1_wr[955]),  .coef_in(coef[886]), .rdup_out(a2_wr[443]), .rdlo_out(a2_wr[955]));
			radix2 #(.width(width)) rd_st1_444  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[444]), .rdlo_in(a1_wr[956]),  .coef_in(coef[888]), .rdup_out(a2_wr[444]), .rdlo_out(a2_wr[956]));
			radix2 #(.width(width)) rd_st1_445  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[445]), .rdlo_in(a1_wr[957]),  .coef_in(coef[890]), .rdup_out(a2_wr[445]), .rdlo_out(a2_wr[957]));
			radix2 #(.width(width)) rd_st1_446  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[446]), .rdlo_in(a1_wr[958]),  .coef_in(coef[892]), .rdup_out(a2_wr[446]), .rdlo_out(a2_wr[958]));
			radix2 #(.width(width)) rd_st1_447  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[447]), .rdlo_in(a1_wr[959]),  .coef_in(coef[894]), .rdup_out(a2_wr[447]), .rdlo_out(a2_wr[959]));
			radix2 #(.width(width)) rd_st1_448  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[448]), .rdlo_in(a1_wr[960]),  .coef_in(coef[896]), .rdup_out(a2_wr[448]), .rdlo_out(a2_wr[960]));
			radix2 #(.width(width)) rd_st1_449  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[449]), .rdlo_in(a1_wr[961]),  .coef_in(coef[898]), .rdup_out(a2_wr[449]), .rdlo_out(a2_wr[961]));
			radix2 #(.width(width)) rd_st1_450  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[450]), .rdlo_in(a1_wr[962]),  .coef_in(coef[900]), .rdup_out(a2_wr[450]), .rdlo_out(a2_wr[962]));
			radix2 #(.width(width)) rd_st1_451  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[451]), .rdlo_in(a1_wr[963]),  .coef_in(coef[902]), .rdup_out(a2_wr[451]), .rdlo_out(a2_wr[963]));
			radix2 #(.width(width)) rd_st1_452  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[452]), .rdlo_in(a1_wr[964]),  .coef_in(coef[904]), .rdup_out(a2_wr[452]), .rdlo_out(a2_wr[964]));
			radix2 #(.width(width)) rd_st1_453  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[453]), .rdlo_in(a1_wr[965]),  .coef_in(coef[906]), .rdup_out(a2_wr[453]), .rdlo_out(a2_wr[965]));
			radix2 #(.width(width)) rd_st1_454  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[454]), .rdlo_in(a1_wr[966]),  .coef_in(coef[908]), .rdup_out(a2_wr[454]), .rdlo_out(a2_wr[966]));
			radix2 #(.width(width)) rd_st1_455  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[455]), .rdlo_in(a1_wr[967]),  .coef_in(coef[910]), .rdup_out(a2_wr[455]), .rdlo_out(a2_wr[967]));
			radix2 #(.width(width)) rd_st1_456  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[456]), .rdlo_in(a1_wr[968]),  .coef_in(coef[912]), .rdup_out(a2_wr[456]), .rdlo_out(a2_wr[968]));
			radix2 #(.width(width)) rd_st1_457  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[457]), .rdlo_in(a1_wr[969]),  .coef_in(coef[914]), .rdup_out(a2_wr[457]), .rdlo_out(a2_wr[969]));
			radix2 #(.width(width)) rd_st1_458  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[458]), .rdlo_in(a1_wr[970]),  .coef_in(coef[916]), .rdup_out(a2_wr[458]), .rdlo_out(a2_wr[970]));
			radix2 #(.width(width)) rd_st1_459  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[459]), .rdlo_in(a1_wr[971]),  .coef_in(coef[918]), .rdup_out(a2_wr[459]), .rdlo_out(a2_wr[971]));
			radix2 #(.width(width)) rd_st1_460  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[460]), .rdlo_in(a1_wr[972]),  .coef_in(coef[920]), .rdup_out(a2_wr[460]), .rdlo_out(a2_wr[972]));
			radix2 #(.width(width)) rd_st1_461  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[461]), .rdlo_in(a1_wr[973]),  .coef_in(coef[922]), .rdup_out(a2_wr[461]), .rdlo_out(a2_wr[973]));
			radix2 #(.width(width)) rd_st1_462  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[462]), .rdlo_in(a1_wr[974]),  .coef_in(coef[924]), .rdup_out(a2_wr[462]), .rdlo_out(a2_wr[974]));
			radix2 #(.width(width)) rd_st1_463  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[463]), .rdlo_in(a1_wr[975]),  .coef_in(coef[926]), .rdup_out(a2_wr[463]), .rdlo_out(a2_wr[975]));
			radix2 #(.width(width)) rd_st1_464  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[464]), .rdlo_in(a1_wr[976]),  .coef_in(coef[928]), .rdup_out(a2_wr[464]), .rdlo_out(a2_wr[976]));
			radix2 #(.width(width)) rd_st1_465  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[465]), .rdlo_in(a1_wr[977]),  .coef_in(coef[930]), .rdup_out(a2_wr[465]), .rdlo_out(a2_wr[977]));
			radix2 #(.width(width)) rd_st1_466  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[466]), .rdlo_in(a1_wr[978]),  .coef_in(coef[932]), .rdup_out(a2_wr[466]), .rdlo_out(a2_wr[978]));
			radix2 #(.width(width)) rd_st1_467  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[467]), .rdlo_in(a1_wr[979]),  .coef_in(coef[934]), .rdup_out(a2_wr[467]), .rdlo_out(a2_wr[979]));
			radix2 #(.width(width)) rd_st1_468  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[468]), .rdlo_in(a1_wr[980]),  .coef_in(coef[936]), .rdup_out(a2_wr[468]), .rdlo_out(a2_wr[980]));
			radix2 #(.width(width)) rd_st1_469  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[469]), .rdlo_in(a1_wr[981]),  .coef_in(coef[938]), .rdup_out(a2_wr[469]), .rdlo_out(a2_wr[981]));
			radix2 #(.width(width)) rd_st1_470  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[470]), .rdlo_in(a1_wr[982]),  .coef_in(coef[940]), .rdup_out(a2_wr[470]), .rdlo_out(a2_wr[982]));
			radix2 #(.width(width)) rd_st1_471  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[471]), .rdlo_in(a1_wr[983]),  .coef_in(coef[942]), .rdup_out(a2_wr[471]), .rdlo_out(a2_wr[983]));
			radix2 #(.width(width)) rd_st1_472  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[472]), .rdlo_in(a1_wr[984]),  .coef_in(coef[944]), .rdup_out(a2_wr[472]), .rdlo_out(a2_wr[984]));
			radix2 #(.width(width)) rd_st1_473  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[473]), .rdlo_in(a1_wr[985]),  .coef_in(coef[946]), .rdup_out(a2_wr[473]), .rdlo_out(a2_wr[985]));
			radix2 #(.width(width)) rd_st1_474  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[474]), .rdlo_in(a1_wr[986]),  .coef_in(coef[948]), .rdup_out(a2_wr[474]), .rdlo_out(a2_wr[986]));
			radix2 #(.width(width)) rd_st1_475  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[475]), .rdlo_in(a1_wr[987]),  .coef_in(coef[950]), .rdup_out(a2_wr[475]), .rdlo_out(a2_wr[987]));
			radix2 #(.width(width)) rd_st1_476  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[476]), .rdlo_in(a1_wr[988]),  .coef_in(coef[952]), .rdup_out(a2_wr[476]), .rdlo_out(a2_wr[988]));
			radix2 #(.width(width)) rd_st1_477  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[477]), .rdlo_in(a1_wr[989]),  .coef_in(coef[954]), .rdup_out(a2_wr[477]), .rdlo_out(a2_wr[989]));
			radix2 #(.width(width)) rd_st1_478  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[478]), .rdlo_in(a1_wr[990]),  .coef_in(coef[956]), .rdup_out(a2_wr[478]), .rdlo_out(a2_wr[990]));
			radix2 #(.width(width)) rd_st1_479  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[479]), .rdlo_in(a1_wr[991]),  .coef_in(coef[958]), .rdup_out(a2_wr[479]), .rdlo_out(a2_wr[991]));
			radix2 #(.width(width)) rd_st1_480  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[480]), .rdlo_in(a1_wr[992]),  .coef_in(coef[960]), .rdup_out(a2_wr[480]), .rdlo_out(a2_wr[992]));
			radix2 #(.width(width)) rd_st1_481  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[481]), .rdlo_in(a1_wr[993]),  .coef_in(coef[962]), .rdup_out(a2_wr[481]), .rdlo_out(a2_wr[993]));
			radix2 #(.width(width)) rd_st1_482  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[482]), .rdlo_in(a1_wr[994]),  .coef_in(coef[964]), .rdup_out(a2_wr[482]), .rdlo_out(a2_wr[994]));
			radix2 #(.width(width)) rd_st1_483  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[483]), .rdlo_in(a1_wr[995]),  .coef_in(coef[966]), .rdup_out(a2_wr[483]), .rdlo_out(a2_wr[995]));
			radix2 #(.width(width)) rd_st1_484  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[484]), .rdlo_in(a1_wr[996]),  .coef_in(coef[968]), .rdup_out(a2_wr[484]), .rdlo_out(a2_wr[996]));
			radix2 #(.width(width)) rd_st1_485  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[485]), .rdlo_in(a1_wr[997]),  .coef_in(coef[970]), .rdup_out(a2_wr[485]), .rdlo_out(a2_wr[997]));
			radix2 #(.width(width)) rd_st1_486  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[486]), .rdlo_in(a1_wr[998]),  .coef_in(coef[972]), .rdup_out(a2_wr[486]), .rdlo_out(a2_wr[998]));
			radix2 #(.width(width)) rd_st1_487  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[487]), .rdlo_in(a1_wr[999]),  .coef_in(coef[974]), .rdup_out(a2_wr[487]), .rdlo_out(a2_wr[999]));
			radix2 #(.width(width)) rd_st1_488  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[488]), .rdlo_in(a1_wr[1000]),  .coef_in(coef[976]), .rdup_out(a2_wr[488]), .rdlo_out(a2_wr[1000]));
			radix2 #(.width(width)) rd_st1_489  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[489]), .rdlo_in(a1_wr[1001]),  .coef_in(coef[978]), .rdup_out(a2_wr[489]), .rdlo_out(a2_wr[1001]));
			radix2 #(.width(width)) rd_st1_490  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[490]), .rdlo_in(a1_wr[1002]),  .coef_in(coef[980]), .rdup_out(a2_wr[490]), .rdlo_out(a2_wr[1002]));
			radix2 #(.width(width)) rd_st1_491  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[491]), .rdlo_in(a1_wr[1003]),  .coef_in(coef[982]), .rdup_out(a2_wr[491]), .rdlo_out(a2_wr[1003]));
			radix2 #(.width(width)) rd_st1_492  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[492]), .rdlo_in(a1_wr[1004]),  .coef_in(coef[984]), .rdup_out(a2_wr[492]), .rdlo_out(a2_wr[1004]));
			radix2 #(.width(width)) rd_st1_493  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[493]), .rdlo_in(a1_wr[1005]),  .coef_in(coef[986]), .rdup_out(a2_wr[493]), .rdlo_out(a2_wr[1005]));
			radix2 #(.width(width)) rd_st1_494  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[494]), .rdlo_in(a1_wr[1006]),  .coef_in(coef[988]), .rdup_out(a2_wr[494]), .rdlo_out(a2_wr[1006]));
			radix2 #(.width(width)) rd_st1_495  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[495]), .rdlo_in(a1_wr[1007]),  .coef_in(coef[990]), .rdup_out(a2_wr[495]), .rdlo_out(a2_wr[1007]));
			radix2 #(.width(width)) rd_st1_496  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[496]), .rdlo_in(a1_wr[1008]),  .coef_in(coef[992]), .rdup_out(a2_wr[496]), .rdlo_out(a2_wr[1008]));
			radix2 #(.width(width)) rd_st1_497  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[497]), .rdlo_in(a1_wr[1009]),  .coef_in(coef[994]), .rdup_out(a2_wr[497]), .rdlo_out(a2_wr[1009]));
			radix2 #(.width(width)) rd_st1_498  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[498]), .rdlo_in(a1_wr[1010]),  .coef_in(coef[996]), .rdup_out(a2_wr[498]), .rdlo_out(a2_wr[1010]));
			radix2 #(.width(width)) rd_st1_499  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[499]), .rdlo_in(a1_wr[1011]),  .coef_in(coef[998]), .rdup_out(a2_wr[499]), .rdlo_out(a2_wr[1011]));
			radix2 #(.width(width)) rd_st1_500  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[500]), .rdlo_in(a1_wr[1012]),  .coef_in(coef[1000]), .rdup_out(a2_wr[500]), .rdlo_out(a2_wr[1012]));
			radix2 #(.width(width)) rd_st1_501  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[501]), .rdlo_in(a1_wr[1013]),  .coef_in(coef[1002]), .rdup_out(a2_wr[501]), .rdlo_out(a2_wr[1013]));
			radix2 #(.width(width)) rd_st1_502  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[502]), .rdlo_in(a1_wr[1014]),  .coef_in(coef[1004]), .rdup_out(a2_wr[502]), .rdlo_out(a2_wr[1014]));
			radix2 #(.width(width)) rd_st1_503  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[503]), .rdlo_in(a1_wr[1015]),  .coef_in(coef[1006]), .rdup_out(a2_wr[503]), .rdlo_out(a2_wr[1015]));
			radix2 #(.width(width)) rd_st1_504  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[504]), .rdlo_in(a1_wr[1016]),  .coef_in(coef[1008]), .rdup_out(a2_wr[504]), .rdlo_out(a2_wr[1016]));
			radix2 #(.width(width)) rd_st1_505  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[505]), .rdlo_in(a1_wr[1017]),  .coef_in(coef[1010]), .rdup_out(a2_wr[505]), .rdlo_out(a2_wr[1017]));
			radix2 #(.width(width)) rd_st1_506  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[506]), .rdlo_in(a1_wr[1018]),  .coef_in(coef[1012]), .rdup_out(a2_wr[506]), .rdlo_out(a2_wr[1018]));
			radix2 #(.width(width)) rd_st1_507  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[507]), .rdlo_in(a1_wr[1019]),  .coef_in(coef[1014]), .rdup_out(a2_wr[507]), .rdlo_out(a2_wr[1019]));
			radix2 #(.width(width)) rd_st1_508  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[508]), .rdlo_in(a1_wr[1020]),  .coef_in(coef[1016]), .rdup_out(a2_wr[508]), .rdlo_out(a2_wr[1020]));
			radix2 #(.width(width)) rd_st1_509  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[509]), .rdlo_in(a1_wr[1021]),  .coef_in(coef[1018]), .rdup_out(a2_wr[509]), .rdlo_out(a2_wr[1021]));
			radix2 #(.width(width)) rd_st1_510  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[510]), .rdlo_in(a1_wr[1022]),  .coef_in(coef[1020]), .rdup_out(a2_wr[510]), .rdlo_out(a2_wr[1022]));
			radix2 #(.width(width)) rd_st1_511  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[511]), .rdlo_in(a1_wr[1023]),  .coef_in(coef[1022]), .rdup_out(a2_wr[511]), .rdlo_out(a2_wr[1023]));
			radix2 #(.width(width)) rd_st1_1024  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1024]), .rdlo_in(a1_wr[1536]),  .coef_in(coef[0]), .rdup_out(a2_wr[1024]), .rdlo_out(a2_wr[1536]));
			radix2 #(.width(width)) rd_st1_1025  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1025]), .rdlo_in(a1_wr[1537]),  .coef_in(coef[2]), .rdup_out(a2_wr[1025]), .rdlo_out(a2_wr[1537]));
			radix2 #(.width(width)) rd_st1_1026  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1026]), .rdlo_in(a1_wr[1538]),  .coef_in(coef[4]), .rdup_out(a2_wr[1026]), .rdlo_out(a2_wr[1538]));
			radix2 #(.width(width)) rd_st1_1027  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1027]), .rdlo_in(a1_wr[1539]),  .coef_in(coef[6]), .rdup_out(a2_wr[1027]), .rdlo_out(a2_wr[1539]));
			radix2 #(.width(width)) rd_st1_1028  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1028]), .rdlo_in(a1_wr[1540]),  .coef_in(coef[8]), .rdup_out(a2_wr[1028]), .rdlo_out(a2_wr[1540]));
			radix2 #(.width(width)) rd_st1_1029  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1029]), .rdlo_in(a1_wr[1541]),  .coef_in(coef[10]), .rdup_out(a2_wr[1029]), .rdlo_out(a2_wr[1541]));
			radix2 #(.width(width)) rd_st1_1030  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1030]), .rdlo_in(a1_wr[1542]),  .coef_in(coef[12]), .rdup_out(a2_wr[1030]), .rdlo_out(a2_wr[1542]));
			radix2 #(.width(width)) rd_st1_1031  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1031]), .rdlo_in(a1_wr[1543]),  .coef_in(coef[14]), .rdup_out(a2_wr[1031]), .rdlo_out(a2_wr[1543]));
			radix2 #(.width(width)) rd_st1_1032  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1032]), .rdlo_in(a1_wr[1544]),  .coef_in(coef[16]), .rdup_out(a2_wr[1032]), .rdlo_out(a2_wr[1544]));
			radix2 #(.width(width)) rd_st1_1033  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1033]), .rdlo_in(a1_wr[1545]),  .coef_in(coef[18]), .rdup_out(a2_wr[1033]), .rdlo_out(a2_wr[1545]));
			radix2 #(.width(width)) rd_st1_1034  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1034]), .rdlo_in(a1_wr[1546]),  .coef_in(coef[20]), .rdup_out(a2_wr[1034]), .rdlo_out(a2_wr[1546]));
			radix2 #(.width(width)) rd_st1_1035  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1035]), .rdlo_in(a1_wr[1547]),  .coef_in(coef[22]), .rdup_out(a2_wr[1035]), .rdlo_out(a2_wr[1547]));
			radix2 #(.width(width)) rd_st1_1036  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1036]), .rdlo_in(a1_wr[1548]),  .coef_in(coef[24]), .rdup_out(a2_wr[1036]), .rdlo_out(a2_wr[1548]));
			radix2 #(.width(width)) rd_st1_1037  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1037]), .rdlo_in(a1_wr[1549]),  .coef_in(coef[26]), .rdup_out(a2_wr[1037]), .rdlo_out(a2_wr[1549]));
			radix2 #(.width(width)) rd_st1_1038  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1038]), .rdlo_in(a1_wr[1550]),  .coef_in(coef[28]), .rdup_out(a2_wr[1038]), .rdlo_out(a2_wr[1550]));
			radix2 #(.width(width)) rd_st1_1039  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1039]), .rdlo_in(a1_wr[1551]),  .coef_in(coef[30]), .rdup_out(a2_wr[1039]), .rdlo_out(a2_wr[1551]));
			radix2 #(.width(width)) rd_st1_1040  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1040]), .rdlo_in(a1_wr[1552]),  .coef_in(coef[32]), .rdup_out(a2_wr[1040]), .rdlo_out(a2_wr[1552]));
			radix2 #(.width(width)) rd_st1_1041  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1041]), .rdlo_in(a1_wr[1553]),  .coef_in(coef[34]), .rdup_out(a2_wr[1041]), .rdlo_out(a2_wr[1553]));
			radix2 #(.width(width)) rd_st1_1042  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1042]), .rdlo_in(a1_wr[1554]),  .coef_in(coef[36]), .rdup_out(a2_wr[1042]), .rdlo_out(a2_wr[1554]));
			radix2 #(.width(width)) rd_st1_1043  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1043]), .rdlo_in(a1_wr[1555]),  .coef_in(coef[38]), .rdup_out(a2_wr[1043]), .rdlo_out(a2_wr[1555]));
			radix2 #(.width(width)) rd_st1_1044  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1044]), .rdlo_in(a1_wr[1556]),  .coef_in(coef[40]), .rdup_out(a2_wr[1044]), .rdlo_out(a2_wr[1556]));
			radix2 #(.width(width)) rd_st1_1045  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1045]), .rdlo_in(a1_wr[1557]),  .coef_in(coef[42]), .rdup_out(a2_wr[1045]), .rdlo_out(a2_wr[1557]));
			radix2 #(.width(width)) rd_st1_1046  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1046]), .rdlo_in(a1_wr[1558]),  .coef_in(coef[44]), .rdup_out(a2_wr[1046]), .rdlo_out(a2_wr[1558]));
			radix2 #(.width(width)) rd_st1_1047  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1047]), .rdlo_in(a1_wr[1559]),  .coef_in(coef[46]), .rdup_out(a2_wr[1047]), .rdlo_out(a2_wr[1559]));
			radix2 #(.width(width)) rd_st1_1048  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1048]), .rdlo_in(a1_wr[1560]),  .coef_in(coef[48]), .rdup_out(a2_wr[1048]), .rdlo_out(a2_wr[1560]));
			radix2 #(.width(width)) rd_st1_1049  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1049]), .rdlo_in(a1_wr[1561]),  .coef_in(coef[50]), .rdup_out(a2_wr[1049]), .rdlo_out(a2_wr[1561]));
			radix2 #(.width(width)) rd_st1_1050  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1050]), .rdlo_in(a1_wr[1562]),  .coef_in(coef[52]), .rdup_out(a2_wr[1050]), .rdlo_out(a2_wr[1562]));
			radix2 #(.width(width)) rd_st1_1051  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1051]), .rdlo_in(a1_wr[1563]),  .coef_in(coef[54]), .rdup_out(a2_wr[1051]), .rdlo_out(a2_wr[1563]));
			radix2 #(.width(width)) rd_st1_1052  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1052]), .rdlo_in(a1_wr[1564]),  .coef_in(coef[56]), .rdup_out(a2_wr[1052]), .rdlo_out(a2_wr[1564]));
			radix2 #(.width(width)) rd_st1_1053  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1053]), .rdlo_in(a1_wr[1565]),  .coef_in(coef[58]), .rdup_out(a2_wr[1053]), .rdlo_out(a2_wr[1565]));
			radix2 #(.width(width)) rd_st1_1054  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1054]), .rdlo_in(a1_wr[1566]),  .coef_in(coef[60]), .rdup_out(a2_wr[1054]), .rdlo_out(a2_wr[1566]));
			radix2 #(.width(width)) rd_st1_1055  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1055]), .rdlo_in(a1_wr[1567]),  .coef_in(coef[62]), .rdup_out(a2_wr[1055]), .rdlo_out(a2_wr[1567]));
			radix2 #(.width(width)) rd_st1_1056  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1056]), .rdlo_in(a1_wr[1568]),  .coef_in(coef[64]), .rdup_out(a2_wr[1056]), .rdlo_out(a2_wr[1568]));
			radix2 #(.width(width)) rd_st1_1057  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1057]), .rdlo_in(a1_wr[1569]),  .coef_in(coef[66]), .rdup_out(a2_wr[1057]), .rdlo_out(a2_wr[1569]));
			radix2 #(.width(width)) rd_st1_1058  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1058]), .rdlo_in(a1_wr[1570]),  .coef_in(coef[68]), .rdup_out(a2_wr[1058]), .rdlo_out(a2_wr[1570]));
			radix2 #(.width(width)) rd_st1_1059  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1059]), .rdlo_in(a1_wr[1571]),  .coef_in(coef[70]), .rdup_out(a2_wr[1059]), .rdlo_out(a2_wr[1571]));
			radix2 #(.width(width)) rd_st1_1060  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1060]), .rdlo_in(a1_wr[1572]),  .coef_in(coef[72]), .rdup_out(a2_wr[1060]), .rdlo_out(a2_wr[1572]));
			radix2 #(.width(width)) rd_st1_1061  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1061]), .rdlo_in(a1_wr[1573]),  .coef_in(coef[74]), .rdup_out(a2_wr[1061]), .rdlo_out(a2_wr[1573]));
			radix2 #(.width(width)) rd_st1_1062  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1062]), .rdlo_in(a1_wr[1574]),  .coef_in(coef[76]), .rdup_out(a2_wr[1062]), .rdlo_out(a2_wr[1574]));
			radix2 #(.width(width)) rd_st1_1063  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1063]), .rdlo_in(a1_wr[1575]),  .coef_in(coef[78]), .rdup_out(a2_wr[1063]), .rdlo_out(a2_wr[1575]));
			radix2 #(.width(width)) rd_st1_1064  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1064]), .rdlo_in(a1_wr[1576]),  .coef_in(coef[80]), .rdup_out(a2_wr[1064]), .rdlo_out(a2_wr[1576]));
			radix2 #(.width(width)) rd_st1_1065  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1065]), .rdlo_in(a1_wr[1577]),  .coef_in(coef[82]), .rdup_out(a2_wr[1065]), .rdlo_out(a2_wr[1577]));
			radix2 #(.width(width)) rd_st1_1066  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1066]), .rdlo_in(a1_wr[1578]),  .coef_in(coef[84]), .rdup_out(a2_wr[1066]), .rdlo_out(a2_wr[1578]));
			radix2 #(.width(width)) rd_st1_1067  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1067]), .rdlo_in(a1_wr[1579]),  .coef_in(coef[86]), .rdup_out(a2_wr[1067]), .rdlo_out(a2_wr[1579]));
			radix2 #(.width(width)) rd_st1_1068  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1068]), .rdlo_in(a1_wr[1580]),  .coef_in(coef[88]), .rdup_out(a2_wr[1068]), .rdlo_out(a2_wr[1580]));
			radix2 #(.width(width)) rd_st1_1069  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1069]), .rdlo_in(a1_wr[1581]),  .coef_in(coef[90]), .rdup_out(a2_wr[1069]), .rdlo_out(a2_wr[1581]));
			radix2 #(.width(width)) rd_st1_1070  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1070]), .rdlo_in(a1_wr[1582]),  .coef_in(coef[92]), .rdup_out(a2_wr[1070]), .rdlo_out(a2_wr[1582]));
			radix2 #(.width(width)) rd_st1_1071  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1071]), .rdlo_in(a1_wr[1583]),  .coef_in(coef[94]), .rdup_out(a2_wr[1071]), .rdlo_out(a2_wr[1583]));
			radix2 #(.width(width)) rd_st1_1072  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1072]), .rdlo_in(a1_wr[1584]),  .coef_in(coef[96]), .rdup_out(a2_wr[1072]), .rdlo_out(a2_wr[1584]));
			radix2 #(.width(width)) rd_st1_1073  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1073]), .rdlo_in(a1_wr[1585]),  .coef_in(coef[98]), .rdup_out(a2_wr[1073]), .rdlo_out(a2_wr[1585]));
			radix2 #(.width(width)) rd_st1_1074  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1074]), .rdlo_in(a1_wr[1586]),  .coef_in(coef[100]), .rdup_out(a2_wr[1074]), .rdlo_out(a2_wr[1586]));
			radix2 #(.width(width)) rd_st1_1075  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1075]), .rdlo_in(a1_wr[1587]),  .coef_in(coef[102]), .rdup_out(a2_wr[1075]), .rdlo_out(a2_wr[1587]));
			radix2 #(.width(width)) rd_st1_1076  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1076]), .rdlo_in(a1_wr[1588]),  .coef_in(coef[104]), .rdup_out(a2_wr[1076]), .rdlo_out(a2_wr[1588]));
			radix2 #(.width(width)) rd_st1_1077  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1077]), .rdlo_in(a1_wr[1589]),  .coef_in(coef[106]), .rdup_out(a2_wr[1077]), .rdlo_out(a2_wr[1589]));
			radix2 #(.width(width)) rd_st1_1078  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1078]), .rdlo_in(a1_wr[1590]),  .coef_in(coef[108]), .rdup_out(a2_wr[1078]), .rdlo_out(a2_wr[1590]));
			radix2 #(.width(width)) rd_st1_1079  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1079]), .rdlo_in(a1_wr[1591]),  .coef_in(coef[110]), .rdup_out(a2_wr[1079]), .rdlo_out(a2_wr[1591]));
			radix2 #(.width(width)) rd_st1_1080  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1080]), .rdlo_in(a1_wr[1592]),  .coef_in(coef[112]), .rdup_out(a2_wr[1080]), .rdlo_out(a2_wr[1592]));
			radix2 #(.width(width)) rd_st1_1081  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1081]), .rdlo_in(a1_wr[1593]),  .coef_in(coef[114]), .rdup_out(a2_wr[1081]), .rdlo_out(a2_wr[1593]));
			radix2 #(.width(width)) rd_st1_1082  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1082]), .rdlo_in(a1_wr[1594]),  .coef_in(coef[116]), .rdup_out(a2_wr[1082]), .rdlo_out(a2_wr[1594]));
			radix2 #(.width(width)) rd_st1_1083  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1083]), .rdlo_in(a1_wr[1595]),  .coef_in(coef[118]), .rdup_out(a2_wr[1083]), .rdlo_out(a2_wr[1595]));
			radix2 #(.width(width)) rd_st1_1084  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1084]), .rdlo_in(a1_wr[1596]),  .coef_in(coef[120]), .rdup_out(a2_wr[1084]), .rdlo_out(a2_wr[1596]));
			radix2 #(.width(width)) rd_st1_1085  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1085]), .rdlo_in(a1_wr[1597]),  .coef_in(coef[122]), .rdup_out(a2_wr[1085]), .rdlo_out(a2_wr[1597]));
			radix2 #(.width(width)) rd_st1_1086  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1086]), .rdlo_in(a1_wr[1598]),  .coef_in(coef[124]), .rdup_out(a2_wr[1086]), .rdlo_out(a2_wr[1598]));
			radix2 #(.width(width)) rd_st1_1087  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1087]), .rdlo_in(a1_wr[1599]),  .coef_in(coef[126]), .rdup_out(a2_wr[1087]), .rdlo_out(a2_wr[1599]));
			radix2 #(.width(width)) rd_st1_1088  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1088]), .rdlo_in(a1_wr[1600]),  .coef_in(coef[128]), .rdup_out(a2_wr[1088]), .rdlo_out(a2_wr[1600]));
			radix2 #(.width(width)) rd_st1_1089  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1089]), .rdlo_in(a1_wr[1601]),  .coef_in(coef[130]), .rdup_out(a2_wr[1089]), .rdlo_out(a2_wr[1601]));
			radix2 #(.width(width)) rd_st1_1090  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1090]), .rdlo_in(a1_wr[1602]),  .coef_in(coef[132]), .rdup_out(a2_wr[1090]), .rdlo_out(a2_wr[1602]));
			radix2 #(.width(width)) rd_st1_1091  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1091]), .rdlo_in(a1_wr[1603]),  .coef_in(coef[134]), .rdup_out(a2_wr[1091]), .rdlo_out(a2_wr[1603]));
			radix2 #(.width(width)) rd_st1_1092  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1092]), .rdlo_in(a1_wr[1604]),  .coef_in(coef[136]), .rdup_out(a2_wr[1092]), .rdlo_out(a2_wr[1604]));
			radix2 #(.width(width)) rd_st1_1093  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1093]), .rdlo_in(a1_wr[1605]),  .coef_in(coef[138]), .rdup_out(a2_wr[1093]), .rdlo_out(a2_wr[1605]));
			radix2 #(.width(width)) rd_st1_1094  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1094]), .rdlo_in(a1_wr[1606]),  .coef_in(coef[140]), .rdup_out(a2_wr[1094]), .rdlo_out(a2_wr[1606]));
			radix2 #(.width(width)) rd_st1_1095  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1095]), .rdlo_in(a1_wr[1607]),  .coef_in(coef[142]), .rdup_out(a2_wr[1095]), .rdlo_out(a2_wr[1607]));
			radix2 #(.width(width)) rd_st1_1096  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1096]), .rdlo_in(a1_wr[1608]),  .coef_in(coef[144]), .rdup_out(a2_wr[1096]), .rdlo_out(a2_wr[1608]));
			radix2 #(.width(width)) rd_st1_1097  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1097]), .rdlo_in(a1_wr[1609]),  .coef_in(coef[146]), .rdup_out(a2_wr[1097]), .rdlo_out(a2_wr[1609]));
			radix2 #(.width(width)) rd_st1_1098  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1098]), .rdlo_in(a1_wr[1610]),  .coef_in(coef[148]), .rdup_out(a2_wr[1098]), .rdlo_out(a2_wr[1610]));
			radix2 #(.width(width)) rd_st1_1099  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1099]), .rdlo_in(a1_wr[1611]),  .coef_in(coef[150]), .rdup_out(a2_wr[1099]), .rdlo_out(a2_wr[1611]));
			radix2 #(.width(width)) rd_st1_1100  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1100]), .rdlo_in(a1_wr[1612]),  .coef_in(coef[152]), .rdup_out(a2_wr[1100]), .rdlo_out(a2_wr[1612]));
			radix2 #(.width(width)) rd_st1_1101  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1101]), .rdlo_in(a1_wr[1613]),  .coef_in(coef[154]), .rdup_out(a2_wr[1101]), .rdlo_out(a2_wr[1613]));
			radix2 #(.width(width)) rd_st1_1102  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1102]), .rdlo_in(a1_wr[1614]),  .coef_in(coef[156]), .rdup_out(a2_wr[1102]), .rdlo_out(a2_wr[1614]));
			radix2 #(.width(width)) rd_st1_1103  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1103]), .rdlo_in(a1_wr[1615]),  .coef_in(coef[158]), .rdup_out(a2_wr[1103]), .rdlo_out(a2_wr[1615]));
			radix2 #(.width(width)) rd_st1_1104  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1104]), .rdlo_in(a1_wr[1616]),  .coef_in(coef[160]), .rdup_out(a2_wr[1104]), .rdlo_out(a2_wr[1616]));
			radix2 #(.width(width)) rd_st1_1105  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1105]), .rdlo_in(a1_wr[1617]),  .coef_in(coef[162]), .rdup_out(a2_wr[1105]), .rdlo_out(a2_wr[1617]));
			radix2 #(.width(width)) rd_st1_1106  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1106]), .rdlo_in(a1_wr[1618]),  .coef_in(coef[164]), .rdup_out(a2_wr[1106]), .rdlo_out(a2_wr[1618]));
			radix2 #(.width(width)) rd_st1_1107  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1107]), .rdlo_in(a1_wr[1619]),  .coef_in(coef[166]), .rdup_out(a2_wr[1107]), .rdlo_out(a2_wr[1619]));
			radix2 #(.width(width)) rd_st1_1108  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1108]), .rdlo_in(a1_wr[1620]),  .coef_in(coef[168]), .rdup_out(a2_wr[1108]), .rdlo_out(a2_wr[1620]));
			radix2 #(.width(width)) rd_st1_1109  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1109]), .rdlo_in(a1_wr[1621]),  .coef_in(coef[170]), .rdup_out(a2_wr[1109]), .rdlo_out(a2_wr[1621]));
			radix2 #(.width(width)) rd_st1_1110  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1110]), .rdlo_in(a1_wr[1622]),  .coef_in(coef[172]), .rdup_out(a2_wr[1110]), .rdlo_out(a2_wr[1622]));
			radix2 #(.width(width)) rd_st1_1111  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1111]), .rdlo_in(a1_wr[1623]),  .coef_in(coef[174]), .rdup_out(a2_wr[1111]), .rdlo_out(a2_wr[1623]));
			radix2 #(.width(width)) rd_st1_1112  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1112]), .rdlo_in(a1_wr[1624]),  .coef_in(coef[176]), .rdup_out(a2_wr[1112]), .rdlo_out(a2_wr[1624]));
			radix2 #(.width(width)) rd_st1_1113  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1113]), .rdlo_in(a1_wr[1625]),  .coef_in(coef[178]), .rdup_out(a2_wr[1113]), .rdlo_out(a2_wr[1625]));
			radix2 #(.width(width)) rd_st1_1114  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1114]), .rdlo_in(a1_wr[1626]),  .coef_in(coef[180]), .rdup_out(a2_wr[1114]), .rdlo_out(a2_wr[1626]));
			radix2 #(.width(width)) rd_st1_1115  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1115]), .rdlo_in(a1_wr[1627]),  .coef_in(coef[182]), .rdup_out(a2_wr[1115]), .rdlo_out(a2_wr[1627]));
			radix2 #(.width(width)) rd_st1_1116  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1116]), .rdlo_in(a1_wr[1628]),  .coef_in(coef[184]), .rdup_out(a2_wr[1116]), .rdlo_out(a2_wr[1628]));
			radix2 #(.width(width)) rd_st1_1117  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1117]), .rdlo_in(a1_wr[1629]),  .coef_in(coef[186]), .rdup_out(a2_wr[1117]), .rdlo_out(a2_wr[1629]));
			radix2 #(.width(width)) rd_st1_1118  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1118]), .rdlo_in(a1_wr[1630]),  .coef_in(coef[188]), .rdup_out(a2_wr[1118]), .rdlo_out(a2_wr[1630]));
			radix2 #(.width(width)) rd_st1_1119  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1119]), .rdlo_in(a1_wr[1631]),  .coef_in(coef[190]), .rdup_out(a2_wr[1119]), .rdlo_out(a2_wr[1631]));
			radix2 #(.width(width)) rd_st1_1120  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1120]), .rdlo_in(a1_wr[1632]),  .coef_in(coef[192]), .rdup_out(a2_wr[1120]), .rdlo_out(a2_wr[1632]));
			radix2 #(.width(width)) rd_st1_1121  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1121]), .rdlo_in(a1_wr[1633]),  .coef_in(coef[194]), .rdup_out(a2_wr[1121]), .rdlo_out(a2_wr[1633]));
			radix2 #(.width(width)) rd_st1_1122  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1122]), .rdlo_in(a1_wr[1634]),  .coef_in(coef[196]), .rdup_out(a2_wr[1122]), .rdlo_out(a2_wr[1634]));
			radix2 #(.width(width)) rd_st1_1123  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1123]), .rdlo_in(a1_wr[1635]),  .coef_in(coef[198]), .rdup_out(a2_wr[1123]), .rdlo_out(a2_wr[1635]));
			radix2 #(.width(width)) rd_st1_1124  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1124]), .rdlo_in(a1_wr[1636]),  .coef_in(coef[200]), .rdup_out(a2_wr[1124]), .rdlo_out(a2_wr[1636]));
			radix2 #(.width(width)) rd_st1_1125  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1125]), .rdlo_in(a1_wr[1637]),  .coef_in(coef[202]), .rdup_out(a2_wr[1125]), .rdlo_out(a2_wr[1637]));
			radix2 #(.width(width)) rd_st1_1126  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1126]), .rdlo_in(a1_wr[1638]),  .coef_in(coef[204]), .rdup_out(a2_wr[1126]), .rdlo_out(a2_wr[1638]));
			radix2 #(.width(width)) rd_st1_1127  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1127]), .rdlo_in(a1_wr[1639]),  .coef_in(coef[206]), .rdup_out(a2_wr[1127]), .rdlo_out(a2_wr[1639]));
			radix2 #(.width(width)) rd_st1_1128  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1128]), .rdlo_in(a1_wr[1640]),  .coef_in(coef[208]), .rdup_out(a2_wr[1128]), .rdlo_out(a2_wr[1640]));
			radix2 #(.width(width)) rd_st1_1129  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1129]), .rdlo_in(a1_wr[1641]),  .coef_in(coef[210]), .rdup_out(a2_wr[1129]), .rdlo_out(a2_wr[1641]));
			radix2 #(.width(width)) rd_st1_1130  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1130]), .rdlo_in(a1_wr[1642]),  .coef_in(coef[212]), .rdup_out(a2_wr[1130]), .rdlo_out(a2_wr[1642]));
			radix2 #(.width(width)) rd_st1_1131  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1131]), .rdlo_in(a1_wr[1643]),  .coef_in(coef[214]), .rdup_out(a2_wr[1131]), .rdlo_out(a2_wr[1643]));
			radix2 #(.width(width)) rd_st1_1132  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1132]), .rdlo_in(a1_wr[1644]),  .coef_in(coef[216]), .rdup_out(a2_wr[1132]), .rdlo_out(a2_wr[1644]));
			radix2 #(.width(width)) rd_st1_1133  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1133]), .rdlo_in(a1_wr[1645]),  .coef_in(coef[218]), .rdup_out(a2_wr[1133]), .rdlo_out(a2_wr[1645]));
			radix2 #(.width(width)) rd_st1_1134  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1134]), .rdlo_in(a1_wr[1646]),  .coef_in(coef[220]), .rdup_out(a2_wr[1134]), .rdlo_out(a2_wr[1646]));
			radix2 #(.width(width)) rd_st1_1135  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1135]), .rdlo_in(a1_wr[1647]),  .coef_in(coef[222]), .rdup_out(a2_wr[1135]), .rdlo_out(a2_wr[1647]));
			radix2 #(.width(width)) rd_st1_1136  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1136]), .rdlo_in(a1_wr[1648]),  .coef_in(coef[224]), .rdup_out(a2_wr[1136]), .rdlo_out(a2_wr[1648]));
			radix2 #(.width(width)) rd_st1_1137  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1137]), .rdlo_in(a1_wr[1649]),  .coef_in(coef[226]), .rdup_out(a2_wr[1137]), .rdlo_out(a2_wr[1649]));
			radix2 #(.width(width)) rd_st1_1138  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1138]), .rdlo_in(a1_wr[1650]),  .coef_in(coef[228]), .rdup_out(a2_wr[1138]), .rdlo_out(a2_wr[1650]));
			radix2 #(.width(width)) rd_st1_1139  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1139]), .rdlo_in(a1_wr[1651]),  .coef_in(coef[230]), .rdup_out(a2_wr[1139]), .rdlo_out(a2_wr[1651]));
			radix2 #(.width(width)) rd_st1_1140  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1140]), .rdlo_in(a1_wr[1652]),  .coef_in(coef[232]), .rdup_out(a2_wr[1140]), .rdlo_out(a2_wr[1652]));
			radix2 #(.width(width)) rd_st1_1141  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1141]), .rdlo_in(a1_wr[1653]),  .coef_in(coef[234]), .rdup_out(a2_wr[1141]), .rdlo_out(a2_wr[1653]));
			radix2 #(.width(width)) rd_st1_1142  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1142]), .rdlo_in(a1_wr[1654]),  .coef_in(coef[236]), .rdup_out(a2_wr[1142]), .rdlo_out(a2_wr[1654]));
			radix2 #(.width(width)) rd_st1_1143  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1143]), .rdlo_in(a1_wr[1655]),  .coef_in(coef[238]), .rdup_out(a2_wr[1143]), .rdlo_out(a2_wr[1655]));
			radix2 #(.width(width)) rd_st1_1144  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1144]), .rdlo_in(a1_wr[1656]),  .coef_in(coef[240]), .rdup_out(a2_wr[1144]), .rdlo_out(a2_wr[1656]));
			radix2 #(.width(width)) rd_st1_1145  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1145]), .rdlo_in(a1_wr[1657]),  .coef_in(coef[242]), .rdup_out(a2_wr[1145]), .rdlo_out(a2_wr[1657]));
			radix2 #(.width(width)) rd_st1_1146  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1146]), .rdlo_in(a1_wr[1658]),  .coef_in(coef[244]), .rdup_out(a2_wr[1146]), .rdlo_out(a2_wr[1658]));
			radix2 #(.width(width)) rd_st1_1147  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1147]), .rdlo_in(a1_wr[1659]),  .coef_in(coef[246]), .rdup_out(a2_wr[1147]), .rdlo_out(a2_wr[1659]));
			radix2 #(.width(width)) rd_st1_1148  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1148]), .rdlo_in(a1_wr[1660]),  .coef_in(coef[248]), .rdup_out(a2_wr[1148]), .rdlo_out(a2_wr[1660]));
			radix2 #(.width(width)) rd_st1_1149  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1149]), .rdlo_in(a1_wr[1661]),  .coef_in(coef[250]), .rdup_out(a2_wr[1149]), .rdlo_out(a2_wr[1661]));
			radix2 #(.width(width)) rd_st1_1150  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1150]), .rdlo_in(a1_wr[1662]),  .coef_in(coef[252]), .rdup_out(a2_wr[1150]), .rdlo_out(a2_wr[1662]));
			radix2 #(.width(width)) rd_st1_1151  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1151]), .rdlo_in(a1_wr[1663]),  .coef_in(coef[254]), .rdup_out(a2_wr[1151]), .rdlo_out(a2_wr[1663]));
			radix2 #(.width(width)) rd_st1_1152  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1152]), .rdlo_in(a1_wr[1664]),  .coef_in(coef[256]), .rdup_out(a2_wr[1152]), .rdlo_out(a2_wr[1664]));
			radix2 #(.width(width)) rd_st1_1153  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1153]), .rdlo_in(a1_wr[1665]),  .coef_in(coef[258]), .rdup_out(a2_wr[1153]), .rdlo_out(a2_wr[1665]));
			radix2 #(.width(width)) rd_st1_1154  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1154]), .rdlo_in(a1_wr[1666]),  .coef_in(coef[260]), .rdup_out(a2_wr[1154]), .rdlo_out(a2_wr[1666]));
			radix2 #(.width(width)) rd_st1_1155  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1155]), .rdlo_in(a1_wr[1667]),  .coef_in(coef[262]), .rdup_out(a2_wr[1155]), .rdlo_out(a2_wr[1667]));
			radix2 #(.width(width)) rd_st1_1156  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1156]), .rdlo_in(a1_wr[1668]),  .coef_in(coef[264]), .rdup_out(a2_wr[1156]), .rdlo_out(a2_wr[1668]));
			radix2 #(.width(width)) rd_st1_1157  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1157]), .rdlo_in(a1_wr[1669]),  .coef_in(coef[266]), .rdup_out(a2_wr[1157]), .rdlo_out(a2_wr[1669]));
			radix2 #(.width(width)) rd_st1_1158  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1158]), .rdlo_in(a1_wr[1670]),  .coef_in(coef[268]), .rdup_out(a2_wr[1158]), .rdlo_out(a2_wr[1670]));
			radix2 #(.width(width)) rd_st1_1159  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1159]), .rdlo_in(a1_wr[1671]),  .coef_in(coef[270]), .rdup_out(a2_wr[1159]), .rdlo_out(a2_wr[1671]));
			radix2 #(.width(width)) rd_st1_1160  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1160]), .rdlo_in(a1_wr[1672]),  .coef_in(coef[272]), .rdup_out(a2_wr[1160]), .rdlo_out(a2_wr[1672]));
			radix2 #(.width(width)) rd_st1_1161  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1161]), .rdlo_in(a1_wr[1673]),  .coef_in(coef[274]), .rdup_out(a2_wr[1161]), .rdlo_out(a2_wr[1673]));
			radix2 #(.width(width)) rd_st1_1162  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1162]), .rdlo_in(a1_wr[1674]),  .coef_in(coef[276]), .rdup_out(a2_wr[1162]), .rdlo_out(a2_wr[1674]));
			radix2 #(.width(width)) rd_st1_1163  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1163]), .rdlo_in(a1_wr[1675]),  .coef_in(coef[278]), .rdup_out(a2_wr[1163]), .rdlo_out(a2_wr[1675]));
			radix2 #(.width(width)) rd_st1_1164  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1164]), .rdlo_in(a1_wr[1676]),  .coef_in(coef[280]), .rdup_out(a2_wr[1164]), .rdlo_out(a2_wr[1676]));
			radix2 #(.width(width)) rd_st1_1165  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1165]), .rdlo_in(a1_wr[1677]),  .coef_in(coef[282]), .rdup_out(a2_wr[1165]), .rdlo_out(a2_wr[1677]));
			radix2 #(.width(width)) rd_st1_1166  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1166]), .rdlo_in(a1_wr[1678]),  .coef_in(coef[284]), .rdup_out(a2_wr[1166]), .rdlo_out(a2_wr[1678]));
			radix2 #(.width(width)) rd_st1_1167  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1167]), .rdlo_in(a1_wr[1679]),  .coef_in(coef[286]), .rdup_out(a2_wr[1167]), .rdlo_out(a2_wr[1679]));
			radix2 #(.width(width)) rd_st1_1168  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1168]), .rdlo_in(a1_wr[1680]),  .coef_in(coef[288]), .rdup_out(a2_wr[1168]), .rdlo_out(a2_wr[1680]));
			radix2 #(.width(width)) rd_st1_1169  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1169]), .rdlo_in(a1_wr[1681]),  .coef_in(coef[290]), .rdup_out(a2_wr[1169]), .rdlo_out(a2_wr[1681]));
			radix2 #(.width(width)) rd_st1_1170  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1170]), .rdlo_in(a1_wr[1682]),  .coef_in(coef[292]), .rdup_out(a2_wr[1170]), .rdlo_out(a2_wr[1682]));
			radix2 #(.width(width)) rd_st1_1171  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1171]), .rdlo_in(a1_wr[1683]),  .coef_in(coef[294]), .rdup_out(a2_wr[1171]), .rdlo_out(a2_wr[1683]));
			radix2 #(.width(width)) rd_st1_1172  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1172]), .rdlo_in(a1_wr[1684]),  .coef_in(coef[296]), .rdup_out(a2_wr[1172]), .rdlo_out(a2_wr[1684]));
			radix2 #(.width(width)) rd_st1_1173  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1173]), .rdlo_in(a1_wr[1685]),  .coef_in(coef[298]), .rdup_out(a2_wr[1173]), .rdlo_out(a2_wr[1685]));
			radix2 #(.width(width)) rd_st1_1174  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1174]), .rdlo_in(a1_wr[1686]),  .coef_in(coef[300]), .rdup_out(a2_wr[1174]), .rdlo_out(a2_wr[1686]));
			radix2 #(.width(width)) rd_st1_1175  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1175]), .rdlo_in(a1_wr[1687]),  .coef_in(coef[302]), .rdup_out(a2_wr[1175]), .rdlo_out(a2_wr[1687]));
			radix2 #(.width(width)) rd_st1_1176  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1176]), .rdlo_in(a1_wr[1688]),  .coef_in(coef[304]), .rdup_out(a2_wr[1176]), .rdlo_out(a2_wr[1688]));
			radix2 #(.width(width)) rd_st1_1177  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1177]), .rdlo_in(a1_wr[1689]),  .coef_in(coef[306]), .rdup_out(a2_wr[1177]), .rdlo_out(a2_wr[1689]));
			radix2 #(.width(width)) rd_st1_1178  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1178]), .rdlo_in(a1_wr[1690]),  .coef_in(coef[308]), .rdup_out(a2_wr[1178]), .rdlo_out(a2_wr[1690]));
			radix2 #(.width(width)) rd_st1_1179  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1179]), .rdlo_in(a1_wr[1691]),  .coef_in(coef[310]), .rdup_out(a2_wr[1179]), .rdlo_out(a2_wr[1691]));
			radix2 #(.width(width)) rd_st1_1180  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1180]), .rdlo_in(a1_wr[1692]),  .coef_in(coef[312]), .rdup_out(a2_wr[1180]), .rdlo_out(a2_wr[1692]));
			radix2 #(.width(width)) rd_st1_1181  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1181]), .rdlo_in(a1_wr[1693]),  .coef_in(coef[314]), .rdup_out(a2_wr[1181]), .rdlo_out(a2_wr[1693]));
			radix2 #(.width(width)) rd_st1_1182  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1182]), .rdlo_in(a1_wr[1694]),  .coef_in(coef[316]), .rdup_out(a2_wr[1182]), .rdlo_out(a2_wr[1694]));
			radix2 #(.width(width)) rd_st1_1183  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1183]), .rdlo_in(a1_wr[1695]),  .coef_in(coef[318]), .rdup_out(a2_wr[1183]), .rdlo_out(a2_wr[1695]));
			radix2 #(.width(width)) rd_st1_1184  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1184]), .rdlo_in(a1_wr[1696]),  .coef_in(coef[320]), .rdup_out(a2_wr[1184]), .rdlo_out(a2_wr[1696]));
			radix2 #(.width(width)) rd_st1_1185  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1185]), .rdlo_in(a1_wr[1697]),  .coef_in(coef[322]), .rdup_out(a2_wr[1185]), .rdlo_out(a2_wr[1697]));
			radix2 #(.width(width)) rd_st1_1186  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1186]), .rdlo_in(a1_wr[1698]),  .coef_in(coef[324]), .rdup_out(a2_wr[1186]), .rdlo_out(a2_wr[1698]));
			radix2 #(.width(width)) rd_st1_1187  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1187]), .rdlo_in(a1_wr[1699]),  .coef_in(coef[326]), .rdup_out(a2_wr[1187]), .rdlo_out(a2_wr[1699]));
			radix2 #(.width(width)) rd_st1_1188  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1188]), .rdlo_in(a1_wr[1700]),  .coef_in(coef[328]), .rdup_out(a2_wr[1188]), .rdlo_out(a2_wr[1700]));
			radix2 #(.width(width)) rd_st1_1189  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1189]), .rdlo_in(a1_wr[1701]),  .coef_in(coef[330]), .rdup_out(a2_wr[1189]), .rdlo_out(a2_wr[1701]));
			radix2 #(.width(width)) rd_st1_1190  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1190]), .rdlo_in(a1_wr[1702]),  .coef_in(coef[332]), .rdup_out(a2_wr[1190]), .rdlo_out(a2_wr[1702]));
			radix2 #(.width(width)) rd_st1_1191  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1191]), .rdlo_in(a1_wr[1703]),  .coef_in(coef[334]), .rdup_out(a2_wr[1191]), .rdlo_out(a2_wr[1703]));
			radix2 #(.width(width)) rd_st1_1192  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1192]), .rdlo_in(a1_wr[1704]),  .coef_in(coef[336]), .rdup_out(a2_wr[1192]), .rdlo_out(a2_wr[1704]));
			radix2 #(.width(width)) rd_st1_1193  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1193]), .rdlo_in(a1_wr[1705]),  .coef_in(coef[338]), .rdup_out(a2_wr[1193]), .rdlo_out(a2_wr[1705]));
			radix2 #(.width(width)) rd_st1_1194  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1194]), .rdlo_in(a1_wr[1706]),  .coef_in(coef[340]), .rdup_out(a2_wr[1194]), .rdlo_out(a2_wr[1706]));
			radix2 #(.width(width)) rd_st1_1195  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1195]), .rdlo_in(a1_wr[1707]),  .coef_in(coef[342]), .rdup_out(a2_wr[1195]), .rdlo_out(a2_wr[1707]));
			radix2 #(.width(width)) rd_st1_1196  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1196]), .rdlo_in(a1_wr[1708]),  .coef_in(coef[344]), .rdup_out(a2_wr[1196]), .rdlo_out(a2_wr[1708]));
			radix2 #(.width(width)) rd_st1_1197  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1197]), .rdlo_in(a1_wr[1709]),  .coef_in(coef[346]), .rdup_out(a2_wr[1197]), .rdlo_out(a2_wr[1709]));
			radix2 #(.width(width)) rd_st1_1198  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1198]), .rdlo_in(a1_wr[1710]),  .coef_in(coef[348]), .rdup_out(a2_wr[1198]), .rdlo_out(a2_wr[1710]));
			radix2 #(.width(width)) rd_st1_1199  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1199]), .rdlo_in(a1_wr[1711]),  .coef_in(coef[350]), .rdup_out(a2_wr[1199]), .rdlo_out(a2_wr[1711]));
			radix2 #(.width(width)) rd_st1_1200  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1200]), .rdlo_in(a1_wr[1712]),  .coef_in(coef[352]), .rdup_out(a2_wr[1200]), .rdlo_out(a2_wr[1712]));
			radix2 #(.width(width)) rd_st1_1201  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1201]), .rdlo_in(a1_wr[1713]),  .coef_in(coef[354]), .rdup_out(a2_wr[1201]), .rdlo_out(a2_wr[1713]));
			radix2 #(.width(width)) rd_st1_1202  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1202]), .rdlo_in(a1_wr[1714]),  .coef_in(coef[356]), .rdup_out(a2_wr[1202]), .rdlo_out(a2_wr[1714]));
			radix2 #(.width(width)) rd_st1_1203  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1203]), .rdlo_in(a1_wr[1715]),  .coef_in(coef[358]), .rdup_out(a2_wr[1203]), .rdlo_out(a2_wr[1715]));
			radix2 #(.width(width)) rd_st1_1204  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1204]), .rdlo_in(a1_wr[1716]),  .coef_in(coef[360]), .rdup_out(a2_wr[1204]), .rdlo_out(a2_wr[1716]));
			radix2 #(.width(width)) rd_st1_1205  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1205]), .rdlo_in(a1_wr[1717]),  .coef_in(coef[362]), .rdup_out(a2_wr[1205]), .rdlo_out(a2_wr[1717]));
			radix2 #(.width(width)) rd_st1_1206  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1206]), .rdlo_in(a1_wr[1718]),  .coef_in(coef[364]), .rdup_out(a2_wr[1206]), .rdlo_out(a2_wr[1718]));
			radix2 #(.width(width)) rd_st1_1207  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1207]), .rdlo_in(a1_wr[1719]),  .coef_in(coef[366]), .rdup_out(a2_wr[1207]), .rdlo_out(a2_wr[1719]));
			radix2 #(.width(width)) rd_st1_1208  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1208]), .rdlo_in(a1_wr[1720]),  .coef_in(coef[368]), .rdup_out(a2_wr[1208]), .rdlo_out(a2_wr[1720]));
			radix2 #(.width(width)) rd_st1_1209  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1209]), .rdlo_in(a1_wr[1721]),  .coef_in(coef[370]), .rdup_out(a2_wr[1209]), .rdlo_out(a2_wr[1721]));
			radix2 #(.width(width)) rd_st1_1210  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1210]), .rdlo_in(a1_wr[1722]),  .coef_in(coef[372]), .rdup_out(a2_wr[1210]), .rdlo_out(a2_wr[1722]));
			radix2 #(.width(width)) rd_st1_1211  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1211]), .rdlo_in(a1_wr[1723]),  .coef_in(coef[374]), .rdup_out(a2_wr[1211]), .rdlo_out(a2_wr[1723]));
			radix2 #(.width(width)) rd_st1_1212  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1212]), .rdlo_in(a1_wr[1724]),  .coef_in(coef[376]), .rdup_out(a2_wr[1212]), .rdlo_out(a2_wr[1724]));
			radix2 #(.width(width)) rd_st1_1213  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1213]), .rdlo_in(a1_wr[1725]),  .coef_in(coef[378]), .rdup_out(a2_wr[1213]), .rdlo_out(a2_wr[1725]));
			radix2 #(.width(width)) rd_st1_1214  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1214]), .rdlo_in(a1_wr[1726]),  .coef_in(coef[380]), .rdup_out(a2_wr[1214]), .rdlo_out(a2_wr[1726]));
			radix2 #(.width(width)) rd_st1_1215  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1215]), .rdlo_in(a1_wr[1727]),  .coef_in(coef[382]), .rdup_out(a2_wr[1215]), .rdlo_out(a2_wr[1727]));
			radix2 #(.width(width)) rd_st1_1216  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1216]), .rdlo_in(a1_wr[1728]),  .coef_in(coef[384]), .rdup_out(a2_wr[1216]), .rdlo_out(a2_wr[1728]));
			radix2 #(.width(width)) rd_st1_1217  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1217]), .rdlo_in(a1_wr[1729]),  .coef_in(coef[386]), .rdup_out(a2_wr[1217]), .rdlo_out(a2_wr[1729]));
			radix2 #(.width(width)) rd_st1_1218  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1218]), .rdlo_in(a1_wr[1730]),  .coef_in(coef[388]), .rdup_out(a2_wr[1218]), .rdlo_out(a2_wr[1730]));
			radix2 #(.width(width)) rd_st1_1219  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1219]), .rdlo_in(a1_wr[1731]),  .coef_in(coef[390]), .rdup_out(a2_wr[1219]), .rdlo_out(a2_wr[1731]));
			radix2 #(.width(width)) rd_st1_1220  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1220]), .rdlo_in(a1_wr[1732]),  .coef_in(coef[392]), .rdup_out(a2_wr[1220]), .rdlo_out(a2_wr[1732]));
			radix2 #(.width(width)) rd_st1_1221  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1221]), .rdlo_in(a1_wr[1733]),  .coef_in(coef[394]), .rdup_out(a2_wr[1221]), .rdlo_out(a2_wr[1733]));
			radix2 #(.width(width)) rd_st1_1222  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1222]), .rdlo_in(a1_wr[1734]),  .coef_in(coef[396]), .rdup_out(a2_wr[1222]), .rdlo_out(a2_wr[1734]));
			radix2 #(.width(width)) rd_st1_1223  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1223]), .rdlo_in(a1_wr[1735]),  .coef_in(coef[398]), .rdup_out(a2_wr[1223]), .rdlo_out(a2_wr[1735]));
			radix2 #(.width(width)) rd_st1_1224  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1224]), .rdlo_in(a1_wr[1736]),  .coef_in(coef[400]), .rdup_out(a2_wr[1224]), .rdlo_out(a2_wr[1736]));
			radix2 #(.width(width)) rd_st1_1225  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1225]), .rdlo_in(a1_wr[1737]),  .coef_in(coef[402]), .rdup_out(a2_wr[1225]), .rdlo_out(a2_wr[1737]));
			radix2 #(.width(width)) rd_st1_1226  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1226]), .rdlo_in(a1_wr[1738]),  .coef_in(coef[404]), .rdup_out(a2_wr[1226]), .rdlo_out(a2_wr[1738]));
			radix2 #(.width(width)) rd_st1_1227  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1227]), .rdlo_in(a1_wr[1739]),  .coef_in(coef[406]), .rdup_out(a2_wr[1227]), .rdlo_out(a2_wr[1739]));
			radix2 #(.width(width)) rd_st1_1228  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1228]), .rdlo_in(a1_wr[1740]),  .coef_in(coef[408]), .rdup_out(a2_wr[1228]), .rdlo_out(a2_wr[1740]));
			radix2 #(.width(width)) rd_st1_1229  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1229]), .rdlo_in(a1_wr[1741]),  .coef_in(coef[410]), .rdup_out(a2_wr[1229]), .rdlo_out(a2_wr[1741]));
			radix2 #(.width(width)) rd_st1_1230  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1230]), .rdlo_in(a1_wr[1742]),  .coef_in(coef[412]), .rdup_out(a2_wr[1230]), .rdlo_out(a2_wr[1742]));
			radix2 #(.width(width)) rd_st1_1231  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1231]), .rdlo_in(a1_wr[1743]),  .coef_in(coef[414]), .rdup_out(a2_wr[1231]), .rdlo_out(a2_wr[1743]));
			radix2 #(.width(width)) rd_st1_1232  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1232]), .rdlo_in(a1_wr[1744]),  .coef_in(coef[416]), .rdup_out(a2_wr[1232]), .rdlo_out(a2_wr[1744]));
			radix2 #(.width(width)) rd_st1_1233  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1233]), .rdlo_in(a1_wr[1745]),  .coef_in(coef[418]), .rdup_out(a2_wr[1233]), .rdlo_out(a2_wr[1745]));
			radix2 #(.width(width)) rd_st1_1234  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1234]), .rdlo_in(a1_wr[1746]),  .coef_in(coef[420]), .rdup_out(a2_wr[1234]), .rdlo_out(a2_wr[1746]));
			radix2 #(.width(width)) rd_st1_1235  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1235]), .rdlo_in(a1_wr[1747]),  .coef_in(coef[422]), .rdup_out(a2_wr[1235]), .rdlo_out(a2_wr[1747]));
			radix2 #(.width(width)) rd_st1_1236  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1236]), .rdlo_in(a1_wr[1748]),  .coef_in(coef[424]), .rdup_out(a2_wr[1236]), .rdlo_out(a2_wr[1748]));
			radix2 #(.width(width)) rd_st1_1237  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1237]), .rdlo_in(a1_wr[1749]),  .coef_in(coef[426]), .rdup_out(a2_wr[1237]), .rdlo_out(a2_wr[1749]));
			radix2 #(.width(width)) rd_st1_1238  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1238]), .rdlo_in(a1_wr[1750]),  .coef_in(coef[428]), .rdup_out(a2_wr[1238]), .rdlo_out(a2_wr[1750]));
			radix2 #(.width(width)) rd_st1_1239  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1239]), .rdlo_in(a1_wr[1751]),  .coef_in(coef[430]), .rdup_out(a2_wr[1239]), .rdlo_out(a2_wr[1751]));
			radix2 #(.width(width)) rd_st1_1240  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1240]), .rdlo_in(a1_wr[1752]),  .coef_in(coef[432]), .rdup_out(a2_wr[1240]), .rdlo_out(a2_wr[1752]));
			radix2 #(.width(width)) rd_st1_1241  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1241]), .rdlo_in(a1_wr[1753]),  .coef_in(coef[434]), .rdup_out(a2_wr[1241]), .rdlo_out(a2_wr[1753]));
			radix2 #(.width(width)) rd_st1_1242  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1242]), .rdlo_in(a1_wr[1754]),  .coef_in(coef[436]), .rdup_out(a2_wr[1242]), .rdlo_out(a2_wr[1754]));
			radix2 #(.width(width)) rd_st1_1243  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1243]), .rdlo_in(a1_wr[1755]),  .coef_in(coef[438]), .rdup_out(a2_wr[1243]), .rdlo_out(a2_wr[1755]));
			radix2 #(.width(width)) rd_st1_1244  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1244]), .rdlo_in(a1_wr[1756]),  .coef_in(coef[440]), .rdup_out(a2_wr[1244]), .rdlo_out(a2_wr[1756]));
			radix2 #(.width(width)) rd_st1_1245  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1245]), .rdlo_in(a1_wr[1757]),  .coef_in(coef[442]), .rdup_out(a2_wr[1245]), .rdlo_out(a2_wr[1757]));
			radix2 #(.width(width)) rd_st1_1246  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1246]), .rdlo_in(a1_wr[1758]),  .coef_in(coef[444]), .rdup_out(a2_wr[1246]), .rdlo_out(a2_wr[1758]));
			radix2 #(.width(width)) rd_st1_1247  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1247]), .rdlo_in(a1_wr[1759]),  .coef_in(coef[446]), .rdup_out(a2_wr[1247]), .rdlo_out(a2_wr[1759]));
			radix2 #(.width(width)) rd_st1_1248  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1248]), .rdlo_in(a1_wr[1760]),  .coef_in(coef[448]), .rdup_out(a2_wr[1248]), .rdlo_out(a2_wr[1760]));
			radix2 #(.width(width)) rd_st1_1249  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1249]), .rdlo_in(a1_wr[1761]),  .coef_in(coef[450]), .rdup_out(a2_wr[1249]), .rdlo_out(a2_wr[1761]));
			radix2 #(.width(width)) rd_st1_1250  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1250]), .rdlo_in(a1_wr[1762]),  .coef_in(coef[452]), .rdup_out(a2_wr[1250]), .rdlo_out(a2_wr[1762]));
			radix2 #(.width(width)) rd_st1_1251  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1251]), .rdlo_in(a1_wr[1763]),  .coef_in(coef[454]), .rdup_out(a2_wr[1251]), .rdlo_out(a2_wr[1763]));
			radix2 #(.width(width)) rd_st1_1252  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1252]), .rdlo_in(a1_wr[1764]),  .coef_in(coef[456]), .rdup_out(a2_wr[1252]), .rdlo_out(a2_wr[1764]));
			radix2 #(.width(width)) rd_st1_1253  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1253]), .rdlo_in(a1_wr[1765]),  .coef_in(coef[458]), .rdup_out(a2_wr[1253]), .rdlo_out(a2_wr[1765]));
			radix2 #(.width(width)) rd_st1_1254  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1254]), .rdlo_in(a1_wr[1766]),  .coef_in(coef[460]), .rdup_out(a2_wr[1254]), .rdlo_out(a2_wr[1766]));
			radix2 #(.width(width)) rd_st1_1255  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1255]), .rdlo_in(a1_wr[1767]),  .coef_in(coef[462]), .rdup_out(a2_wr[1255]), .rdlo_out(a2_wr[1767]));
			radix2 #(.width(width)) rd_st1_1256  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1256]), .rdlo_in(a1_wr[1768]),  .coef_in(coef[464]), .rdup_out(a2_wr[1256]), .rdlo_out(a2_wr[1768]));
			radix2 #(.width(width)) rd_st1_1257  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1257]), .rdlo_in(a1_wr[1769]),  .coef_in(coef[466]), .rdup_out(a2_wr[1257]), .rdlo_out(a2_wr[1769]));
			radix2 #(.width(width)) rd_st1_1258  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1258]), .rdlo_in(a1_wr[1770]),  .coef_in(coef[468]), .rdup_out(a2_wr[1258]), .rdlo_out(a2_wr[1770]));
			radix2 #(.width(width)) rd_st1_1259  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1259]), .rdlo_in(a1_wr[1771]),  .coef_in(coef[470]), .rdup_out(a2_wr[1259]), .rdlo_out(a2_wr[1771]));
			radix2 #(.width(width)) rd_st1_1260  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1260]), .rdlo_in(a1_wr[1772]),  .coef_in(coef[472]), .rdup_out(a2_wr[1260]), .rdlo_out(a2_wr[1772]));
			radix2 #(.width(width)) rd_st1_1261  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1261]), .rdlo_in(a1_wr[1773]),  .coef_in(coef[474]), .rdup_out(a2_wr[1261]), .rdlo_out(a2_wr[1773]));
			radix2 #(.width(width)) rd_st1_1262  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1262]), .rdlo_in(a1_wr[1774]),  .coef_in(coef[476]), .rdup_out(a2_wr[1262]), .rdlo_out(a2_wr[1774]));
			radix2 #(.width(width)) rd_st1_1263  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1263]), .rdlo_in(a1_wr[1775]),  .coef_in(coef[478]), .rdup_out(a2_wr[1263]), .rdlo_out(a2_wr[1775]));
			radix2 #(.width(width)) rd_st1_1264  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1264]), .rdlo_in(a1_wr[1776]),  .coef_in(coef[480]), .rdup_out(a2_wr[1264]), .rdlo_out(a2_wr[1776]));
			radix2 #(.width(width)) rd_st1_1265  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1265]), .rdlo_in(a1_wr[1777]),  .coef_in(coef[482]), .rdup_out(a2_wr[1265]), .rdlo_out(a2_wr[1777]));
			radix2 #(.width(width)) rd_st1_1266  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1266]), .rdlo_in(a1_wr[1778]),  .coef_in(coef[484]), .rdup_out(a2_wr[1266]), .rdlo_out(a2_wr[1778]));
			radix2 #(.width(width)) rd_st1_1267  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1267]), .rdlo_in(a1_wr[1779]),  .coef_in(coef[486]), .rdup_out(a2_wr[1267]), .rdlo_out(a2_wr[1779]));
			radix2 #(.width(width)) rd_st1_1268  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1268]), .rdlo_in(a1_wr[1780]),  .coef_in(coef[488]), .rdup_out(a2_wr[1268]), .rdlo_out(a2_wr[1780]));
			radix2 #(.width(width)) rd_st1_1269  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1269]), .rdlo_in(a1_wr[1781]),  .coef_in(coef[490]), .rdup_out(a2_wr[1269]), .rdlo_out(a2_wr[1781]));
			radix2 #(.width(width)) rd_st1_1270  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1270]), .rdlo_in(a1_wr[1782]),  .coef_in(coef[492]), .rdup_out(a2_wr[1270]), .rdlo_out(a2_wr[1782]));
			radix2 #(.width(width)) rd_st1_1271  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1271]), .rdlo_in(a1_wr[1783]),  .coef_in(coef[494]), .rdup_out(a2_wr[1271]), .rdlo_out(a2_wr[1783]));
			radix2 #(.width(width)) rd_st1_1272  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1272]), .rdlo_in(a1_wr[1784]),  .coef_in(coef[496]), .rdup_out(a2_wr[1272]), .rdlo_out(a2_wr[1784]));
			radix2 #(.width(width)) rd_st1_1273  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1273]), .rdlo_in(a1_wr[1785]),  .coef_in(coef[498]), .rdup_out(a2_wr[1273]), .rdlo_out(a2_wr[1785]));
			radix2 #(.width(width)) rd_st1_1274  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1274]), .rdlo_in(a1_wr[1786]),  .coef_in(coef[500]), .rdup_out(a2_wr[1274]), .rdlo_out(a2_wr[1786]));
			radix2 #(.width(width)) rd_st1_1275  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1275]), .rdlo_in(a1_wr[1787]),  .coef_in(coef[502]), .rdup_out(a2_wr[1275]), .rdlo_out(a2_wr[1787]));
			radix2 #(.width(width)) rd_st1_1276  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1276]), .rdlo_in(a1_wr[1788]),  .coef_in(coef[504]), .rdup_out(a2_wr[1276]), .rdlo_out(a2_wr[1788]));
			radix2 #(.width(width)) rd_st1_1277  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1277]), .rdlo_in(a1_wr[1789]),  .coef_in(coef[506]), .rdup_out(a2_wr[1277]), .rdlo_out(a2_wr[1789]));
			radix2 #(.width(width)) rd_st1_1278  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1278]), .rdlo_in(a1_wr[1790]),  .coef_in(coef[508]), .rdup_out(a2_wr[1278]), .rdlo_out(a2_wr[1790]));
			radix2 #(.width(width)) rd_st1_1279  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1279]), .rdlo_in(a1_wr[1791]),  .coef_in(coef[510]), .rdup_out(a2_wr[1279]), .rdlo_out(a2_wr[1791]));
			radix2 #(.width(width)) rd_st1_1280  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1280]), .rdlo_in(a1_wr[1792]),  .coef_in(coef[512]), .rdup_out(a2_wr[1280]), .rdlo_out(a2_wr[1792]));
			radix2 #(.width(width)) rd_st1_1281  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1281]), .rdlo_in(a1_wr[1793]),  .coef_in(coef[514]), .rdup_out(a2_wr[1281]), .rdlo_out(a2_wr[1793]));
			radix2 #(.width(width)) rd_st1_1282  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1282]), .rdlo_in(a1_wr[1794]),  .coef_in(coef[516]), .rdup_out(a2_wr[1282]), .rdlo_out(a2_wr[1794]));
			radix2 #(.width(width)) rd_st1_1283  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1283]), .rdlo_in(a1_wr[1795]),  .coef_in(coef[518]), .rdup_out(a2_wr[1283]), .rdlo_out(a2_wr[1795]));
			radix2 #(.width(width)) rd_st1_1284  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1284]), .rdlo_in(a1_wr[1796]),  .coef_in(coef[520]), .rdup_out(a2_wr[1284]), .rdlo_out(a2_wr[1796]));
			radix2 #(.width(width)) rd_st1_1285  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1285]), .rdlo_in(a1_wr[1797]),  .coef_in(coef[522]), .rdup_out(a2_wr[1285]), .rdlo_out(a2_wr[1797]));
			radix2 #(.width(width)) rd_st1_1286  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1286]), .rdlo_in(a1_wr[1798]),  .coef_in(coef[524]), .rdup_out(a2_wr[1286]), .rdlo_out(a2_wr[1798]));
			radix2 #(.width(width)) rd_st1_1287  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1287]), .rdlo_in(a1_wr[1799]),  .coef_in(coef[526]), .rdup_out(a2_wr[1287]), .rdlo_out(a2_wr[1799]));
			radix2 #(.width(width)) rd_st1_1288  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1288]), .rdlo_in(a1_wr[1800]),  .coef_in(coef[528]), .rdup_out(a2_wr[1288]), .rdlo_out(a2_wr[1800]));
			radix2 #(.width(width)) rd_st1_1289  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1289]), .rdlo_in(a1_wr[1801]),  .coef_in(coef[530]), .rdup_out(a2_wr[1289]), .rdlo_out(a2_wr[1801]));
			radix2 #(.width(width)) rd_st1_1290  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1290]), .rdlo_in(a1_wr[1802]),  .coef_in(coef[532]), .rdup_out(a2_wr[1290]), .rdlo_out(a2_wr[1802]));
			radix2 #(.width(width)) rd_st1_1291  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1291]), .rdlo_in(a1_wr[1803]),  .coef_in(coef[534]), .rdup_out(a2_wr[1291]), .rdlo_out(a2_wr[1803]));
			radix2 #(.width(width)) rd_st1_1292  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1292]), .rdlo_in(a1_wr[1804]),  .coef_in(coef[536]), .rdup_out(a2_wr[1292]), .rdlo_out(a2_wr[1804]));
			radix2 #(.width(width)) rd_st1_1293  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1293]), .rdlo_in(a1_wr[1805]),  .coef_in(coef[538]), .rdup_out(a2_wr[1293]), .rdlo_out(a2_wr[1805]));
			radix2 #(.width(width)) rd_st1_1294  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1294]), .rdlo_in(a1_wr[1806]),  .coef_in(coef[540]), .rdup_out(a2_wr[1294]), .rdlo_out(a2_wr[1806]));
			radix2 #(.width(width)) rd_st1_1295  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1295]), .rdlo_in(a1_wr[1807]),  .coef_in(coef[542]), .rdup_out(a2_wr[1295]), .rdlo_out(a2_wr[1807]));
			radix2 #(.width(width)) rd_st1_1296  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1296]), .rdlo_in(a1_wr[1808]),  .coef_in(coef[544]), .rdup_out(a2_wr[1296]), .rdlo_out(a2_wr[1808]));
			radix2 #(.width(width)) rd_st1_1297  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1297]), .rdlo_in(a1_wr[1809]),  .coef_in(coef[546]), .rdup_out(a2_wr[1297]), .rdlo_out(a2_wr[1809]));
			radix2 #(.width(width)) rd_st1_1298  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1298]), .rdlo_in(a1_wr[1810]),  .coef_in(coef[548]), .rdup_out(a2_wr[1298]), .rdlo_out(a2_wr[1810]));
			radix2 #(.width(width)) rd_st1_1299  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1299]), .rdlo_in(a1_wr[1811]),  .coef_in(coef[550]), .rdup_out(a2_wr[1299]), .rdlo_out(a2_wr[1811]));
			radix2 #(.width(width)) rd_st1_1300  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1300]), .rdlo_in(a1_wr[1812]),  .coef_in(coef[552]), .rdup_out(a2_wr[1300]), .rdlo_out(a2_wr[1812]));
			radix2 #(.width(width)) rd_st1_1301  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1301]), .rdlo_in(a1_wr[1813]),  .coef_in(coef[554]), .rdup_out(a2_wr[1301]), .rdlo_out(a2_wr[1813]));
			radix2 #(.width(width)) rd_st1_1302  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1302]), .rdlo_in(a1_wr[1814]),  .coef_in(coef[556]), .rdup_out(a2_wr[1302]), .rdlo_out(a2_wr[1814]));
			radix2 #(.width(width)) rd_st1_1303  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1303]), .rdlo_in(a1_wr[1815]),  .coef_in(coef[558]), .rdup_out(a2_wr[1303]), .rdlo_out(a2_wr[1815]));
			radix2 #(.width(width)) rd_st1_1304  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1304]), .rdlo_in(a1_wr[1816]),  .coef_in(coef[560]), .rdup_out(a2_wr[1304]), .rdlo_out(a2_wr[1816]));
			radix2 #(.width(width)) rd_st1_1305  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1305]), .rdlo_in(a1_wr[1817]),  .coef_in(coef[562]), .rdup_out(a2_wr[1305]), .rdlo_out(a2_wr[1817]));
			radix2 #(.width(width)) rd_st1_1306  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1306]), .rdlo_in(a1_wr[1818]),  .coef_in(coef[564]), .rdup_out(a2_wr[1306]), .rdlo_out(a2_wr[1818]));
			radix2 #(.width(width)) rd_st1_1307  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1307]), .rdlo_in(a1_wr[1819]),  .coef_in(coef[566]), .rdup_out(a2_wr[1307]), .rdlo_out(a2_wr[1819]));
			radix2 #(.width(width)) rd_st1_1308  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1308]), .rdlo_in(a1_wr[1820]),  .coef_in(coef[568]), .rdup_out(a2_wr[1308]), .rdlo_out(a2_wr[1820]));
			radix2 #(.width(width)) rd_st1_1309  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1309]), .rdlo_in(a1_wr[1821]),  .coef_in(coef[570]), .rdup_out(a2_wr[1309]), .rdlo_out(a2_wr[1821]));
			radix2 #(.width(width)) rd_st1_1310  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1310]), .rdlo_in(a1_wr[1822]),  .coef_in(coef[572]), .rdup_out(a2_wr[1310]), .rdlo_out(a2_wr[1822]));
			radix2 #(.width(width)) rd_st1_1311  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1311]), .rdlo_in(a1_wr[1823]),  .coef_in(coef[574]), .rdup_out(a2_wr[1311]), .rdlo_out(a2_wr[1823]));
			radix2 #(.width(width)) rd_st1_1312  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1312]), .rdlo_in(a1_wr[1824]),  .coef_in(coef[576]), .rdup_out(a2_wr[1312]), .rdlo_out(a2_wr[1824]));
			radix2 #(.width(width)) rd_st1_1313  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1313]), .rdlo_in(a1_wr[1825]),  .coef_in(coef[578]), .rdup_out(a2_wr[1313]), .rdlo_out(a2_wr[1825]));
			radix2 #(.width(width)) rd_st1_1314  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1314]), .rdlo_in(a1_wr[1826]),  .coef_in(coef[580]), .rdup_out(a2_wr[1314]), .rdlo_out(a2_wr[1826]));
			radix2 #(.width(width)) rd_st1_1315  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1315]), .rdlo_in(a1_wr[1827]),  .coef_in(coef[582]), .rdup_out(a2_wr[1315]), .rdlo_out(a2_wr[1827]));
			radix2 #(.width(width)) rd_st1_1316  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1316]), .rdlo_in(a1_wr[1828]),  .coef_in(coef[584]), .rdup_out(a2_wr[1316]), .rdlo_out(a2_wr[1828]));
			radix2 #(.width(width)) rd_st1_1317  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1317]), .rdlo_in(a1_wr[1829]),  .coef_in(coef[586]), .rdup_out(a2_wr[1317]), .rdlo_out(a2_wr[1829]));
			radix2 #(.width(width)) rd_st1_1318  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1318]), .rdlo_in(a1_wr[1830]),  .coef_in(coef[588]), .rdup_out(a2_wr[1318]), .rdlo_out(a2_wr[1830]));
			radix2 #(.width(width)) rd_st1_1319  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1319]), .rdlo_in(a1_wr[1831]),  .coef_in(coef[590]), .rdup_out(a2_wr[1319]), .rdlo_out(a2_wr[1831]));
			radix2 #(.width(width)) rd_st1_1320  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1320]), .rdlo_in(a1_wr[1832]),  .coef_in(coef[592]), .rdup_out(a2_wr[1320]), .rdlo_out(a2_wr[1832]));
			radix2 #(.width(width)) rd_st1_1321  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1321]), .rdlo_in(a1_wr[1833]),  .coef_in(coef[594]), .rdup_out(a2_wr[1321]), .rdlo_out(a2_wr[1833]));
			radix2 #(.width(width)) rd_st1_1322  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1322]), .rdlo_in(a1_wr[1834]),  .coef_in(coef[596]), .rdup_out(a2_wr[1322]), .rdlo_out(a2_wr[1834]));
			radix2 #(.width(width)) rd_st1_1323  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1323]), .rdlo_in(a1_wr[1835]),  .coef_in(coef[598]), .rdup_out(a2_wr[1323]), .rdlo_out(a2_wr[1835]));
			radix2 #(.width(width)) rd_st1_1324  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1324]), .rdlo_in(a1_wr[1836]),  .coef_in(coef[600]), .rdup_out(a2_wr[1324]), .rdlo_out(a2_wr[1836]));
			radix2 #(.width(width)) rd_st1_1325  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1325]), .rdlo_in(a1_wr[1837]),  .coef_in(coef[602]), .rdup_out(a2_wr[1325]), .rdlo_out(a2_wr[1837]));
			radix2 #(.width(width)) rd_st1_1326  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1326]), .rdlo_in(a1_wr[1838]),  .coef_in(coef[604]), .rdup_out(a2_wr[1326]), .rdlo_out(a2_wr[1838]));
			radix2 #(.width(width)) rd_st1_1327  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1327]), .rdlo_in(a1_wr[1839]),  .coef_in(coef[606]), .rdup_out(a2_wr[1327]), .rdlo_out(a2_wr[1839]));
			radix2 #(.width(width)) rd_st1_1328  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1328]), .rdlo_in(a1_wr[1840]),  .coef_in(coef[608]), .rdup_out(a2_wr[1328]), .rdlo_out(a2_wr[1840]));
			radix2 #(.width(width)) rd_st1_1329  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1329]), .rdlo_in(a1_wr[1841]),  .coef_in(coef[610]), .rdup_out(a2_wr[1329]), .rdlo_out(a2_wr[1841]));
			radix2 #(.width(width)) rd_st1_1330  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1330]), .rdlo_in(a1_wr[1842]),  .coef_in(coef[612]), .rdup_out(a2_wr[1330]), .rdlo_out(a2_wr[1842]));
			radix2 #(.width(width)) rd_st1_1331  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1331]), .rdlo_in(a1_wr[1843]),  .coef_in(coef[614]), .rdup_out(a2_wr[1331]), .rdlo_out(a2_wr[1843]));
			radix2 #(.width(width)) rd_st1_1332  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1332]), .rdlo_in(a1_wr[1844]),  .coef_in(coef[616]), .rdup_out(a2_wr[1332]), .rdlo_out(a2_wr[1844]));
			radix2 #(.width(width)) rd_st1_1333  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1333]), .rdlo_in(a1_wr[1845]),  .coef_in(coef[618]), .rdup_out(a2_wr[1333]), .rdlo_out(a2_wr[1845]));
			radix2 #(.width(width)) rd_st1_1334  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1334]), .rdlo_in(a1_wr[1846]),  .coef_in(coef[620]), .rdup_out(a2_wr[1334]), .rdlo_out(a2_wr[1846]));
			radix2 #(.width(width)) rd_st1_1335  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1335]), .rdlo_in(a1_wr[1847]),  .coef_in(coef[622]), .rdup_out(a2_wr[1335]), .rdlo_out(a2_wr[1847]));
			radix2 #(.width(width)) rd_st1_1336  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1336]), .rdlo_in(a1_wr[1848]),  .coef_in(coef[624]), .rdup_out(a2_wr[1336]), .rdlo_out(a2_wr[1848]));
			radix2 #(.width(width)) rd_st1_1337  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1337]), .rdlo_in(a1_wr[1849]),  .coef_in(coef[626]), .rdup_out(a2_wr[1337]), .rdlo_out(a2_wr[1849]));
			radix2 #(.width(width)) rd_st1_1338  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1338]), .rdlo_in(a1_wr[1850]),  .coef_in(coef[628]), .rdup_out(a2_wr[1338]), .rdlo_out(a2_wr[1850]));
			radix2 #(.width(width)) rd_st1_1339  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1339]), .rdlo_in(a1_wr[1851]),  .coef_in(coef[630]), .rdup_out(a2_wr[1339]), .rdlo_out(a2_wr[1851]));
			radix2 #(.width(width)) rd_st1_1340  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1340]), .rdlo_in(a1_wr[1852]),  .coef_in(coef[632]), .rdup_out(a2_wr[1340]), .rdlo_out(a2_wr[1852]));
			radix2 #(.width(width)) rd_st1_1341  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1341]), .rdlo_in(a1_wr[1853]),  .coef_in(coef[634]), .rdup_out(a2_wr[1341]), .rdlo_out(a2_wr[1853]));
			radix2 #(.width(width)) rd_st1_1342  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1342]), .rdlo_in(a1_wr[1854]),  .coef_in(coef[636]), .rdup_out(a2_wr[1342]), .rdlo_out(a2_wr[1854]));
			radix2 #(.width(width)) rd_st1_1343  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1343]), .rdlo_in(a1_wr[1855]),  .coef_in(coef[638]), .rdup_out(a2_wr[1343]), .rdlo_out(a2_wr[1855]));
			radix2 #(.width(width)) rd_st1_1344  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1344]), .rdlo_in(a1_wr[1856]),  .coef_in(coef[640]), .rdup_out(a2_wr[1344]), .rdlo_out(a2_wr[1856]));
			radix2 #(.width(width)) rd_st1_1345  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1345]), .rdlo_in(a1_wr[1857]),  .coef_in(coef[642]), .rdup_out(a2_wr[1345]), .rdlo_out(a2_wr[1857]));
			radix2 #(.width(width)) rd_st1_1346  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1346]), .rdlo_in(a1_wr[1858]),  .coef_in(coef[644]), .rdup_out(a2_wr[1346]), .rdlo_out(a2_wr[1858]));
			radix2 #(.width(width)) rd_st1_1347  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1347]), .rdlo_in(a1_wr[1859]),  .coef_in(coef[646]), .rdup_out(a2_wr[1347]), .rdlo_out(a2_wr[1859]));
			radix2 #(.width(width)) rd_st1_1348  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1348]), .rdlo_in(a1_wr[1860]),  .coef_in(coef[648]), .rdup_out(a2_wr[1348]), .rdlo_out(a2_wr[1860]));
			radix2 #(.width(width)) rd_st1_1349  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1349]), .rdlo_in(a1_wr[1861]),  .coef_in(coef[650]), .rdup_out(a2_wr[1349]), .rdlo_out(a2_wr[1861]));
			radix2 #(.width(width)) rd_st1_1350  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1350]), .rdlo_in(a1_wr[1862]),  .coef_in(coef[652]), .rdup_out(a2_wr[1350]), .rdlo_out(a2_wr[1862]));
			radix2 #(.width(width)) rd_st1_1351  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1351]), .rdlo_in(a1_wr[1863]),  .coef_in(coef[654]), .rdup_out(a2_wr[1351]), .rdlo_out(a2_wr[1863]));
			radix2 #(.width(width)) rd_st1_1352  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1352]), .rdlo_in(a1_wr[1864]),  .coef_in(coef[656]), .rdup_out(a2_wr[1352]), .rdlo_out(a2_wr[1864]));
			radix2 #(.width(width)) rd_st1_1353  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1353]), .rdlo_in(a1_wr[1865]),  .coef_in(coef[658]), .rdup_out(a2_wr[1353]), .rdlo_out(a2_wr[1865]));
			radix2 #(.width(width)) rd_st1_1354  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1354]), .rdlo_in(a1_wr[1866]),  .coef_in(coef[660]), .rdup_out(a2_wr[1354]), .rdlo_out(a2_wr[1866]));
			radix2 #(.width(width)) rd_st1_1355  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1355]), .rdlo_in(a1_wr[1867]),  .coef_in(coef[662]), .rdup_out(a2_wr[1355]), .rdlo_out(a2_wr[1867]));
			radix2 #(.width(width)) rd_st1_1356  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1356]), .rdlo_in(a1_wr[1868]),  .coef_in(coef[664]), .rdup_out(a2_wr[1356]), .rdlo_out(a2_wr[1868]));
			radix2 #(.width(width)) rd_st1_1357  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1357]), .rdlo_in(a1_wr[1869]),  .coef_in(coef[666]), .rdup_out(a2_wr[1357]), .rdlo_out(a2_wr[1869]));
			radix2 #(.width(width)) rd_st1_1358  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1358]), .rdlo_in(a1_wr[1870]),  .coef_in(coef[668]), .rdup_out(a2_wr[1358]), .rdlo_out(a2_wr[1870]));
			radix2 #(.width(width)) rd_st1_1359  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1359]), .rdlo_in(a1_wr[1871]),  .coef_in(coef[670]), .rdup_out(a2_wr[1359]), .rdlo_out(a2_wr[1871]));
			radix2 #(.width(width)) rd_st1_1360  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1360]), .rdlo_in(a1_wr[1872]),  .coef_in(coef[672]), .rdup_out(a2_wr[1360]), .rdlo_out(a2_wr[1872]));
			radix2 #(.width(width)) rd_st1_1361  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1361]), .rdlo_in(a1_wr[1873]),  .coef_in(coef[674]), .rdup_out(a2_wr[1361]), .rdlo_out(a2_wr[1873]));
			radix2 #(.width(width)) rd_st1_1362  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1362]), .rdlo_in(a1_wr[1874]),  .coef_in(coef[676]), .rdup_out(a2_wr[1362]), .rdlo_out(a2_wr[1874]));
			radix2 #(.width(width)) rd_st1_1363  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1363]), .rdlo_in(a1_wr[1875]),  .coef_in(coef[678]), .rdup_out(a2_wr[1363]), .rdlo_out(a2_wr[1875]));
			radix2 #(.width(width)) rd_st1_1364  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1364]), .rdlo_in(a1_wr[1876]),  .coef_in(coef[680]), .rdup_out(a2_wr[1364]), .rdlo_out(a2_wr[1876]));
			radix2 #(.width(width)) rd_st1_1365  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1365]), .rdlo_in(a1_wr[1877]),  .coef_in(coef[682]), .rdup_out(a2_wr[1365]), .rdlo_out(a2_wr[1877]));
			radix2 #(.width(width)) rd_st1_1366  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1366]), .rdlo_in(a1_wr[1878]),  .coef_in(coef[684]), .rdup_out(a2_wr[1366]), .rdlo_out(a2_wr[1878]));
			radix2 #(.width(width)) rd_st1_1367  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1367]), .rdlo_in(a1_wr[1879]),  .coef_in(coef[686]), .rdup_out(a2_wr[1367]), .rdlo_out(a2_wr[1879]));
			radix2 #(.width(width)) rd_st1_1368  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1368]), .rdlo_in(a1_wr[1880]),  .coef_in(coef[688]), .rdup_out(a2_wr[1368]), .rdlo_out(a2_wr[1880]));
			radix2 #(.width(width)) rd_st1_1369  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1369]), .rdlo_in(a1_wr[1881]),  .coef_in(coef[690]), .rdup_out(a2_wr[1369]), .rdlo_out(a2_wr[1881]));
			radix2 #(.width(width)) rd_st1_1370  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1370]), .rdlo_in(a1_wr[1882]),  .coef_in(coef[692]), .rdup_out(a2_wr[1370]), .rdlo_out(a2_wr[1882]));
			radix2 #(.width(width)) rd_st1_1371  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1371]), .rdlo_in(a1_wr[1883]),  .coef_in(coef[694]), .rdup_out(a2_wr[1371]), .rdlo_out(a2_wr[1883]));
			radix2 #(.width(width)) rd_st1_1372  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1372]), .rdlo_in(a1_wr[1884]),  .coef_in(coef[696]), .rdup_out(a2_wr[1372]), .rdlo_out(a2_wr[1884]));
			radix2 #(.width(width)) rd_st1_1373  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1373]), .rdlo_in(a1_wr[1885]),  .coef_in(coef[698]), .rdup_out(a2_wr[1373]), .rdlo_out(a2_wr[1885]));
			radix2 #(.width(width)) rd_st1_1374  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1374]), .rdlo_in(a1_wr[1886]),  .coef_in(coef[700]), .rdup_out(a2_wr[1374]), .rdlo_out(a2_wr[1886]));
			radix2 #(.width(width)) rd_st1_1375  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1375]), .rdlo_in(a1_wr[1887]),  .coef_in(coef[702]), .rdup_out(a2_wr[1375]), .rdlo_out(a2_wr[1887]));
			radix2 #(.width(width)) rd_st1_1376  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1376]), .rdlo_in(a1_wr[1888]),  .coef_in(coef[704]), .rdup_out(a2_wr[1376]), .rdlo_out(a2_wr[1888]));
			radix2 #(.width(width)) rd_st1_1377  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1377]), .rdlo_in(a1_wr[1889]),  .coef_in(coef[706]), .rdup_out(a2_wr[1377]), .rdlo_out(a2_wr[1889]));
			radix2 #(.width(width)) rd_st1_1378  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1378]), .rdlo_in(a1_wr[1890]),  .coef_in(coef[708]), .rdup_out(a2_wr[1378]), .rdlo_out(a2_wr[1890]));
			radix2 #(.width(width)) rd_st1_1379  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1379]), .rdlo_in(a1_wr[1891]),  .coef_in(coef[710]), .rdup_out(a2_wr[1379]), .rdlo_out(a2_wr[1891]));
			radix2 #(.width(width)) rd_st1_1380  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1380]), .rdlo_in(a1_wr[1892]),  .coef_in(coef[712]), .rdup_out(a2_wr[1380]), .rdlo_out(a2_wr[1892]));
			radix2 #(.width(width)) rd_st1_1381  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1381]), .rdlo_in(a1_wr[1893]),  .coef_in(coef[714]), .rdup_out(a2_wr[1381]), .rdlo_out(a2_wr[1893]));
			radix2 #(.width(width)) rd_st1_1382  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1382]), .rdlo_in(a1_wr[1894]),  .coef_in(coef[716]), .rdup_out(a2_wr[1382]), .rdlo_out(a2_wr[1894]));
			radix2 #(.width(width)) rd_st1_1383  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1383]), .rdlo_in(a1_wr[1895]),  .coef_in(coef[718]), .rdup_out(a2_wr[1383]), .rdlo_out(a2_wr[1895]));
			radix2 #(.width(width)) rd_st1_1384  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1384]), .rdlo_in(a1_wr[1896]),  .coef_in(coef[720]), .rdup_out(a2_wr[1384]), .rdlo_out(a2_wr[1896]));
			radix2 #(.width(width)) rd_st1_1385  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1385]), .rdlo_in(a1_wr[1897]),  .coef_in(coef[722]), .rdup_out(a2_wr[1385]), .rdlo_out(a2_wr[1897]));
			radix2 #(.width(width)) rd_st1_1386  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1386]), .rdlo_in(a1_wr[1898]),  .coef_in(coef[724]), .rdup_out(a2_wr[1386]), .rdlo_out(a2_wr[1898]));
			radix2 #(.width(width)) rd_st1_1387  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1387]), .rdlo_in(a1_wr[1899]),  .coef_in(coef[726]), .rdup_out(a2_wr[1387]), .rdlo_out(a2_wr[1899]));
			radix2 #(.width(width)) rd_st1_1388  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1388]), .rdlo_in(a1_wr[1900]),  .coef_in(coef[728]), .rdup_out(a2_wr[1388]), .rdlo_out(a2_wr[1900]));
			radix2 #(.width(width)) rd_st1_1389  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1389]), .rdlo_in(a1_wr[1901]),  .coef_in(coef[730]), .rdup_out(a2_wr[1389]), .rdlo_out(a2_wr[1901]));
			radix2 #(.width(width)) rd_st1_1390  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1390]), .rdlo_in(a1_wr[1902]),  .coef_in(coef[732]), .rdup_out(a2_wr[1390]), .rdlo_out(a2_wr[1902]));
			radix2 #(.width(width)) rd_st1_1391  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1391]), .rdlo_in(a1_wr[1903]),  .coef_in(coef[734]), .rdup_out(a2_wr[1391]), .rdlo_out(a2_wr[1903]));
			radix2 #(.width(width)) rd_st1_1392  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1392]), .rdlo_in(a1_wr[1904]),  .coef_in(coef[736]), .rdup_out(a2_wr[1392]), .rdlo_out(a2_wr[1904]));
			radix2 #(.width(width)) rd_st1_1393  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1393]), .rdlo_in(a1_wr[1905]),  .coef_in(coef[738]), .rdup_out(a2_wr[1393]), .rdlo_out(a2_wr[1905]));
			radix2 #(.width(width)) rd_st1_1394  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1394]), .rdlo_in(a1_wr[1906]),  .coef_in(coef[740]), .rdup_out(a2_wr[1394]), .rdlo_out(a2_wr[1906]));
			radix2 #(.width(width)) rd_st1_1395  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1395]), .rdlo_in(a1_wr[1907]),  .coef_in(coef[742]), .rdup_out(a2_wr[1395]), .rdlo_out(a2_wr[1907]));
			radix2 #(.width(width)) rd_st1_1396  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1396]), .rdlo_in(a1_wr[1908]),  .coef_in(coef[744]), .rdup_out(a2_wr[1396]), .rdlo_out(a2_wr[1908]));
			radix2 #(.width(width)) rd_st1_1397  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1397]), .rdlo_in(a1_wr[1909]),  .coef_in(coef[746]), .rdup_out(a2_wr[1397]), .rdlo_out(a2_wr[1909]));
			radix2 #(.width(width)) rd_st1_1398  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1398]), .rdlo_in(a1_wr[1910]),  .coef_in(coef[748]), .rdup_out(a2_wr[1398]), .rdlo_out(a2_wr[1910]));
			radix2 #(.width(width)) rd_st1_1399  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1399]), .rdlo_in(a1_wr[1911]),  .coef_in(coef[750]), .rdup_out(a2_wr[1399]), .rdlo_out(a2_wr[1911]));
			radix2 #(.width(width)) rd_st1_1400  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1400]), .rdlo_in(a1_wr[1912]),  .coef_in(coef[752]), .rdup_out(a2_wr[1400]), .rdlo_out(a2_wr[1912]));
			radix2 #(.width(width)) rd_st1_1401  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1401]), .rdlo_in(a1_wr[1913]),  .coef_in(coef[754]), .rdup_out(a2_wr[1401]), .rdlo_out(a2_wr[1913]));
			radix2 #(.width(width)) rd_st1_1402  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1402]), .rdlo_in(a1_wr[1914]),  .coef_in(coef[756]), .rdup_out(a2_wr[1402]), .rdlo_out(a2_wr[1914]));
			radix2 #(.width(width)) rd_st1_1403  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1403]), .rdlo_in(a1_wr[1915]),  .coef_in(coef[758]), .rdup_out(a2_wr[1403]), .rdlo_out(a2_wr[1915]));
			radix2 #(.width(width)) rd_st1_1404  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1404]), .rdlo_in(a1_wr[1916]),  .coef_in(coef[760]), .rdup_out(a2_wr[1404]), .rdlo_out(a2_wr[1916]));
			radix2 #(.width(width)) rd_st1_1405  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1405]), .rdlo_in(a1_wr[1917]),  .coef_in(coef[762]), .rdup_out(a2_wr[1405]), .rdlo_out(a2_wr[1917]));
			radix2 #(.width(width)) rd_st1_1406  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1406]), .rdlo_in(a1_wr[1918]),  .coef_in(coef[764]), .rdup_out(a2_wr[1406]), .rdlo_out(a2_wr[1918]));
			radix2 #(.width(width)) rd_st1_1407  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1407]), .rdlo_in(a1_wr[1919]),  .coef_in(coef[766]), .rdup_out(a2_wr[1407]), .rdlo_out(a2_wr[1919]));
			radix2 #(.width(width)) rd_st1_1408  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1408]), .rdlo_in(a1_wr[1920]),  .coef_in(coef[768]), .rdup_out(a2_wr[1408]), .rdlo_out(a2_wr[1920]));
			radix2 #(.width(width)) rd_st1_1409  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1409]), .rdlo_in(a1_wr[1921]),  .coef_in(coef[770]), .rdup_out(a2_wr[1409]), .rdlo_out(a2_wr[1921]));
			radix2 #(.width(width)) rd_st1_1410  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1410]), .rdlo_in(a1_wr[1922]),  .coef_in(coef[772]), .rdup_out(a2_wr[1410]), .rdlo_out(a2_wr[1922]));
			radix2 #(.width(width)) rd_st1_1411  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1411]), .rdlo_in(a1_wr[1923]),  .coef_in(coef[774]), .rdup_out(a2_wr[1411]), .rdlo_out(a2_wr[1923]));
			radix2 #(.width(width)) rd_st1_1412  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1412]), .rdlo_in(a1_wr[1924]),  .coef_in(coef[776]), .rdup_out(a2_wr[1412]), .rdlo_out(a2_wr[1924]));
			radix2 #(.width(width)) rd_st1_1413  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1413]), .rdlo_in(a1_wr[1925]),  .coef_in(coef[778]), .rdup_out(a2_wr[1413]), .rdlo_out(a2_wr[1925]));
			radix2 #(.width(width)) rd_st1_1414  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1414]), .rdlo_in(a1_wr[1926]),  .coef_in(coef[780]), .rdup_out(a2_wr[1414]), .rdlo_out(a2_wr[1926]));
			radix2 #(.width(width)) rd_st1_1415  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1415]), .rdlo_in(a1_wr[1927]),  .coef_in(coef[782]), .rdup_out(a2_wr[1415]), .rdlo_out(a2_wr[1927]));
			radix2 #(.width(width)) rd_st1_1416  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1416]), .rdlo_in(a1_wr[1928]),  .coef_in(coef[784]), .rdup_out(a2_wr[1416]), .rdlo_out(a2_wr[1928]));
			radix2 #(.width(width)) rd_st1_1417  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1417]), .rdlo_in(a1_wr[1929]),  .coef_in(coef[786]), .rdup_out(a2_wr[1417]), .rdlo_out(a2_wr[1929]));
			radix2 #(.width(width)) rd_st1_1418  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1418]), .rdlo_in(a1_wr[1930]),  .coef_in(coef[788]), .rdup_out(a2_wr[1418]), .rdlo_out(a2_wr[1930]));
			radix2 #(.width(width)) rd_st1_1419  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1419]), .rdlo_in(a1_wr[1931]),  .coef_in(coef[790]), .rdup_out(a2_wr[1419]), .rdlo_out(a2_wr[1931]));
			radix2 #(.width(width)) rd_st1_1420  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1420]), .rdlo_in(a1_wr[1932]),  .coef_in(coef[792]), .rdup_out(a2_wr[1420]), .rdlo_out(a2_wr[1932]));
			radix2 #(.width(width)) rd_st1_1421  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1421]), .rdlo_in(a1_wr[1933]),  .coef_in(coef[794]), .rdup_out(a2_wr[1421]), .rdlo_out(a2_wr[1933]));
			radix2 #(.width(width)) rd_st1_1422  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1422]), .rdlo_in(a1_wr[1934]),  .coef_in(coef[796]), .rdup_out(a2_wr[1422]), .rdlo_out(a2_wr[1934]));
			radix2 #(.width(width)) rd_st1_1423  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1423]), .rdlo_in(a1_wr[1935]),  .coef_in(coef[798]), .rdup_out(a2_wr[1423]), .rdlo_out(a2_wr[1935]));
			radix2 #(.width(width)) rd_st1_1424  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1424]), .rdlo_in(a1_wr[1936]),  .coef_in(coef[800]), .rdup_out(a2_wr[1424]), .rdlo_out(a2_wr[1936]));
			radix2 #(.width(width)) rd_st1_1425  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1425]), .rdlo_in(a1_wr[1937]),  .coef_in(coef[802]), .rdup_out(a2_wr[1425]), .rdlo_out(a2_wr[1937]));
			radix2 #(.width(width)) rd_st1_1426  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1426]), .rdlo_in(a1_wr[1938]),  .coef_in(coef[804]), .rdup_out(a2_wr[1426]), .rdlo_out(a2_wr[1938]));
			radix2 #(.width(width)) rd_st1_1427  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1427]), .rdlo_in(a1_wr[1939]),  .coef_in(coef[806]), .rdup_out(a2_wr[1427]), .rdlo_out(a2_wr[1939]));
			radix2 #(.width(width)) rd_st1_1428  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1428]), .rdlo_in(a1_wr[1940]),  .coef_in(coef[808]), .rdup_out(a2_wr[1428]), .rdlo_out(a2_wr[1940]));
			radix2 #(.width(width)) rd_st1_1429  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1429]), .rdlo_in(a1_wr[1941]),  .coef_in(coef[810]), .rdup_out(a2_wr[1429]), .rdlo_out(a2_wr[1941]));
			radix2 #(.width(width)) rd_st1_1430  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1430]), .rdlo_in(a1_wr[1942]),  .coef_in(coef[812]), .rdup_out(a2_wr[1430]), .rdlo_out(a2_wr[1942]));
			radix2 #(.width(width)) rd_st1_1431  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1431]), .rdlo_in(a1_wr[1943]),  .coef_in(coef[814]), .rdup_out(a2_wr[1431]), .rdlo_out(a2_wr[1943]));
			radix2 #(.width(width)) rd_st1_1432  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1432]), .rdlo_in(a1_wr[1944]),  .coef_in(coef[816]), .rdup_out(a2_wr[1432]), .rdlo_out(a2_wr[1944]));
			radix2 #(.width(width)) rd_st1_1433  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1433]), .rdlo_in(a1_wr[1945]),  .coef_in(coef[818]), .rdup_out(a2_wr[1433]), .rdlo_out(a2_wr[1945]));
			radix2 #(.width(width)) rd_st1_1434  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1434]), .rdlo_in(a1_wr[1946]),  .coef_in(coef[820]), .rdup_out(a2_wr[1434]), .rdlo_out(a2_wr[1946]));
			radix2 #(.width(width)) rd_st1_1435  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1435]), .rdlo_in(a1_wr[1947]),  .coef_in(coef[822]), .rdup_out(a2_wr[1435]), .rdlo_out(a2_wr[1947]));
			radix2 #(.width(width)) rd_st1_1436  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1436]), .rdlo_in(a1_wr[1948]),  .coef_in(coef[824]), .rdup_out(a2_wr[1436]), .rdlo_out(a2_wr[1948]));
			radix2 #(.width(width)) rd_st1_1437  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1437]), .rdlo_in(a1_wr[1949]),  .coef_in(coef[826]), .rdup_out(a2_wr[1437]), .rdlo_out(a2_wr[1949]));
			radix2 #(.width(width)) rd_st1_1438  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1438]), .rdlo_in(a1_wr[1950]),  .coef_in(coef[828]), .rdup_out(a2_wr[1438]), .rdlo_out(a2_wr[1950]));
			radix2 #(.width(width)) rd_st1_1439  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1439]), .rdlo_in(a1_wr[1951]),  .coef_in(coef[830]), .rdup_out(a2_wr[1439]), .rdlo_out(a2_wr[1951]));
			radix2 #(.width(width)) rd_st1_1440  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1440]), .rdlo_in(a1_wr[1952]),  .coef_in(coef[832]), .rdup_out(a2_wr[1440]), .rdlo_out(a2_wr[1952]));
			radix2 #(.width(width)) rd_st1_1441  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1441]), .rdlo_in(a1_wr[1953]),  .coef_in(coef[834]), .rdup_out(a2_wr[1441]), .rdlo_out(a2_wr[1953]));
			radix2 #(.width(width)) rd_st1_1442  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1442]), .rdlo_in(a1_wr[1954]),  .coef_in(coef[836]), .rdup_out(a2_wr[1442]), .rdlo_out(a2_wr[1954]));
			radix2 #(.width(width)) rd_st1_1443  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1443]), .rdlo_in(a1_wr[1955]),  .coef_in(coef[838]), .rdup_out(a2_wr[1443]), .rdlo_out(a2_wr[1955]));
			radix2 #(.width(width)) rd_st1_1444  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1444]), .rdlo_in(a1_wr[1956]),  .coef_in(coef[840]), .rdup_out(a2_wr[1444]), .rdlo_out(a2_wr[1956]));
			radix2 #(.width(width)) rd_st1_1445  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1445]), .rdlo_in(a1_wr[1957]),  .coef_in(coef[842]), .rdup_out(a2_wr[1445]), .rdlo_out(a2_wr[1957]));
			radix2 #(.width(width)) rd_st1_1446  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1446]), .rdlo_in(a1_wr[1958]),  .coef_in(coef[844]), .rdup_out(a2_wr[1446]), .rdlo_out(a2_wr[1958]));
			radix2 #(.width(width)) rd_st1_1447  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1447]), .rdlo_in(a1_wr[1959]),  .coef_in(coef[846]), .rdup_out(a2_wr[1447]), .rdlo_out(a2_wr[1959]));
			radix2 #(.width(width)) rd_st1_1448  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1448]), .rdlo_in(a1_wr[1960]),  .coef_in(coef[848]), .rdup_out(a2_wr[1448]), .rdlo_out(a2_wr[1960]));
			radix2 #(.width(width)) rd_st1_1449  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1449]), .rdlo_in(a1_wr[1961]),  .coef_in(coef[850]), .rdup_out(a2_wr[1449]), .rdlo_out(a2_wr[1961]));
			radix2 #(.width(width)) rd_st1_1450  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1450]), .rdlo_in(a1_wr[1962]),  .coef_in(coef[852]), .rdup_out(a2_wr[1450]), .rdlo_out(a2_wr[1962]));
			radix2 #(.width(width)) rd_st1_1451  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1451]), .rdlo_in(a1_wr[1963]),  .coef_in(coef[854]), .rdup_out(a2_wr[1451]), .rdlo_out(a2_wr[1963]));
			radix2 #(.width(width)) rd_st1_1452  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1452]), .rdlo_in(a1_wr[1964]),  .coef_in(coef[856]), .rdup_out(a2_wr[1452]), .rdlo_out(a2_wr[1964]));
			radix2 #(.width(width)) rd_st1_1453  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1453]), .rdlo_in(a1_wr[1965]),  .coef_in(coef[858]), .rdup_out(a2_wr[1453]), .rdlo_out(a2_wr[1965]));
			radix2 #(.width(width)) rd_st1_1454  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1454]), .rdlo_in(a1_wr[1966]),  .coef_in(coef[860]), .rdup_out(a2_wr[1454]), .rdlo_out(a2_wr[1966]));
			radix2 #(.width(width)) rd_st1_1455  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1455]), .rdlo_in(a1_wr[1967]),  .coef_in(coef[862]), .rdup_out(a2_wr[1455]), .rdlo_out(a2_wr[1967]));
			radix2 #(.width(width)) rd_st1_1456  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1456]), .rdlo_in(a1_wr[1968]),  .coef_in(coef[864]), .rdup_out(a2_wr[1456]), .rdlo_out(a2_wr[1968]));
			radix2 #(.width(width)) rd_st1_1457  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1457]), .rdlo_in(a1_wr[1969]),  .coef_in(coef[866]), .rdup_out(a2_wr[1457]), .rdlo_out(a2_wr[1969]));
			radix2 #(.width(width)) rd_st1_1458  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1458]), .rdlo_in(a1_wr[1970]),  .coef_in(coef[868]), .rdup_out(a2_wr[1458]), .rdlo_out(a2_wr[1970]));
			radix2 #(.width(width)) rd_st1_1459  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1459]), .rdlo_in(a1_wr[1971]),  .coef_in(coef[870]), .rdup_out(a2_wr[1459]), .rdlo_out(a2_wr[1971]));
			radix2 #(.width(width)) rd_st1_1460  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1460]), .rdlo_in(a1_wr[1972]),  .coef_in(coef[872]), .rdup_out(a2_wr[1460]), .rdlo_out(a2_wr[1972]));
			radix2 #(.width(width)) rd_st1_1461  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1461]), .rdlo_in(a1_wr[1973]),  .coef_in(coef[874]), .rdup_out(a2_wr[1461]), .rdlo_out(a2_wr[1973]));
			radix2 #(.width(width)) rd_st1_1462  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1462]), .rdlo_in(a1_wr[1974]),  .coef_in(coef[876]), .rdup_out(a2_wr[1462]), .rdlo_out(a2_wr[1974]));
			radix2 #(.width(width)) rd_st1_1463  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1463]), .rdlo_in(a1_wr[1975]),  .coef_in(coef[878]), .rdup_out(a2_wr[1463]), .rdlo_out(a2_wr[1975]));
			radix2 #(.width(width)) rd_st1_1464  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1464]), .rdlo_in(a1_wr[1976]),  .coef_in(coef[880]), .rdup_out(a2_wr[1464]), .rdlo_out(a2_wr[1976]));
			radix2 #(.width(width)) rd_st1_1465  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1465]), .rdlo_in(a1_wr[1977]),  .coef_in(coef[882]), .rdup_out(a2_wr[1465]), .rdlo_out(a2_wr[1977]));
			radix2 #(.width(width)) rd_st1_1466  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1466]), .rdlo_in(a1_wr[1978]),  .coef_in(coef[884]), .rdup_out(a2_wr[1466]), .rdlo_out(a2_wr[1978]));
			radix2 #(.width(width)) rd_st1_1467  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1467]), .rdlo_in(a1_wr[1979]),  .coef_in(coef[886]), .rdup_out(a2_wr[1467]), .rdlo_out(a2_wr[1979]));
			radix2 #(.width(width)) rd_st1_1468  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1468]), .rdlo_in(a1_wr[1980]),  .coef_in(coef[888]), .rdup_out(a2_wr[1468]), .rdlo_out(a2_wr[1980]));
			radix2 #(.width(width)) rd_st1_1469  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1469]), .rdlo_in(a1_wr[1981]),  .coef_in(coef[890]), .rdup_out(a2_wr[1469]), .rdlo_out(a2_wr[1981]));
			radix2 #(.width(width)) rd_st1_1470  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1470]), .rdlo_in(a1_wr[1982]),  .coef_in(coef[892]), .rdup_out(a2_wr[1470]), .rdlo_out(a2_wr[1982]));
			radix2 #(.width(width)) rd_st1_1471  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1471]), .rdlo_in(a1_wr[1983]),  .coef_in(coef[894]), .rdup_out(a2_wr[1471]), .rdlo_out(a2_wr[1983]));
			radix2 #(.width(width)) rd_st1_1472  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1472]), .rdlo_in(a1_wr[1984]),  .coef_in(coef[896]), .rdup_out(a2_wr[1472]), .rdlo_out(a2_wr[1984]));
			radix2 #(.width(width)) rd_st1_1473  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1473]), .rdlo_in(a1_wr[1985]),  .coef_in(coef[898]), .rdup_out(a2_wr[1473]), .rdlo_out(a2_wr[1985]));
			radix2 #(.width(width)) rd_st1_1474  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1474]), .rdlo_in(a1_wr[1986]),  .coef_in(coef[900]), .rdup_out(a2_wr[1474]), .rdlo_out(a2_wr[1986]));
			radix2 #(.width(width)) rd_st1_1475  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1475]), .rdlo_in(a1_wr[1987]),  .coef_in(coef[902]), .rdup_out(a2_wr[1475]), .rdlo_out(a2_wr[1987]));
			radix2 #(.width(width)) rd_st1_1476  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1476]), .rdlo_in(a1_wr[1988]),  .coef_in(coef[904]), .rdup_out(a2_wr[1476]), .rdlo_out(a2_wr[1988]));
			radix2 #(.width(width)) rd_st1_1477  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1477]), .rdlo_in(a1_wr[1989]),  .coef_in(coef[906]), .rdup_out(a2_wr[1477]), .rdlo_out(a2_wr[1989]));
			radix2 #(.width(width)) rd_st1_1478  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1478]), .rdlo_in(a1_wr[1990]),  .coef_in(coef[908]), .rdup_out(a2_wr[1478]), .rdlo_out(a2_wr[1990]));
			radix2 #(.width(width)) rd_st1_1479  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1479]), .rdlo_in(a1_wr[1991]),  .coef_in(coef[910]), .rdup_out(a2_wr[1479]), .rdlo_out(a2_wr[1991]));
			radix2 #(.width(width)) rd_st1_1480  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1480]), .rdlo_in(a1_wr[1992]),  .coef_in(coef[912]), .rdup_out(a2_wr[1480]), .rdlo_out(a2_wr[1992]));
			radix2 #(.width(width)) rd_st1_1481  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1481]), .rdlo_in(a1_wr[1993]),  .coef_in(coef[914]), .rdup_out(a2_wr[1481]), .rdlo_out(a2_wr[1993]));
			radix2 #(.width(width)) rd_st1_1482  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1482]), .rdlo_in(a1_wr[1994]),  .coef_in(coef[916]), .rdup_out(a2_wr[1482]), .rdlo_out(a2_wr[1994]));
			radix2 #(.width(width)) rd_st1_1483  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1483]), .rdlo_in(a1_wr[1995]),  .coef_in(coef[918]), .rdup_out(a2_wr[1483]), .rdlo_out(a2_wr[1995]));
			radix2 #(.width(width)) rd_st1_1484  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1484]), .rdlo_in(a1_wr[1996]),  .coef_in(coef[920]), .rdup_out(a2_wr[1484]), .rdlo_out(a2_wr[1996]));
			radix2 #(.width(width)) rd_st1_1485  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1485]), .rdlo_in(a1_wr[1997]),  .coef_in(coef[922]), .rdup_out(a2_wr[1485]), .rdlo_out(a2_wr[1997]));
			radix2 #(.width(width)) rd_st1_1486  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1486]), .rdlo_in(a1_wr[1998]),  .coef_in(coef[924]), .rdup_out(a2_wr[1486]), .rdlo_out(a2_wr[1998]));
			radix2 #(.width(width)) rd_st1_1487  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1487]), .rdlo_in(a1_wr[1999]),  .coef_in(coef[926]), .rdup_out(a2_wr[1487]), .rdlo_out(a2_wr[1999]));
			radix2 #(.width(width)) rd_st1_1488  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1488]), .rdlo_in(a1_wr[2000]),  .coef_in(coef[928]), .rdup_out(a2_wr[1488]), .rdlo_out(a2_wr[2000]));
			radix2 #(.width(width)) rd_st1_1489  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1489]), .rdlo_in(a1_wr[2001]),  .coef_in(coef[930]), .rdup_out(a2_wr[1489]), .rdlo_out(a2_wr[2001]));
			radix2 #(.width(width)) rd_st1_1490  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1490]), .rdlo_in(a1_wr[2002]),  .coef_in(coef[932]), .rdup_out(a2_wr[1490]), .rdlo_out(a2_wr[2002]));
			radix2 #(.width(width)) rd_st1_1491  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1491]), .rdlo_in(a1_wr[2003]),  .coef_in(coef[934]), .rdup_out(a2_wr[1491]), .rdlo_out(a2_wr[2003]));
			radix2 #(.width(width)) rd_st1_1492  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1492]), .rdlo_in(a1_wr[2004]),  .coef_in(coef[936]), .rdup_out(a2_wr[1492]), .rdlo_out(a2_wr[2004]));
			radix2 #(.width(width)) rd_st1_1493  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1493]), .rdlo_in(a1_wr[2005]),  .coef_in(coef[938]), .rdup_out(a2_wr[1493]), .rdlo_out(a2_wr[2005]));
			radix2 #(.width(width)) rd_st1_1494  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1494]), .rdlo_in(a1_wr[2006]),  .coef_in(coef[940]), .rdup_out(a2_wr[1494]), .rdlo_out(a2_wr[2006]));
			radix2 #(.width(width)) rd_st1_1495  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1495]), .rdlo_in(a1_wr[2007]),  .coef_in(coef[942]), .rdup_out(a2_wr[1495]), .rdlo_out(a2_wr[2007]));
			radix2 #(.width(width)) rd_st1_1496  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1496]), .rdlo_in(a1_wr[2008]),  .coef_in(coef[944]), .rdup_out(a2_wr[1496]), .rdlo_out(a2_wr[2008]));
			radix2 #(.width(width)) rd_st1_1497  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1497]), .rdlo_in(a1_wr[2009]),  .coef_in(coef[946]), .rdup_out(a2_wr[1497]), .rdlo_out(a2_wr[2009]));
			radix2 #(.width(width)) rd_st1_1498  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1498]), .rdlo_in(a1_wr[2010]),  .coef_in(coef[948]), .rdup_out(a2_wr[1498]), .rdlo_out(a2_wr[2010]));
			radix2 #(.width(width)) rd_st1_1499  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1499]), .rdlo_in(a1_wr[2011]),  .coef_in(coef[950]), .rdup_out(a2_wr[1499]), .rdlo_out(a2_wr[2011]));
			radix2 #(.width(width)) rd_st1_1500  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1500]), .rdlo_in(a1_wr[2012]),  .coef_in(coef[952]), .rdup_out(a2_wr[1500]), .rdlo_out(a2_wr[2012]));
			radix2 #(.width(width)) rd_st1_1501  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1501]), .rdlo_in(a1_wr[2013]),  .coef_in(coef[954]), .rdup_out(a2_wr[1501]), .rdlo_out(a2_wr[2013]));
			radix2 #(.width(width)) rd_st1_1502  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1502]), .rdlo_in(a1_wr[2014]),  .coef_in(coef[956]), .rdup_out(a2_wr[1502]), .rdlo_out(a2_wr[2014]));
			radix2 #(.width(width)) rd_st1_1503  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1503]), .rdlo_in(a1_wr[2015]),  .coef_in(coef[958]), .rdup_out(a2_wr[1503]), .rdlo_out(a2_wr[2015]));
			radix2 #(.width(width)) rd_st1_1504  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1504]), .rdlo_in(a1_wr[2016]),  .coef_in(coef[960]), .rdup_out(a2_wr[1504]), .rdlo_out(a2_wr[2016]));
			radix2 #(.width(width)) rd_st1_1505  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1505]), .rdlo_in(a1_wr[2017]),  .coef_in(coef[962]), .rdup_out(a2_wr[1505]), .rdlo_out(a2_wr[2017]));
			radix2 #(.width(width)) rd_st1_1506  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1506]), .rdlo_in(a1_wr[2018]),  .coef_in(coef[964]), .rdup_out(a2_wr[1506]), .rdlo_out(a2_wr[2018]));
			radix2 #(.width(width)) rd_st1_1507  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1507]), .rdlo_in(a1_wr[2019]),  .coef_in(coef[966]), .rdup_out(a2_wr[1507]), .rdlo_out(a2_wr[2019]));
			radix2 #(.width(width)) rd_st1_1508  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1508]), .rdlo_in(a1_wr[2020]),  .coef_in(coef[968]), .rdup_out(a2_wr[1508]), .rdlo_out(a2_wr[2020]));
			radix2 #(.width(width)) rd_st1_1509  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1509]), .rdlo_in(a1_wr[2021]),  .coef_in(coef[970]), .rdup_out(a2_wr[1509]), .rdlo_out(a2_wr[2021]));
			radix2 #(.width(width)) rd_st1_1510  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1510]), .rdlo_in(a1_wr[2022]),  .coef_in(coef[972]), .rdup_out(a2_wr[1510]), .rdlo_out(a2_wr[2022]));
			radix2 #(.width(width)) rd_st1_1511  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1511]), .rdlo_in(a1_wr[2023]),  .coef_in(coef[974]), .rdup_out(a2_wr[1511]), .rdlo_out(a2_wr[2023]));
			radix2 #(.width(width)) rd_st1_1512  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1512]), .rdlo_in(a1_wr[2024]),  .coef_in(coef[976]), .rdup_out(a2_wr[1512]), .rdlo_out(a2_wr[2024]));
			radix2 #(.width(width)) rd_st1_1513  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1513]), .rdlo_in(a1_wr[2025]),  .coef_in(coef[978]), .rdup_out(a2_wr[1513]), .rdlo_out(a2_wr[2025]));
			radix2 #(.width(width)) rd_st1_1514  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1514]), .rdlo_in(a1_wr[2026]),  .coef_in(coef[980]), .rdup_out(a2_wr[1514]), .rdlo_out(a2_wr[2026]));
			radix2 #(.width(width)) rd_st1_1515  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1515]), .rdlo_in(a1_wr[2027]),  .coef_in(coef[982]), .rdup_out(a2_wr[1515]), .rdlo_out(a2_wr[2027]));
			radix2 #(.width(width)) rd_st1_1516  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1516]), .rdlo_in(a1_wr[2028]),  .coef_in(coef[984]), .rdup_out(a2_wr[1516]), .rdlo_out(a2_wr[2028]));
			radix2 #(.width(width)) rd_st1_1517  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1517]), .rdlo_in(a1_wr[2029]),  .coef_in(coef[986]), .rdup_out(a2_wr[1517]), .rdlo_out(a2_wr[2029]));
			radix2 #(.width(width)) rd_st1_1518  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1518]), .rdlo_in(a1_wr[2030]),  .coef_in(coef[988]), .rdup_out(a2_wr[1518]), .rdlo_out(a2_wr[2030]));
			radix2 #(.width(width)) rd_st1_1519  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1519]), .rdlo_in(a1_wr[2031]),  .coef_in(coef[990]), .rdup_out(a2_wr[1519]), .rdlo_out(a2_wr[2031]));
			radix2 #(.width(width)) rd_st1_1520  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1520]), .rdlo_in(a1_wr[2032]),  .coef_in(coef[992]), .rdup_out(a2_wr[1520]), .rdlo_out(a2_wr[2032]));
			radix2 #(.width(width)) rd_st1_1521  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1521]), .rdlo_in(a1_wr[2033]),  .coef_in(coef[994]), .rdup_out(a2_wr[1521]), .rdlo_out(a2_wr[2033]));
			radix2 #(.width(width)) rd_st1_1522  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1522]), .rdlo_in(a1_wr[2034]),  .coef_in(coef[996]), .rdup_out(a2_wr[1522]), .rdlo_out(a2_wr[2034]));
			radix2 #(.width(width)) rd_st1_1523  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1523]), .rdlo_in(a1_wr[2035]),  .coef_in(coef[998]), .rdup_out(a2_wr[1523]), .rdlo_out(a2_wr[2035]));
			radix2 #(.width(width)) rd_st1_1524  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1524]), .rdlo_in(a1_wr[2036]),  .coef_in(coef[1000]), .rdup_out(a2_wr[1524]), .rdlo_out(a2_wr[2036]));
			radix2 #(.width(width)) rd_st1_1525  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1525]), .rdlo_in(a1_wr[2037]),  .coef_in(coef[1002]), .rdup_out(a2_wr[1525]), .rdlo_out(a2_wr[2037]));
			radix2 #(.width(width)) rd_st1_1526  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1526]), .rdlo_in(a1_wr[2038]),  .coef_in(coef[1004]), .rdup_out(a2_wr[1526]), .rdlo_out(a2_wr[2038]));
			radix2 #(.width(width)) rd_st1_1527  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1527]), .rdlo_in(a1_wr[2039]),  .coef_in(coef[1006]), .rdup_out(a2_wr[1527]), .rdlo_out(a2_wr[2039]));
			radix2 #(.width(width)) rd_st1_1528  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1528]), .rdlo_in(a1_wr[2040]),  .coef_in(coef[1008]), .rdup_out(a2_wr[1528]), .rdlo_out(a2_wr[2040]));
			radix2 #(.width(width)) rd_st1_1529  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1529]), .rdlo_in(a1_wr[2041]),  .coef_in(coef[1010]), .rdup_out(a2_wr[1529]), .rdlo_out(a2_wr[2041]));
			radix2 #(.width(width)) rd_st1_1530  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1530]), .rdlo_in(a1_wr[2042]),  .coef_in(coef[1012]), .rdup_out(a2_wr[1530]), .rdlo_out(a2_wr[2042]));
			radix2 #(.width(width)) rd_st1_1531  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1531]), .rdlo_in(a1_wr[2043]),  .coef_in(coef[1014]), .rdup_out(a2_wr[1531]), .rdlo_out(a2_wr[2043]));
			radix2 #(.width(width)) rd_st1_1532  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1532]), .rdlo_in(a1_wr[2044]),  .coef_in(coef[1016]), .rdup_out(a2_wr[1532]), .rdlo_out(a2_wr[2044]));
			radix2 #(.width(width)) rd_st1_1533  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1533]), .rdlo_in(a1_wr[2045]),  .coef_in(coef[1018]), .rdup_out(a2_wr[1533]), .rdlo_out(a2_wr[2045]));
			radix2 #(.width(width)) rd_st1_1534  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1534]), .rdlo_in(a1_wr[2046]),  .coef_in(coef[1020]), .rdup_out(a2_wr[1534]), .rdlo_out(a2_wr[2046]));
			radix2 #(.width(width)) rd_st1_1535  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a1_wr[1535]), .rdlo_in(a1_wr[2047]),  .coef_in(coef[1022]), .rdup_out(a2_wr[1535]), .rdlo_out(a2_wr[2047]));

		//--- radix stage 2
			radix2 #(.width(width)) rd_st2_0   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[0]), .rdlo_in(a2_wr[256]),  .coef_in(coef[0]), .rdup_out(a3_wr[0]), .rdlo_out(a3_wr[256]));
			radix2 #(.width(width)) rd_st2_1   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1]), .rdlo_in(a2_wr[257]),  .coef_in(coef[4]), .rdup_out(a3_wr[1]), .rdlo_out(a3_wr[257]));
			radix2 #(.width(width)) rd_st2_2   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[2]), .rdlo_in(a2_wr[258]),  .coef_in(coef[8]), .rdup_out(a3_wr[2]), .rdlo_out(a3_wr[258]));
			radix2 #(.width(width)) rd_st2_3   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[3]), .rdlo_in(a2_wr[259]),  .coef_in(coef[12]), .rdup_out(a3_wr[3]), .rdlo_out(a3_wr[259]));
			radix2 #(.width(width)) rd_st2_4   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[4]), .rdlo_in(a2_wr[260]),  .coef_in(coef[16]), .rdup_out(a3_wr[4]), .rdlo_out(a3_wr[260]));
			radix2 #(.width(width)) rd_st2_5   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[5]), .rdlo_in(a2_wr[261]),  .coef_in(coef[20]), .rdup_out(a3_wr[5]), .rdlo_out(a3_wr[261]));
			radix2 #(.width(width)) rd_st2_6   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[6]), .rdlo_in(a2_wr[262]),  .coef_in(coef[24]), .rdup_out(a3_wr[6]), .rdlo_out(a3_wr[262]));
			radix2 #(.width(width)) rd_st2_7   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[7]), .rdlo_in(a2_wr[263]),  .coef_in(coef[28]), .rdup_out(a3_wr[7]), .rdlo_out(a3_wr[263]));
			radix2 #(.width(width)) rd_st2_8   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[8]), .rdlo_in(a2_wr[264]),  .coef_in(coef[32]), .rdup_out(a3_wr[8]), .rdlo_out(a3_wr[264]));
			radix2 #(.width(width)) rd_st2_9   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[9]), .rdlo_in(a2_wr[265]),  .coef_in(coef[36]), .rdup_out(a3_wr[9]), .rdlo_out(a3_wr[265]));
			radix2 #(.width(width)) rd_st2_10  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[10]), .rdlo_in(a2_wr[266]),  .coef_in(coef[40]), .rdup_out(a3_wr[10]), .rdlo_out(a3_wr[266]));
			radix2 #(.width(width)) rd_st2_11  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[11]), .rdlo_in(a2_wr[267]),  .coef_in(coef[44]), .rdup_out(a3_wr[11]), .rdlo_out(a3_wr[267]));
			radix2 #(.width(width)) rd_st2_12  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[12]), .rdlo_in(a2_wr[268]),  .coef_in(coef[48]), .rdup_out(a3_wr[12]), .rdlo_out(a3_wr[268]));
			radix2 #(.width(width)) rd_st2_13  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[13]), .rdlo_in(a2_wr[269]),  .coef_in(coef[52]), .rdup_out(a3_wr[13]), .rdlo_out(a3_wr[269]));
			radix2 #(.width(width)) rd_st2_14  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[14]), .rdlo_in(a2_wr[270]),  .coef_in(coef[56]), .rdup_out(a3_wr[14]), .rdlo_out(a3_wr[270]));
			radix2 #(.width(width)) rd_st2_15  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[15]), .rdlo_in(a2_wr[271]),  .coef_in(coef[60]), .rdup_out(a3_wr[15]), .rdlo_out(a3_wr[271]));
			radix2 #(.width(width)) rd_st2_16  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[16]), .rdlo_in(a2_wr[272]),  .coef_in(coef[64]), .rdup_out(a3_wr[16]), .rdlo_out(a3_wr[272]));
			radix2 #(.width(width)) rd_st2_17  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[17]), .rdlo_in(a2_wr[273]),  .coef_in(coef[68]), .rdup_out(a3_wr[17]), .rdlo_out(a3_wr[273]));
			radix2 #(.width(width)) rd_st2_18  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[18]), .rdlo_in(a2_wr[274]),  .coef_in(coef[72]), .rdup_out(a3_wr[18]), .rdlo_out(a3_wr[274]));
			radix2 #(.width(width)) rd_st2_19  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[19]), .rdlo_in(a2_wr[275]),  .coef_in(coef[76]), .rdup_out(a3_wr[19]), .rdlo_out(a3_wr[275]));
			radix2 #(.width(width)) rd_st2_20  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[20]), .rdlo_in(a2_wr[276]),  .coef_in(coef[80]), .rdup_out(a3_wr[20]), .rdlo_out(a3_wr[276]));
			radix2 #(.width(width)) rd_st2_21  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[21]), .rdlo_in(a2_wr[277]),  .coef_in(coef[84]), .rdup_out(a3_wr[21]), .rdlo_out(a3_wr[277]));
			radix2 #(.width(width)) rd_st2_22  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[22]), .rdlo_in(a2_wr[278]),  .coef_in(coef[88]), .rdup_out(a3_wr[22]), .rdlo_out(a3_wr[278]));
			radix2 #(.width(width)) rd_st2_23  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[23]), .rdlo_in(a2_wr[279]),  .coef_in(coef[92]), .rdup_out(a3_wr[23]), .rdlo_out(a3_wr[279]));
			radix2 #(.width(width)) rd_st2_24  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[24]), .rdlo_in(a2_wr[280]),  .coef_in(coef[96]), .rdup_out(a3_wr[24]), .rdlo_out(a3_wr[280]));
			radix2 #(.width(width)) rd_st2_25  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[25]), .rdlo_in(a2_wr[281]),  .coef_in(coef[100]), .rdup_out(a3_wr[25]), .rdlo_out(a3_wr[281]));
			radix2 #(.width(width)) rd_st2_26  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[26]), .rdlo_in(a2_wr[282]),  .coef_in(coef[104]), .rdup_out(a3_wr[26]), .rdlo_out(a3_wr[282]));
			radix2 #(.width(width)) rd_st2_27  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[27]), .rdlo_in(a2_wr[283]),  .coef_in(coef[108]), .rdup_out(a3_wr[27]), .rdlo_out(a3_wr[283]));
			radix2 #(.width(width)) rd_st2_28  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[28]), .rdlo_in(a2_wr[284]),  .coef_in(coef[112]), .rdup_out(a3_wr[28]), .rdlo_out(a3_wr[284]));
			radix2 #(.width(width)) rd_st2_29  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[29]), .rdlo_in(a2_wr[285]),  .coef_in(coef[116]), .rdup_out(a3_wr[29]), .rdlo_out(a3_wr[285]));
			radix2 #(.width(width)) rd_st2_30  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[30]), .rdlo_in(a2_wr[286]),  .coef_in(coef[120]), .rdup_out(a3_wr[30]), .rdlo_out(a3_wr[286]));
			radix2 #(.width(width)) rd_st2_31  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[31]), .rdlo_in(a2_wr[287]),  .coef_in(coef[124]), .rdup_out(a3_wr[31]), .rdlo_out(a3_wr[287]));
			radix2 #(.width(width)) rd_st2_32  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[32]), .rdlo_in(a2_wr[288]),  .coef_in(coef[128]), .rdup_out(a3_wr[32]), .rdlo_out(a3_wr[288]));
			radix2 #(.width(width)) rd_st2_33  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[33]), .rdlo_in(a2_wr[289]),  .coef_in(coef[132]), .rdup_out(a3_wr[33]), .rdlo_out(a3_wr[289]));
			radix2 #(.width(width)) rd_st2_34  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[34]), .rdlo_in(a2_wr[290]),  .coef_in(coef[136]), .rdup_out(a3_wr[34]), .rdlo_out(a3_wr[290]));
			radix2 #(.width(width)) rd_st2_35  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[35]), .rdlo_in(a2_wr[291]),  .coef_in(coef[140]), .rdup_out(a3_wr[35]), .rdlo_out(a3_wr[291]));
			radix2 #(.width(width)) rd_st2_36  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[36]), .rdlo_in(a2_wr[292]),  .coef_in(coef[144]), .rdup_out(a3_wr[36]), .rdlo_out(a3_wr[292]));
			radix2 #(.width(width)) rd_st2_37  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[37]), .rdlo_in(a2_wr[293]),  .coef_in(coef[148]), .rdup_out(a3_wr[37]), .rdlo_out(a3_wr[293]));
			radix2 #(.width(width)) rd_st2_38  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[38]), .rdlo_in(a2_wr[294]),  .coef_in(coef[152]), .rdup_out(a3_wr[38]), .rdlo_out(a3_wr[294]));
			radix2 #(.width(width)) rd_st2_39  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[39]), .rdlo_in(a2_wr[295]),  .coef_in(coef[156]), .rdup_out(a3_wr[39]), .rdlo_out(a3_wr[295]));
			radix2 #(.width(width)) rd_st2_40  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[40]), .rdlo_in(a2_wr[296]),  .coef_in(coef[160]), .rdup_out(a3_wr[40]), .rdlo_out(a3_wr[296]));
			radix2 #(.width(width)) rd_st2_41  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[41]), .rdlo_in(a2_wr[297]),  .coef_in(coef[164]), .rdup_out(a3_wr[41]), .rdlo_out(a3_wr[297]));
			radix2 #(.width(width)) rd_st2_42  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[42]), .rdlo_in(a2_wr[298]),  .coef_in(coef[168]), .rdup_out(a3_wr[42]), .rdlo_out(a3_wr[298]));
			radix2 #(.width(width)) rd_st2_43  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[43]), .rdlo_in(a2_wr[299]),  .coef_in(coef[172]), .rdup_out(a3_wr[43]), .rdlo_out(a3_wr[299]));
			radix2 #(.width(width)) rd_st2_44  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[44]), .rdlo_in(a2_wr[300]),  .coef_in(coef[176]), .rdup_out(a3_wr[44]), .rdlo_out(a3_wr[300]));
			radix2 #(.width(width)) rd_st2_45  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[45]), .rdlo_in(a2_wr[301]),  .coef_in(coef[180]), .rdup_out(a3_wr[45]), .rdlo_out(a3_wr[301]));
			radix2 #(.width(width)) rd_st2_46  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[46]), .rdlo_in(a2_wr[302]),  .coef_in(coef[184]), .rdup_out(a3_wr[46]), .rdlo_out(a3_wr[302]));
			radix2 #(.width(width)) rd_st2_47  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[47]), .rdlo_in(a2_wr[303]),  .coef_in(coef[188]), .rdup_out(a3_wr[47]), .rdlo_out(a3_wr[303]));
			radix2 #(.width(width)) rd_st2_48  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[48]), .rdlo_in(a2_wr[304]),  .coef_in(coef[192]), .rdup_out(a3_wr[48]), .rdlo_out(a3_wr[304]));
			radix2 #(.width(width)) rd_st2_49  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[49]), .rdlo_in(a2_wr[305]),  .coef_in(coef[196]), .rdup_out(a3_wr[49]), .rdlo_out(a3_wr[305]));
			radix2 #(.width(width)) rd_st2_50  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[50]), .rdlo_in(a2_wr[306]),  .coef_in(coef[200]), .rdup_out(a3_wr[50]), .rdlo_out(a3_wr[306]));
			radix2 #(.width(width)) rd_st2_51  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[51]), .rdlo_in(a2_wr[307]),  .coef_in(coef[204]), .rdup_out(a3_wr[51]), .rdlo_out(a3_wr[307]));
			radix2 #(.width(width)) rd_st2_52  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[52]), .rdlo_in(a2_wr[308]),  .coef_in(coef[208]), .rdup_out(a3_wr[52]), .rdlo_out(a3_wr[308]));
			radix2 #(.width(width)) rd_st2_53  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[53]), .rdlo_in(a2_wr[309]),  .coef_in(coef[212]), .rdup_out(a3_wr[53]), .rdlo_out(a3_wr[309]));
			radix2 #(.width(width)) rd_st2_54  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[54]), .rdlo_in(a2_wr[310]),  .coef_in(coef[216]), .rdup_out(a3_wr[54]), .rdlo_out(a3_wr[310]));
			radix2 #(.width(width)) rd_st2_55  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[55]), .rdlo_in(a2_wr[311]),  .coef_in(coef[220]), .rdup_out(a3_wr[55]), .rdlo_out(a3_wr[311]));
			radix2 #(.width(width)) rd_st2_56  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[56]), .rdlo_in(a2_wr[312]),  .coef_in(coef[224]), .rdup_out(a3_wr[56]), .rdlo_out(a3_wr[312]));
			radix2 #(.width(width)) rd_st2_57  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[57]), .rdlo_in(a2_wr[313]),  .coef_in(coef[228]), .rdup_out(a3_wr[57]), .rdlo_out(a3_wr[313]));
			radix2 #(.width(width)) rd_st2_58  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[58]), .rdlo_in(a2_wr[314]),  .coef_in(coef[232]), .rdup_out(a3_wr[58]), .rdlo_out(a3_wr[314]));
			radix2 #(.width(width)) rd_st2_59  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[59]), .rdlo_in(a2_wr[315]),  .coef_in(coef[236]), .rdup_out(a3_wr[59]), .rdlo_out(a3_wr[315]));
			radix2 #(.width(width)) rd_st2_60  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[60]), .rdlo_in(a2_wr[316]),  .coef_in(coef[240]), .rdup_out(a3_wr[60]), .rdlo_out(a3_wr[316]));
			radix2 #(.width(width)) rd_st2_61  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[61]), .rdlo_in(a2_wr[317]),  .coef_in(coef[244]), .rdup_out(a3_wr[61]), .rdlo_out(a3_wr[317]));
			radix2 #(.width(width)) rd_st2_62  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[62]), .rdlo_in(a2_wr[318]),  .coef_in(coef[248]), .rdup_out(a3_wr[62]), .rdlo_out(a3_wr[318]));
			radix2 #(.width(width)) rd_st2_63  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[63]), .rdlo_in(a2_wr[319]),  .coef_in(coef[252]), .rdup_out(a3_wr[63]), .rdlo_out(a3_wr[319]));
			radix2 #(.width(width)) rd_st2_64  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[64]), .rdlo_in(a2_wr[320]),  .coef_in(coef[256]), .rdup_out(a3_wr[64]), .rdlo_out(a3_wr[320]));
			radix2 #(.width(width)) rd_st2_65  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[65]), .rdlo_in(a2_wr[321]),  .coef_in(coef[260]), .rdup_out(a3_wr[65]), .rdlo_out(a3_wr[321]));
			radix2 #(.width(width)) rd_st2_66  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[66]), .rdlo_in(a2_wr[322]),  .coef_in(coef[264]), .rdup_out(a3_wr[66]), .rdlo_out(a3_wr[322]));
			radix2 #(.width(width)) rd_st2_67  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[67]), .rdlo_in(a2_wr[323]),  .coef_in(coef[268]), .rdup_out(a3_wr[67]), .rdlo_out(a3_wr[323]));
			radix2 #(.width(width)) rd_st2_68  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[68]), .rdlo_in(a2_wr[324]),  .coef_in(coef[272]), .rdup_out(a3_wr[68]), .rdlo_out(a3_wr[324]));
			radix2 #(.width(width)) rd_st2_69  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[69]), .rdlo_in(a2_wr[325]),  .coef_in(coef[276]), .rdup_out(a3_wr[69]), .rdlo_out(a3_wr[325]));
			radix2 #(.width(width)) rd_st2_70  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[70]), .rdlo_in(a2_wr[326]),  .coef_in(coef[280]), .rdup_out(a3_wr[70]), .rdlo_out(a3_wr[326]));
			radix2 #(.width(width)) rd_st2_71  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[71]), .rdlo_in(a2_wr[327]),  .coef_in(coef[284]), .rdup_out(a3_wr[71]), .rdlo_out(a3_wr[327]));
			radix2 #(.width(width)) rd_st2_72  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[72]), .rdlo_in(a2_wr[328]),  .coef_in(coef[288]), .rdup_out(a3_wr[72]), .rdlo_out(a3_wr[328]));
			radix2 #(.width(width)) rd_st2_73  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[73]), .rdlo_in(a2_wr[329]),  .coef_in(coef[292]), .rdup_out(a3_wr[73]), .rdlo_out(a3_wr[329]));
			radix2 #(.width(width)) rd_st2_74  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[74]), .rdlo_in(a2_wr[330]),  .coef_in(coef[296]), .rdup_out(a3_wr[74]), .rdlo_out(a3_wr[330]));
			radix2 #(.width(width)) rd_st2_75  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[75]), .rdlo_in(a2_wr[331]),  .coef_in(coef[300]), .rdup_out(a3_wr[75]), .rdlo_out(a3_wr[331]));
			radix2 #(.width(width)) rd_st2_76  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[76]), .rdlo_in(a2_wr[332]),  .coef_in(coef[304]), .rdup_out(a3_wr[76]), .rdlo_out(a3_wr[332]));
			radix2 #(.width(width)) rd_st2_77  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[77]), .rdlo_in(a2_wr[333]),  .coef_in(coef[308]), .rdup_out(a3_wr[77]), .rdlo_out(a3_wr[333]));
			radix2 #(.width(width)) rd_st2_78  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[78]), .rdlo_in(a2_wr[334]),  .coef_in(coef[312]), .rdup_out(a3_wr[78]), .rdlo_out(a3_wr[334]));
			radix2 #(.width(width)) rd_st2_79  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[79]), .rdlo_in(a2_wr[335]),  .coef_in(coef[316]), .rdup_out(a3_wr[79]), .rdlo_out(a3_wr[335]));
			radix2 #(.width(width)) rd_st2_80  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[80]), .rdlo_in(a2_wr[336]),  .coef_in(coef[320]), .rdup_out(a3_wr[80]), .rdlo_out(a3_wr[336]));
			radix2 #(.width(width)) rd_st2_81  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[81]), .rdlo_in(a2_wr[337]),  .coef_in(coef[324]), .rdup_out(a3_wr[81]), .rdlo_out(a3_wr[337]));
			radix2 #(.width(width)) rd_st2_82  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[82]), .rdlo_in(a2_wr[338]),  .coef_in(coef[328]), .rdup_out(a3_wr[82]), .rdlo_out(a3_wr[338]));
			radix2 #(.width(width)) rd_st2_83  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[83]), .rdlo_in(a2_wr[339]),  .coef_in(coef[332]), .rdup_out(a3_wr[83]), .rdlo_out(a3_wr[339]));
			radix2 #(.width(width)) rd_st2_84  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[84]), .rdlo_in(a2_wr[340]),  .coef_in(coef[336]), .rdup_out(a3_wr[84]), .rdlo_out(a3_wr[340]));
			radix2 #(.width(width)) rd_st2_85  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[85]), .rdlo_in(a2_wr[341]),  .coef_in(coef[340]), .rdup_out(a3_wr[85]), .rdlo_out(a3_wr[341]));
			radix2 #(.width(width)) rd_st2_86  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[86]), .rdlo_in(a2_wr[342]),  .coef_in(coef[344]), .rdup_out(a3_wr[86]), .rdlo_out(a3_wr[342]));
			radix2 #(.width(width)) rd_st2_87  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[87]), .rdlo_in(a2_wr[343]),  .coef_in(coef[348]), .rdup_out(a3_wr[87]), .rdlo_out(a3_wr[343]));
			radix2 #(.width(width)) rd_st2_88  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[88]), .rdlo_in(a2_wr[344]),  .coef_in(coef[352]), .rdup_out(a3_wr[88]), .rdlo_out(a3_wr[344]));
			radix2 #(.width(width)) rd_st2_89  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[89]), .rdlo_in(a2_wr[345]),  .coef_in(coef[356]), .rdup_out(a3_wr[89]), .rdlo_out(a3_wr[345]));
			radix2 #(.width(width)) rd_st2_90  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[90]), .rdlo_in(a2_wr[346]),  .coef_in(coef[360]), .rdup_out(a3_wr[90]), .rdlo_out(a3_wr[346]));
			radix2 #(.width(width)) rd_st2_91  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[91]), .rdlo_in(a2_wr[347]),  .coef_in(coef[364]), .rdup_out(a3_wr[91]), .rdlo_out(a3_wr[347]));
			radix2 #(.width(width)) rd_st2_92  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[92]), .rdlo_in(a2_wr[348]),  .coef_in(coef[368]), .rdup_out(a3_wr[92]), .rdlo_out(a3_wr[348]));
			radix2 #(.width(width)) rd_st2_93  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[93]), .rdlo_in(a2_wr[349]),  .coef_in(coef[372]), .rdup_out(a3_wr[93]), .rdlo_out(a3_wr[349]));
			radix2 #(.width(width)) rd_st2_94  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[94]), .rdlo_in(a2_wr[350]),  .coef_in(coef[376]), .rdup_out(a3_wr[94]), .rdlo_out(a3_wr[350]));
			radix2 #(.width(width)) rd_st2_95  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[95]), .rdlo_in(a2_wr[351]),  .coef_in(coef[380]), .rdup_out(a3_wr[95]), .rdlo_out(a3_wr[351]));
			radix2 #(.width(width)) rd_st2_96  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[96]), .rdlo_in(a2_wr[352]),  .coef_in(coef[384]), .rdup_out(a3_wr[96]), .rdlo_out(a3_wr[352]));
			radix2 #(.width(width)) rd_st2_97  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[97]), .rdlo_in(a2_wr[353]),  .coef_in(coef[388]), .rdup_out(a3_wr[97]), .rdlo_out(a3_wr[353]));
			radix2 #(.width(width)) rd_st2_98  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[98]), .rdlo_in(a2_wr[354]),  .coef_in(coef[392]), .rdup_out(a3_wr[98]), .rdlo_out(a3_wr[354]));
			radix2 #(.width(width)) rd_st2_99  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[99]), .rdlo_in(a2_wr[355]),  .coef_in(coef[396]), .rdup_out(a3_wr[99]), .rdlo_out(a3_wr[355]));
			radix2 #(.width(width)) rd_st2_100  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[100]), .rdlo_in(a2_wr[356]),  .coef_in(coef[400]), .rdup_out(a3_wr[100]), .rdlo_out(a3_wr[356]));
			radix2 #(.width(width)) rd_st2_101  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[101]), .rdlo_in(a2_wr[357]),  .coef_in(coef[404]), .rdup_out(a3_wr[101]), .rdlo_out(a3_wr[357]));
			radix2 #(.width(width)) rd_st2_102  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[102]), .rdlo_in(a2_wr[358]),  .coef_in(coef[408]), .rdup_out(a3_wr[102]), .rdlo_out(a3_wr[358]));
			radix2 #(.width(width)) rd_st2_103  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[103]), .rdlo_in(a2_wr[359]),  .coef_in(coef[412]), .rdup_out(a3_wr[103]), .rdlo_out(a3_wr[359]));
			radix2 #(.width(width)) rd_st2_104  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[104]), .rdlo_in(a2_wr[360]),  .coef_in(coef[416]), .rdup_out(a3_wr[104]), .rdlo_out(a3_wr[360]));
			radix2 #(.width(width)) rd_st2_105  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[105]), .rdlo_in(a2_wr[361]),  .coef_in(coef[420]), .rdup_out(a3_wr[105]), .rdlo_out(a3_wr[361]));
			radix2 #(.width(width)) rd_st2_106  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[106]), .rdlo_in(a2_wr[362]),  .coef_in(coef[424]), .rdup_out(a3_wr[106]), .rdlo_out(a3_wr[362]));
			radix2 #(.width(width)) rd_st2_107  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[107]), .rdlo_in(a2_wr[363]),  .coef_in(coef[428]), .rdup_out(a3_wr[107]), .rdlo_out(a3_wr[363]));
			radix2 #(.width(width)) rd_st2_108  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[108]), .rdlo_in(a2_wr[364]),  .coef_in(coef[432]), .rdup_out(a3_wr[108]), .rdlo_out(a3_wr[364]));
			radix2 #(.width(width)) rd_st2_109  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[109]), .rdlo_in(a2_wr[365]),  .coef_in(coef[436]), .rdup_out(a3_wr[109]), .rdlo_out(a3_wr[365]));
			radix2 #(.width(width)) rd_st2_110  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[110]), .rdlo_in(a2_wr[366]),  .coef_in(coef[440]), .rdup_out(a3_wr[110]), .rdlo_out(a3_wr[366]));
			radix2 #(.width(width)) rd_st2_111  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[111]), .rdlo_in(a2_wr[367]),  .coef_in(coef[444]), .rdup_out(a3_wr[111]), .rdlo_out(a3_wr[367]));
			radix2 #(.width(width)) rd_st2_112  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[112]), .rdlo_in(a2_wr[368]),  .coef_in(coef[448]), .rdup_out(a3_wr[112]), .rdlo_out(a3_wr[368]));
			radix2 #(.width(width)) rd_st2_113  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[113]), .rdlo_in(a2_wr[369]),  .coef_in(coef[452]), .rdup_out(a3_wr[113]), .rdlo_out(a3_wr[369]));
			radix2 #(.width(width)) rd_st2_114  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[114]), .rdlo_in(a2_wr[370]),  .coef_in(coef[456]), .rdup_out(a3_wr[114]), .rdlo_out(a3_wr[370]));
			radix2 #(.width(width)) rd_st2_115  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[115]), .rdlo_in(a2_wr[371]),  .coef_in(coef[460]), .rdup_out(a3_wr[115]), .rdlo_out(a3_wr[371]));
			radix2 #(.width(width)) rd_st2_116  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[116]), .rdlo_in(a2_wr[372]),  .coef_in(coef[464]), .rdup_out(a3_wr[116]), .rdlo_out(a3_wr[372]));
			radix2 #(.width(width)) rd_st2_117  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[117]), .rdlo_in(a2_wr[373]),  .coef_in(coef[468]), .rdup_out(a3_wr[117]), .rdlo_out(a3_wr[373]));
			radix2 #(.width(width)) rd_st2_118  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[118]), .rdlo_in(a2_wr[374]),  .coef_in(coef[472]), .rdup_out(a3_wr[118]), .rdlo_out(a3_wr[374]));
			radix2 #(.width(width)) rd_st2_119  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[119]), .rdlo_in(a2_wr[375]),  .coef_in(coef[476]), .rdup_out(a3_wr[119]), .rdlo_out(a3_wr[375]));
			radix2 #(.width(width)) rd_st2_120  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[120]), .rdlo_in(a2_wr[376]),  .coef_in(coef[480]), .rdup_out(a3_wr[120]), .rdlo_out(a3_wr[376]));
			radix2 #(.width(width)) rd_st2_121  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[121]), .rdlo_in(a2_wr[377]),  .coef_in(coef[484]), .rdup_out(a3_wr[121]), .rdlo_out(a3_wr[377]));
			radix2 #(.width(width)) rd_st2_122  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[122]), .rdlo_in(a2_wr[378]),  .coef_in(coef[488]), .rdup_out(a3_wr[122]), .rdlo_out(a3_wr[378]));
			radix2 #(.width(width)) rd_st2_123  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[123]), .rdlo_in(a2_wr[379]),  .coef_in(coef[492]), .rdup_out(a3_wr[123]), .rdlo_out(a3_wr[379]));
			radix2 #(.width(width)) rd_st2_124  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[124]), .rdlo_in(a2_wr[380]),  .coef_in(coef[496]), .rdup_out(a3_wr[124]), .rdlo_out(a3_wr[380]));
			radix2 #(.width(width)) rd_st2_125  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[125]), .rdlo_in(a2_wr[381]),  .coef_in(coef[500]), .rdup_out(a3_wr[125]), .rdlo_out(a3_wr[381]));
			radix2 #(.width(width)) rd_st2_126  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[126]), .rdlo_in(a2_wr[382]),  .coef_in(coef[504]), .rdup_out(a3_wr[126]), .rdlo_out(a3_wr[382]));
			radix2 #(.width(width)) rd_st2_127  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[127]), .rdlo_in(a2_wr[383]),  .coef_in(coef[508]), .rdup_out(a3_wr[127]), .rdlo_out(a3_wr[383]));
			radix2 #(.width(width)) rd_st2_128  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[128]), .rdlo_in(a2_wr[384]),  .coef_in(coef[512]), .rdup_out(a3_wr[128]), .rdlo_out(a3_wr[384]));
			radix2 #(.width(width)) rd_st2_129  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[129]), .rdlo_in(a2_wr[385]),  .coef_in(coef[516]), .rdup_out(a3_wr[129]), .rdlo_out(a3_wr[385]));
			radix2 #(.width(width)) rd_st2_130  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[130]), .rdlo_in(a2_wr[386]),  .coef_in(coef[520]), .rdup_out(a3_wr[130]), .rdlo_out(a3_wr[386]));
			radix2 #(.width(width)) rd_st2_131  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[131]), .rdlo_in(a2_wr[387]),  .coef_in(coef[524]), .rdup_out(a3_wr[131]), .rdlo_out(a3_wr[387]));
			radix2 #(.width(width)) rd_st2_132  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[132]), .rdlo_in(a2_wr[388]),  .coef_in(coef[528]), .rdup_out(a3_wr[132]), .rdlo_out(a3_wr[388]));
			radix2 #(.width(width)) rd_st2_133  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[133]), .rdlo_in(a2_wr[389]),  .coef_in(coef[532]), .rdup_out(a3_wr[133]), .rdlo_out(a3_wr[389]));
			radix2 #(.width(width)) rd_st2_134  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[134]), .rdlo_in(a2_wr[390]),  .coef_in(coef[536]), .rdup_out(a3_wr[134]), .rdlo_out(a3_wr[390]));
			radix2 #(.width(width)) rd_st2_135  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[135]), .rdlo_in(a2_wr[391]),  .coef_in(coef[540]), .rdup_out(a3_wr[135]), .rdlo_out(a3_wr[391]));
			radix2 #(.width(width)) rd_st2_136  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[136]), .rdlo_in(a2_wr[392]),  .coef_in(coef[544]), .rdup_out(a3_wr[136]), .rdlo_out(a3_wr[392]));
			radix2 #(.width(width)) rd_st2_137  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[137]), .rdlo_in(a2_wr[393]),  .coef_in(coef[548]), .rdup_out(a3_wr[137]), .rdlo_out(a3_wr[393]));
			radix2 #(.width(width)) rd_st2_138  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[138]), .rdlo_in(a2_wr[394]),  .coef_in(coef[552]), .rdup_out(a3_wr[138]), .rdlo_out(a3_wr[394]));
			radix2 #(.width(width)) rd_st2_139  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[139]), .rdlo_in(a2_wr[395]),  .coef_in(coef[556]), .rdup_out(a3_wr[139]), .rdlo_out(a3_wr[395]));
			radix2 #(.width(width)) rd_st2_140  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[140]), .rdlo_in(a2_wr[396]),  .coef_in(coef[560]), .rdup_out(a3_wr[140]), .rdlo_out(a3_wr[396]));
			radix2 #(.width(width)) rd_st2_141  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[141]), .rdlo_in(a2_wr[397]),  .coef_in(coef[564]), .rdup_out(a3_wr[141]), .rdlo_out(a3_wr[397]));
			radix2 #(.width(width)) rd_st2_142  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[142]), .rdlo_in(a2_wr[398]),  .coef_in(coef[568]), .rdup_out(a3_wr[142]), .rdlo_out(a3_wr[398]));
			radix2 #(.width(width)) rd_st2_143  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[143]), .rdlo_in(a2_wr[399]),  .coef_in(coef[572]), .rdup_out(a3_wr[143]), .rdlo_out(a3_wr[399]));
			radix2 #(.width(width)) rd_st2_144  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[144]), .rdlo_in(a2_wr[400]),  .coef_in(coef[576]), .rdup_out(a3_wr[144]), .rdlo_out(a3_wr[400]));
			radix2 #(.width(width)) rd_st2_145  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[145]), .rdlo_in(a2_wr[401]),  .coef_in(coef[580]), .rdup_out(a3_wr[145]), .rdlo_out(a3_wr[401]));
			radix2 #(.width(width)) rd_st2_146  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[146]), .rdlo_in(a2_wr[402]),  .coef_in(coef[584]), .rdup_out(a3_wr[146]), .rdlo_out(a3_wr[402]));
			radix2 #(.width(width)) rd_st2_147  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[147]), .rdlo_in(a2_wr[403]),  .coef_in(coef[588]), .rdup_out(a3_wr[147]), .rdlo_out(a3_wr[403]));
			radix2 #(.width(width)) rd_st2_148  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[148]), .rdlo_in(a2_wr[404]),  .coef_in(coef[592]), .rdup_out(a3_wr[148]), .rdlo_out(a3_wr[404]));
			radix2 #(.width(width)) rd_st2_149  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[149]), .rdlo_in(a2_wr[405]),  .coef_in(coef[596]), .rdup_out(a3_wr[149]), .rdlo_out(a3_wr[405]));
			radix2 #(.width(width)) rd_st2_150  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[150]), .rdlo_in(a2_wr[406]),  .coef_in(coef[600]), .rdup_out(a3_wr[150]), .rdlo_out(a3_wr[406]));
			radix2 #(.width(width)) rd_st2_151  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[151]), .rdlo_in(a2_wr[407]),  .coef_in(coef[604]), .rdup_out(a3_wr[151]), .rdlo_out(a3_wr[407]));
			radix2 #(.width(width)) rd_st2_152  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[152]), .rdlo_in(a2_wr[408]),  .coef_in(coef[608]), .rdup_out(a3_wr[152]), .rdlo_out(a3_wr[408]));
			radix2 #(.width(width)) rd_st2_153  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[153]), .rdlo_in(a2_wr[409]),  .coef_in(coef[612]), .rdup_out(a3_wr[153]), .rdlo_out(a3_wr[409]));
			radix2 #(.width(width)) rd_st2_154  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[154]), .rdlo_in(a2_wr[410]),  .coef_in(coef[616]), .rdup_out(a3_wr[154]), .rdlo_out(a3_wr[410]));
			radix2 #(.width(width)) rd_st2_155  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[155]), .rdlo_in(a2_wr[411]),  .coef_in(coef[620]), .rdup_out(a3_wr[155]), .rdlo_out(a3_wr[411]));
			radix2 #(.width(width)) rd_st2_156  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[156]), .rdlo_in(a2_wr[412]),  .coef_in(coef[624]), .rdup_out(a3_wr[156]), .rdlo_out(a3_wr[412]));
			radix2 #(.width(width)) rd_st2_157  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[157]), .rdlo_in(a2_wr[413]),  .coef_in(coef[628]), .rdup_out(a3_wr[157]), .rdlo_out(a3_wr[413]));
			radix2 #(.width(width)) rd_st2_158  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[158]), .rdlo_in(a2_wr[414]),  .coef_in(coef[632]), .rdup_out(a3_wr[158]), .rdlo_out(a3_wr[414]));
			radix2 #(.width(width)) rd_st2_159  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[159]), .rdlo_in(a2_wr[415]),  .coef_in(coef[636]), .rdup_out(a3_wr[159]), .rdlo_out(a3_wr[415]));
			radix2 #(.width(width)) rd_st2_160  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[160]), .rdlo_in(a2_wr[416]),  .coef_in(coef[640]), .rdup_out(a3_wr[160]), .rdlo_out(a3_wr[416]));
			radix2 #(.width(width)) rd_st2_161  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[161]), .rdlo_in(a2_wr[417]),  .coef_in(coef[644]), .rdup_out(a3_wr[161]), .rdlo_out(a3_wr[417]));
			radix2 #(.width(width)) rd_st2_162  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[162]), .rdlo_in(a2_wr[418]),  .coef_in(coef[648]), .rdup_out(a3_wr[162]), .rdlo_out(a3_wr[418]));
			radix2 #(.width(width)) rd_st2_163  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[163]), .rdlo_in(a2_wr[419]),  .coef_in(coef[652]), .rdup_out(a3_wr[163]), .rdlo_out(a3_wr[419]));
			radix2 #(.width(width)) rd_st2_164  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[164]), .rdlo_in(a2_wr[420]),  .coef_in(coef[656]), .rdup_out(a3_wr[164]), .rdlo_out(a3_wr[420]));
			radix2 #(.width(width)) rd_st2_165  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[165]), .rdlo_in(a2_wr[421]),  .coef_in(coef[660]), .rdup_out(a3_wr[165]), .rdlo_out(a3_wr[421]));
			radix2 #(.width(width)) rd_st2_166  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[166]), .rdlo_in(a2_wr[422]),  .coef_in(coef[664]), .rdup_out(a3_wr[166]), .rdlo_out(a3_wr[422]));
			radix2 #(.width(width)) rd_st2_167  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[167]), .rdlo_in(a2_wr[423]),  .coef_in(coef[668]), .rdup_out(a3_wr[167]), .rdlo_out(a3_wr[423]));
			radix2 #(.width(width)) rd_st2_168  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[168]), .rdlo_in(a2_wr[424]),  .coef_in(coef[672]), .rdup_out(a3_wr[168]), .rdlo_out(a3_wr[424]));
			radix2 #(.width(width)) rd_st2_169  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[169]), .rdlo_in(a2_wr[425]),  .coef_in(coef[676]), .rdup_out(a3_wr[169]), .rdlo_out(a3_wr[425]));
			radix2 #(.width(width)) rd_st2_170  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[170]), .rdlo_in(a2_wr[426]),  .coef_in(coef[680]), .rdup_out(a3_wr[170]), .rdlo_out(a3_wr[426]));
			radix2 #(.width(width)) rd_st2_171  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[171]), .rdlo_in(a2_wr[427]),  .coef_in(coef[684]), .rdup_out(a3_wr[171]), .rdlo_out(a3_wr[427]));
			radix2 #(.width(width)) rd_st2_172  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[172]), .rdlo_in(a2_wr[428]),  .coef_in(coef[688]), .rdup_out(a3_wr[172]), .rdlo_out(a3_wr[428]));
			radix2 #(.width(width)) rd_st2_173  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[173]), .rdlo_in(a2_wr[429]),  .coef_in(coef[692]), .rdup_out(a3_wr[173]), .rdlo_out(a3_wr[429]));
			radix2 #(.width(width)) rd_st2_174  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[174]), .rdlo_in(a2_wr[430]),  .coef_in(coef[696]), .rdup_out(a3_wr[174]), .rdlo_out(a3_wr[430]));
			radix2 #(.width(width)) rd_st2_175  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[175]), .rdlo_in(a2_wr[431]),  .coef_in(coef[700]), .rdup_out(a3_wr[175]), .rdlo_out(a3_wr[431]));
			radix2 #(.width(width)) rd_st2_176  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[176]), .rdlo_in(a2_wr[432]),  .coef_in(coef[704]), .rdup_out(a3_wr[176]), .rdlo_out(a3_wr[432]));
			radix2 #(.width(width)) rd_st2_177  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[177]), .rdlo_in(a2_wr[433]),  .coef_in(coef[708]), .rdup_out(a3_wr[177]), .rdlo_out(a3_wr[433]));
			radix2 #(.width(width)) rd_st2_178  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[178]), .rdlo_in(a2_wr[434]),  .coef_in(coef[712]), .rdup_out(a3_wr[178]), .rdlo_out(a3_wr[434]));
			radix2 #(.width(width)) rd_st2_179  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[179]), .rdlo_in(a2_wr[435]),  .coef_in(coef[716]), .rdup_out(a3_wr[179]), .rdlo_out(a3_wr[435]));
			radix2 #(.width(width)) rd_st2_180  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[180]), .rdlo_in(a2_wr[436]),  .coef_in(coef[720]), .rdup_out(a3_wr[180]), .rdlo_out(a3_wr[436]));
			radix2 #(.width(width)) rd_st2_181  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[181]), .rdlo_in(a2_wr[437]),  .coef_in(coef[724]), .rdup_out(a3_wr[181]), .rdlo_out(a3_wr[437]));
			radix2 #(.width(width)) rd_st2_182  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[182]), .rdlo_in(a2_wr[438]),  .coef_in(coef[728]), .rdup_out(a3_wr[182]), .rdlo_out(a3_wr[438]));
			radix2 #(.width(width)) rd_st2_183  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[183]), .rdlo_in(a2_wr[439]),  .coef_in(coef[732]), .rdup_out(a3_wr[183]), .rdlo_out(a3_wr[439]));
			radix2 #(.width(width)) rd_st2_184  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[184]), .rdlo_in(a2_wr[440]),  .coef_in(coef[736]), .rdup_out(a3_wr[184]), .rdlo_out(a3_wr[440]));
			radix2 #(.width(width)) rd_st2_185  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[185]), .rdlo_in(a2_wr[441]),  .coef_in(coef[740]), .rdup_out(a3_wr[185]), .rdlo_out(a3_wr[441]));
			radix2 #(.width(width)) rd_st2_186  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[186]), .rdlo_in(a2_wr[442]),  .coef_in(coef[744]), .rdup_out(a3_wr[186]), .rdlo_out(a3_wr[442]));
			radix2 #(.width(width)) rd_st2_187  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[187]), .rdlo_in(a2_wr[443]),  .coef_in(coef[748]), .rdup_out(a3_wr[187]), .rdlo_out(a3_wr[443]));
			radix2 #(.width(width)) rd_st2_188  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[188]), .rdlo_in(a2_wr[444]),  .coef_in(coef[752]), .rdup_out(a3_wr[188]), .rdlo_out(a3_wr[444]));
			radix2 #(.width(width)) rd_st2_189  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[189]), .rdlo_in(a2_wr[445]),  .coef_in(coef[756]), .rdup_out(a3_wr[189]), .rdlo_out(a3_wr[445]));
			radix2 #(.width(width)) rd_st2_190  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[190]), .rdlo_in(a2_wr[446]),  .coef_in(coef[760]), .rdup_out(a3_wr[190]), .rdlo_out(a3_wr[446]));
			radix2 #(.width(width)) rd_st2_191  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[191]), .rdlo_in(a2_wr[447]),  .coef_in(coef[764]), .rdup_out(a3_wr[191]), .rdlo_out(a3_wr[447]));
			radix2 #(.width(width)) rd_st2_192  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[192]), .rdlo_in(a2_wr[448]),  .coef_in(coef[768]), .rdup_out(a3_wr[192]), .rdlo_out(a3_wr[448]));
			radix2 #(.width(width)) rd_st2_193  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[193]), .rdlo_in(a2_wr[449]),  .coef_in(coef[772]), .rdup_out(a3_wr[193]), .rdlo_out(a3_wr[449]));
			radix2 #(.width(width)) rd_st2_194  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[194]), .rdlo_in(a2_wr[450]),  .coef_in(coef[776]), .rdup_out(a3_wr[194]), .rdlo_out(a3_wr[450]));
			radix2 #(.width(width)) rd_st2_195  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[195]), .rdlo_in(a2_wr[451]),  .coef_in(coef[780]), .rdup_out(a3_wr[195]), .rdlo_out(a3_wr[451]));
			radix2 #(.width(width)) rd_st2_196  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[196]), .rdlo_in(a2_wr[452]),  .coef_in(coef[784]), .rdup_out(a3_wr[196]), .rdlo_out(a3_wr[452]));
			radix2 #(.width(width)) rd_st2_197  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[197]), .rdlo_in(a2_wr[453]),  .coef_in(coef[788]), .rdup_out(a3_wr[197]), .rdlo_out(a3_wr[453]));
			radix2 #(.width(width)) rd_st2_198  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[198]), .rdlo_in(a2_wr[454]),  .coef_in(coef[792]), .rdup_out(a3_wr[198]), .rdlo_out(a3_wr[454]));
			radix2 #(.width(width)) rd_st2_199  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[199]), .rdlo_in(a2_wr[455]),  .coef_in(coef[796]), .rdup_out(a3_wr[199]), .rdlo_out(a3_wr[455]));
			radix2 #(.width(width)) rd_st2_200  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[200]), .rdlo_in(a2_wr[456]),  .coef_in(coef[800]), .rdup_out(a3_wr[200]), .rdlo_out(a3_wr[456]));
			radix2 #(.width(width)) rd_st2_201  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[201]), .rdlo_in(a2_wr[457]),  .coef_in(coef[804]), .rdup_out(a3_wr[201]), .rdlo_out(a3_wr[457]));
			radix2 #(.width(width)) rd_st2_202  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[202]), .rdlo_in(a2_wr[458]),  .coef_in(coef[808]), .rdup_out(a3_wr[202]), .rdlo_out(a3_wr[458]));
			radix2 #(.width(width)) rd_st2_203  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[203]), .rdlo_in(a2_wr[459]),  .coef_in(coef[812]), .rdup_out(a3_wr[203]), .rdlo_out(a3_wr[459]));
			radix2 #(.width(width)) rd_st2_204  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[204]), .rdlo_in(a2_wr[460]),  .coef_in(coef[816]), .rdup_out(a3_wr[204]), .rdlo_out(a3_wr[460]));
			radix2 #(.width(width)) rd_st2_205  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[205]), .rdlo_in(a2_wr[461]),  .coef_in(coef[820]), .rdup_out(a3_wr[205]), .rdlo_out(a3_wr[461]));
			radix2 #(.width(width)) rd_st2_206  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[206]), .rdlo_in(a2_wr[462]),  .coef_in(coef[824]), .rdup_out(a3_wr[206]), .rdlo_out(a3_wr[462]));
			radix2 #(.width(width)) rd_st2_207  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[207]), .rdlo_in(a2_wr[463]),  .coef_in(coef[828]), .rdup_out(a3_wr[207]), .rdlo_out(a3_wr[463]));
			radix2 #(.width(width)) rd_st2_208  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[208]), .rdlo_in(a2_wr[464]),  .coef_in(coef[832]), .rdup_out(a3_wr[208]), .rdlo_out(a3_wr[464]));
			radix2 #(.width(width)) rd_st2_209  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[209]), .rdlo_in(a2_wr[465]),  .coef_in(coef[836]), .rdup_out(a3_wr[209]), .rdlo_out(a3_wr[465]));
			radix2 #(.width(width)) rd_st2_210  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[210]), .rdlo_in(a2_wr[466]),  .coef_in(coef[840]), .rdup_out(a3_wr[210]), .rdlo_out(a3_wr[466]));
			radix2 #(.width(width)) rd_st2_211  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[211]), .rdlo_in(a2_wr[467]),  .coef_in(coef[844]), .rdup_out(a3_wr[211]), .rdlo_out(a3_wr[467]));
			radix2 #(.width(width)) rd_st2_212  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[212]), .rdlo_in(a2_wr[468]),  .coef_in(coef[848]), .rdup_out(a3_wr[212]), .rdlo_out(a3_wr[468]));
			radix2 #(.width(width)) rd_st2_213  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[213]), .rdlo_in(a2_wr[469]),  .coef_in(coef[852]), .rdup_out(a3_wr[213]), .rdlo_out(a3_wr[469]));
			radix2 #(.width(width)) rd_st2_214  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[214]), .rdlo_in(a2_wr[470]),  .coef_in(coef[856]), .rdup_out(a3_wr[214]), .rdlo_out(a3_wr[470]));
			radix2 #(.width(width)) rd_st2_215  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[215]), .rdlo_in(a2_wr[471]),  .coef_in(coef[860]), .rdup_out(a3_wr[215]), .rdlo_out(a3_wr[471]));
			radix2 #(.width(width)) rd_st2_216  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[216]), .rdlo_in(a2_wr[472]),  .coef_in(coef[864]), .rdup_out(a3_wr[216]), .rdlo_out(a3_wr[472]));
			radix2 #(.width(width)) rd_st2_217  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[217]), .rdlo_in(a2_wr[473]),  .coef_in(coef[868]), .rdup_out(a3_wr[217]), .rdlo_out(a3_wr[473]));
			radix2 #(.width(width)) rd_st2_218  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[218]), .rdlo_in(a2_wr[474]),  .coef_in(coef[872]), .rdup_out(a3_wr[218]), .rdlo_out(a3_wr[474]));
			radix2 #(.width(width)) rd_st2_219  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[219]), .rdlo_in(a2_wr[475]),  .coef_in(coef[876]), .rdup_out(a3_wr[219]), .rdlo_out(a3_wr[475]));
			radix2 #(.width(width)) rd_st2_220  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[220]), .rdlo_in(a2_wr[476]),  .coef_in(coef[880]), .rdup_out(a3_wr[220]), .rdlo_out(a3_wr[476]));
			radix2 #(.width(width)) rd_st2_221  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[221]), .rdlo_in(a2_wr[477]),  .coef_in(coef[884]), .rdup_out(a3_wr[221]), .rdlo_out(a3_wr[477]));
			radix2 #(.width(width)) rd_st2_222  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[222]), .rdlo_in(a2_wr[478]),  .coef_in(coef[888]), .rdup_out(a3_wr[222]), .rdlo_out(a3_wr[478]));
			radix2 #(.width(width)) rd_st2_223  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[223]), .rdlo_in(a2_wr[479]),  .coef_in(coef[892]), .rdup_out(a3_wr[223]), .rdlo_out(a3_wr[479]));
			radix2 #(.width(width)) rd_st2_224  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[224]), .rdlo_in(a2_wr[480]),  .coef_in(coef[896]), .rdup_out(a3_wr[224]), .rdlo_out(a3_wr[480]));
			radix2 #(.width(width)) rd_st2_225  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[225]), .rdlo_in(a2_wr[481]),  .coef_in(coef[900]), .rdup_out(a3_wr[225]), .rdlo_out(a3_wr[481]));
			radix2 #(.width(width)) rd_st2_226  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[226]), .rdlo_in(a2_wr[482]),  .coef_in(coef[904]), .rdup_out(a3_wr[226]), .rdlo_out(a3_wr[482]));
			radix2 #(.width(width)) rd_st2_227  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[227]), .rdlo_in(a2_wr[483]),  .coef_in(coef[908]), .rdup_out(a3_wr[227]), .rdlo_out(a3_wr[483]));
			radix2 #(.width(width)) rd_st2_228  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[228]), .rdlo_in(a2_wr[484]),  .coef_in(coef[912]), .rdup_out(a3_wr[228]), .rdlo_out(a3_wr[484]));
			radix2 #(.width(width)) rd_st2_229  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[229]), .rdlo_in(a2_wr[485]),  .coef_in(coef[916]), .rdup_out(a3_wr[229]), .rdlo_out(a3_wr[485]));
			radix2 #(.width(width)) rd_st2_230  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[230]), .rdlo_in(a2_wr[486]),  .coef_in(coef[920]), .rdup_out(a3_wr[230]), .rdlo_out(a3_wr[486]));
			radix2 #(.width(width)) rd_st2_231  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[231]), .rdlo_in(a2_wr[487]),  .coef_in(coef[924]), .rdup_out(a3_wr[231]), .rdlo_out(a3_wr[487]));
			radix2 #(.width(width)) rd_st2_232  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[232]), .rdlo_in(a2_wr[488]),  .coef_in(coef[928]), .rdup_out(a3_wr[232]), .rdlo_out(a3_wr[488]));
			radix2 #(.width(width)) rd_st2_233  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[233]), .rdlo_in(a2_wr[489]),  .coef_in(coef[932]), .rdup_out(a3_wr[233]), .rdlo_out(a3_wr[489]));
			radix2 #(.width(width)) rd_st2_234  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[234]), .rdlo_in(a2_wr[490]),  .coef_in(coef[936]), .rdup_out(a3_wr[234]), .rdlo_out(a3_wr[490]));
			radix2 #(.width(width)) rd_st2_235  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[235]), .rdlo_in(a2_wr[491]),  .coef_in(coef[940]), .rdup_out(a3_wr[235]), .rdlo_out(a3_wr[491]));
			radix2 #(.width(width)) rd_st2_236  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[236]), .rdlo_in(a2_wr[492]),  .coef_in(coef[944]), .rdup_out(a3_wr[236]), .rdlo_out(a3_wr[492]));
			radix2 #(.width(width)) rd_st2_237  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[237]), .rdlo_in(a2_wr[493]),  .coef_in(coef[948]), .rdup_out(a3_wr[237]), .rdlo_out(a3_wr[493]));
			radix2 #(.width(width)) rd_st2_238  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[238]), .rdlo_in(a2_wr[494]),  .coef_in(coef[952]), .rdup_out(a3_wr[238]), .rdlo_out(a3_wr[494]));
			radix2 #(.width(width)) rd_st2_239  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[239]), .rdlo_in(a2_wr[495]),  .coef_in(coef[956]), .rdup_out(a3_wr[239]), .rdlo_out(a3_wr[495]));
			radix2 #(.width(width)) rd_st2_240  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[240]), .rdlo_in(a2_wr[496]),  .coef_in(coef[960]), .rdup_out(a3_wr[240]), .rdlo_out(a3_wr[496]));
			radix2 #(.width(width)) rd_st2_241  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[241]), .rdlo_in(a2_wr[497]),  .coef_in(coef[964]), .rdup_out(a3_wr[241]), .rdlo_out(a3_wr[497]));
			radix2 #(.width(width)) rd_st2_242  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[242]), .rdlo_in(a2_wr[498]),  .coef_in(coef[968]), .rdup_out(a3_wr[242]), .rdlo_out(a3_wr[498]));
			radix2 #(.width(width)) rd_st2_243  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[243]), .rdlo_in(a2_wr[499]),  .coef_in(coef[972]), .rdup_out(a3_wr[243]), .rdlo_out(a3_wr[499]));
			radix2 #(.width(width)) rd_st2_244  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[244]), .rdlo_in(a2_wr[500]),  .coef_in(coef[976]), .rdup_out(a3_wr[244]), .rdlo_out(a3_wr[500]));
			radix2 #(.width(width)) rd_st2_245  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[245]), .rdlo_in(a2_wr[501]),  .coef_in(coef[980]), .rdup_out(a3_wr[245]), .rdlo_out(a3_wr[501]));
			radix2 #(.width(width)) rd_st2_246  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[246]), .rdlo_in(a2_wr[502]),  .coef_in(coef[984]), .rdup_out(a3_wr[246]), .rdlo_out(a3_wr[502]));
			radix2 #(.width(width)) rd_st2_247  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[247]), .rdlo_in(a2_wr[503]),  .coef_in(coef[988]), .rdup_out(a3_wr[247]), .rdlo_out(a3_wr[503]));
			radix2 #(.width(width)) rd_st2_248  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[248]), .rdlo_in(a2_wr[504]),  .coef_in(coef[992]), .rdup_out(a3_wr[248]), .rdlo_out(a3_wr[504]));
			radix2 #(.width(width)) rd_st2_249  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[249]), .rdlo_in(a2_wr[505]),  .coef_in(coef[996]), .rdup_out(a3_wr[249]), .rdlo_out(a3_wr[505]));
			radix2 #(.width(width)) rd_st2_250  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[250]), .rdlo_in(a2_wr[506]),  .coef_in(coef[1000]), .rdup_out(a3_wr[250]), .rdlo_out(a3_wr[506]));
			radix2 #(.width(width)) rd_st2_251  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[251]), .rdlo_in(a2_wr[507]),  .coef_in(coef[1004]), .rdup_out(a3_wr[251]), .rdlo_out(a3_wr[507]));
			radix2 #(.width(width)) rd_st2_252  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[252]), .rdlo_in(a2_wr[508]),  .coef_in(coef[1008]), .rdup_out(a3_wr[252]), .rdlo_out(a3_wr[508]));
			radix2 #(.width(width)) rd_st2_253  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[253]), .rdlo_in(a2_wr[509]),  .coef_in(coef[1012]), .rdup_out(a3_wr[253]), .rdlo_out(a3_wr[509]));
			radix2 #(.width(width)) rd_st2_254  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[254]), .rdlo_in(a2_wr[510]),  .coef_in(coef[1016]), .rdup_out(a3_wr[254]), .rdlo_out(a3_wr[510]));
			radix2 #(.width(width)) rd_st2_255  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[255]), .rdlo_in(a2_wr[511]),  .coef_in(coef[1020]), .rdup_out(a3_wr[255]), .rdlo_out(a3_wr[511]));
			radix2 #(.width(width)) rd_st2_512  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[512]), .rdlo_in(a2_wr[768]),  .coef_in(coef[0]), .rdup_out(a3_wr[512]), .rdlo_out(a3_wr[768]));
			radix2 #(.width(width)) rd_st2_513  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[513]), .rdlo_in(a2_wr[769]),  .coef_in(coef[4]), .rdup_out(a3_wr[513]), .rdlo_out(a3_wr[769]));
			radix2 #(.width(width)) rd_st2_514  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[514]), .rdlo_in(a2_wr[770]),  .coef_in(coef[8]), .rdup_out(a3_wr[514]), .rdlo_out(a3_wr[770]));
			radix2 #(.width(width)) rd_st2_515  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[515]), .rdlo_in(a2_wr[771]),  .coef_in(coef[12]), .rdup_out(a3_wr[515]), .rdlo_out(a3_wr[771]));
			radix2 #(.width(width)) rd_st2_516  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[516]), .rdlo_in(a2_wr[772]),  .coef_in(coef[16]), .rdup_out(a3_wr[516]), .rdlo_out(a3_wr[772]));
			radix2 #(.width(width)) rd_st2_517  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[517]), .rdlo_in(a2_wr[773]),  .coef_in(coef[20]), .rdup_out(a3_wr[517]), .rdlo_out(a3_wr[773]));
			radix2 #(.width(width)) rd_st2_518  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[518]), .rdlo_in(a2_wr[774]),  .coef_in(coef[24]), .rdup_out(a3_wr[518]), .rdlo_out(a3_wr[774]));
			radix2 #(.width(width)) rd_st2_519  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[519]), .rdlo_in(a2_wr[775]),  .coef_in(coef[28]), .rdup_out(a3_wr[519]), .rdlo_out(a3_wr[775]));
			radix2 #(.width(width)) rd_st2_520  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[520]), .rdlo_in(a2_wr[776]),  .coef_in(coef[32]), .rdup_out(a3_wr[520]), .rdlo_out(a3_wr[776]));
			radix2 #(.width(width)) rd_st2_521  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[521]), .rdlo_in(a2_wr[777]),  .coef_in(coef[36]), .rdup_out(a3_wr[521]), .rdlo_out(a3_wr[777]));
			radix2 #(.width(width)) rd_st2_522  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[522]), .rdlo_in(a2_wr[778]),  .coef_in(coef[40]), .rdup_out(a3_wr[522]), .rdlo_out(a3_wr[778]));
			radix2 #(.width(width)) rd_st2_523  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[523]), .rdlo_in(a2_wr[779]),  .coef_in(coef[44]), .rdup_out(a3_wr[523]), .rdlo_out(a3_wr[779]));
			radix2 #(.width(width)) rd_st2_524  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[524]), .rdlo_in(a2_wr[780]),  .coef_in(coef[48]), .rdup_out(a3_wr[524]), .rdlo_out(a3_wr[780]));
			radix2 #(.width(width)) rd_st2_525  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[525]), .rdlo_in(a2_wr[781]),  .coef_in(coef[52]), .rdup_out(a3_wr[525]), .rdlo_out(a3_wr[781]));
			radix2 #(.width(width)) rd_st2_526  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[526]), .rdlo_in(a2_wr[782]),  .coef_in(coef[56]), .rdup_out(a3_wr[526]), .rdlo_out(a3_wr[782]));
			radix2 #(.width(width)) rd_st2_527  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[527]), .rdlo_in(a2_wr[783]),  .coef_in(coef[60]), .rdup_out(a3_wr[527]), .rdlo_out(a3_wr[783]));
			radix2 #(.width(width)) rd_st2_528  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[528]), .rdlo_in(a2_wr[784]),  .coef_in(coef[64]), .rdup_out(a3_wr[528]), .rdlo_out(a3_wr[784]));
			radix2 #(.width(width)) rd_st2_529  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[529]), .rdlo_in(a2_wr[785]),  .coef_in(coef[68]), .rdup_out(a3_wr[529]), .rdlo_out(a3_wr[785]));
			radix2 #(.width(width)) rd_st2_530  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[530]), .rdlo_in(a2_wr[786]),  .coef_in(coef[72]), .rdup_out(a3_wr[530]), .rdlo_out(a3_wr[786]));
			radix2 #(.width(width)) rd_st2_531  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[531]), .rdlo_in(a2_wr[787]),  .coef_in(coef[76]), .rdup_out(a3_wr[531]), .rdlo_out(a3_wr[787]));
			radix2 #(.width(width)) rd_st2_532  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[532]), .rdlo_in(a2_wr[788]),  .coef_in(coef[80]), .rdup_out(a3_wr[532]), .rdlo_out(a3_wr[788]));
			radix2 #(.width(width)) rd_st2_533  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[533]), .rdlo_in(a2_wr[789]),  .coef_in(coef[84]), .rdup_out(a3_wr[533]), .rdlo_out(a3_wr[789]));
			radix2 #(.width(width)) rd_st2_534  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[534]), .rdlo_in(a2_wr[790]),  .coef_in(coef[88]), .rdup_out(a3_wr[534]), .rdlo_out(a3_wr[790]));
			radix2 #(.width(width)) rd_st2_535  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[535]), .rdlo_in(a2_wr[791]),  .coef_in(coef[92]), .rdup_out(a3_wr[535]), .rdlo_out(a3_wr[791]));
			radix2 #(.width(width)) rd_st2_536  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[536]), .rdlo_in(a2_wr[792]),  .coef_in(coef[96]), .rdup_out(a3_wr[536]), .rdlo_out(a3_wr[792]));
			radix2 #(.width(width)) rd_st2_537  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[537]), .rdlo_in(a2_wr[793]),  .coef_in(coef[100]), .rdup_out(a3_wr[537]), .rdlo_out(a3_wr[793]));
			radix2 #(.width(width)) rd_st2_538  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[538]), .rdlo_in(a2_wr[794]),  .coef_in(coef[104]), .rdup_out(a3_wr[538]), .rdlo_out(a3_wr[794]));
			radix2 #(.width(width)) rd_st2_539  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[539]), .rdlo_in(a2_wr[795]),  .coef_in(coef[108]), .rdup_out(a3_wr[539]), .rdlo_out(a3_wr[795]));
			radix2 #(.width(width)) rd_st2_540  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[540]), .rdlo_in(a2_wr[796]),  .coef_in(coef[112]), .rdup_out(a3_wr[540]), .rdlo_out(a3_wr[796]));
			radix2 #(.width(width)) rd_st2_541  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[541]), .rdlo_in(a2_wr[797]),  .coef_in(coef[116]), .rdup_out(a3_wr[541]), .rdlo_out(a3_wr[797]));
			radix2 #(.width(width)) rd_st2_542  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[542]), .rdlo_in(a2_wr[798]),  .coef_in(coef[120]), .rdup_out(a3_wr[542]), .rdlo_out(a3_wr[798]));
			radix2 #(.width(width)) rd_st2_543  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[543]), .rdlo_in(a2_wr[799]),  .coef_in(coef[124]), .rdup_out(a3_wr[543]), .rdlo_out(a3_wr[799]));
			radix2 #(.width(width)) rd_st2_544  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[544]), .rdlo_in(a2_wr[800]),  .coef_in(coef[128]), .rdup_out(a3_wr[544]), .rdlo_out(a3_wr[800]));
			radix2 #(.width(width)) rd_st2_545  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[545]), .rdlo_in(a2_wr[801]),  .coef_in(coef[132]), .rdup_out(a3_wr[545]), .rdlo_out(a3_wr[801]));
			radix2 #(.width(width)) rd_st2_546  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[546]), .rdlo_in(a2_wr[802]),  .coef_in(coef[136]), .rdup_out(a3_wr[546]), .rdlo_out(a3_wr[802]));
			radix2 #(.width(width)) rd_st2_547  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[547]), .rdlo_in(a2_wr[803]),  .coef_in(coef[140]), .rdup_out(a3_wr[547]), .rdlo_out(a3_wr[803]));
			radix2 #(.width(width)) rd_st2_548  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[548]), .rdlo_in(a2_wr[804]),  .coef_in(coef[144]), .rdup_out(a3_wr[548]), .rdlo_out(a3_wr[804]));
			radix2 #(.width(width)) rd_st2_549  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[549]), .rdlo_in(a2_wr[805]),  .coef_in(coef[148]), .rdup_out(a3_wr[549]), .rdlo_out(a3_wr[805]));
			radix2 #(.width(width)) rd_st2_550  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[550]), .rdlo_in(a2_wr[806]),  .coef_in(coef[152]), .rdup_out(a3_wr[550]), .rdlo_out(a3_wr[806]));
			radix2 #(.width(width)) rd_st2_551  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[551]), .rdlo_in(a2_wr[807]),  .coef_in(coef[156]), .rdup_out(a3_wr[551]), .rdlo_out(a3_wr[807]));
			radix2 #(.width(width)) rd_st2_552  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[552]), .rdlo_in(a2_wr[808]),  .coef_in(coef[160]), .rdup_out(a3_wr[552]), .rdlo_out(a3_wr[808]));
			radix2 #(.width(width)) rd_st2_553  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[553]), .rdlo_in(a2_wr[809]),  .coef_in(coef[164]), .rdup_out(a3_wr[553]), .rdlo_out(a3_wr[809]));
			radix2 #(.width(width)) rd_st2_554  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[554]), .rdlo_in(a2_wr[810]),  .coef_in(coef[168]), .rdup_out(a3_wr[554]), .rdlo_out(a3_wr[810]));
			radix2 #(.width(width)) rd_st2_555  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[555]), .rdlo_in(a2_wr[811]),  .coef_in(coef[172]), .rdup_out(a3_wr[555]), .rdlo_out(a3_wr[811]));
			radix2 #(.width(width)) rd_st2_556  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[556]), .rdlo_in(a2_wr[812]),  .coef_in(coef[176]), .rdup_out(a3_wr[556]), .rdlo_out(a3_wr[812]));
			radix2 #(.width(width)) rd_st2_557  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[557]), .rdlo_in(a2_wr[813]),  .coef_in(coef[180]), .rdup_out(a3_wr[557]), .rdlo_out(a3_wr[813]));
			radix2 #(.width(width)) rd_st2_558  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[558]), .rdlo_in(a2_wr[814]),  .coef_in(coef[184]), .rdup_out(a3_wr[558]), .rdlo_out(a3_wr[814]));
			radix2 #(.width(width)) rd_st2_559  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[559]), .rdlo_in(a2_wr[815]),  .coef_in(coef[188]), .rdup_out(a3_wr[559]), .rdlo_out(a3_wr[815]));
			radix2 #(.width(width)) rd_st2_560  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[560]), .rdlo_in(a2_wr[816]),  .coef_in(coef[192]), .rdup_out(a3_wr[560]), .rdlo_out(a3_wr[816]));
			radix2 #(.width(width)) rd_st2_561  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[561]), .rdlo_in(a2_wr[817]),  .coef_in(coef[196]), .rdup_out(a3_wr[561]), .rdlo_out(a3_wr[817]));
			radix2 #(.width(width)) rd_st2_562  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[562]), .rdlo_in(a2_wr[818]),  .coef_in(coef[200]), .rdup_out(a3_wr[562]), .rdlo_out(a3_wr[818]));
			radix2 #(.width(width)) rd_st2_563  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[563]), .rdlo_in(a2_wr[819]),  .coef_in(coef[204]), .rdup_out(a3_wr[563]), .rdlo_out(a3_wr[819]));
			radix2 #(.width(width)) rd_st2_564  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[564]), .rdlo_in(a2_wr[820]),  .coef_in(coef[208]), .rdup_out(a3_wr[564]), .rdlo_out(a3_wr[820]));
			radix2 #(.width(width)) rd_st2_565  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[565]), .rdlo_in(a2_wr[821]),  .coef_in(coef[212]), .rdup_out(a3_wr[565]), .rdlo_out(a3_wr[821]));
			radix2 #(.width(width)) rd_st2_566  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[566]), .rdlo_in(a2_wr[822]),  .coef_in(coef[216]), .rdup_out(a3_wr[566]), .rdlo_out(a3_wr[822]));
			radix2 #(.width(width)) rd_st2_567  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[567]), .rdlo_in(a2_wr[823]),  .coef_in(coef[220]), .rdup_out(a3_wr[567]), .rdlo_out(a3_wr[823]));
			radix2 #(.width(width)) rd_st2_568  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[568]), .rdlo_in(a2_wr[824]),  .coef_in(coef[224]), .rdup_out(a3_wr[568]), .rdlo_out(a3_wr[824]));
			radix2 #(.width(width)) rd_st2_569  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[569]), .rdlo_in(a2_wr[825]),  .coef_in(coef[228]), .rdup_out(a3_wr[569]), .rdlo_out(a3_wr[825]));
			radix2 #(.width(width)) rd_st2_570  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[570]), .rdlo_in(a2_wr[826]),  .coef_in(coef[232]), .rdup_out(a3_wr[570]), .rdlo_out(a3_wr[826]));
			radix2 #(.width(width)) rd_st2_571  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[571]), .rdlo_in(a2_wr[827]),  .coef_in(coef[236]), .rdup_out(a3_wr[571]), .rdlo_out(a3_wr[827]));
			radix2 #(.width(width)) rd_st2_572  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[572]), .rdlo_in(a2_wr[828]),  .coef_in(coef[240]), .rdup_out(a3_wr[572]), .rdlo_out(a3_wr[828]));
			radix2 #(.width(width)) rd_st2_573  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[573]), .rdlo_in(a2_wr[829]),  .coef_in(coef[244]), .rdup_out(a3_wr[573]), .rdlo_out(a3_wr[829]));
			radix2 #(.width(width)) rd_st2_574  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[574]), .rdlo_in(a2_wr[830]),  .coef_in(coef[248]), .rdup_out(a3_wr[574]), .rdlo_out(a3_wr[830]));
			radix2 #(.width(width)) rd_st2_575  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[575]), .rdlo_in(a2_wr[831]),  .coef_in(coef[252]), .rdup_out(a3_wr[575]), .rdlo_out(a3_wr[831]));
			radix2 #(.width(width)) rd_st2_576  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[576]), .rdlo_in(a2_wr[832]),  .coef_in(coef[256]), .rdup_out(a3_wr[576]), .rdlo_out(a3_wr[832]));
			radix2 #(.width(width)) rd_st2_577  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[577]), .rdlo_in(a2_wr[833]),  .coef_in(coef[260]), .rdup_out(a3_wr[577]), .rdlo_out(a3_wr[833]));
			radix2 #(.width(width)) rd_st2_578  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[578]), .rdlo_in(a2_wr[834]),  .coef_in(coef[264]), .rdup_out(a3_wr[578]), .rdlo_out(a3_wr[834]));
			radix2 #(.width(width)) rd_st2_579  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[579]), .rdlo_in(a2_wr[835]),  .coef_in(coef[268]), .rdup_out(a3_wr[579]), .rdlo_out(a3_wr[835]));
			radix2 #(.width(width)) rd_st2_580  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[580]), .rdlo_in(a2_wr[836]),  .coef_in(coef[272]), .rdup_out(a3_wr[580]), .rdlo_out(a3_wr[836]));
			radix2 #(.width(width)) rd_st2_581  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[581]), .rdlo_in(a2_wr[837]),  .coef_in(coef[276]), .rdup_out(a3_wr[581]), .rdlo_out(a3_wr[837]));
			radix2 #(.width(width)) rd_st2_582  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[582]), .rdlo_in(a2_wr[838]),  .coef_in(coef[280]), .rdup_out(a3_wr[582]), .rdlo_out(a3_wr[838]));
			radix2 #(.width(width)) rd_st2_583  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[583]), .rdlo_in(a2_wr[839]),  .coef_in(coef[284]), .rdup_out(a3_wr[583]), .rdlo_out(a3_wr[839]));
			radix2 #(.width(width)) rd_st2_584  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[584]), .rdlo_in(a2_wr[840]),  .coef_in(coef[288]), .rdup_out(a3_wr[584]), .rdlo_out(a3_wr[840]));
			radix2 #(.width(width)) rd_st2_585  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[585]), .rdlo_in(a2_wr[841]),  .coef_in(coef[292]), .rdup_out(a3_wr[585]), .rdlo_out(a3_wr[841]));
			radix2 #(.width(width)) rd_st2_586  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[586]), .rdlo_in(a2_wr[842]),  .coef_in(coef[296]), .rdup_out(a3_wr[586]), .rdlo_out(a3_wr[842]));
			radix2 #(.width(width)) rd_st2_587  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[587]), .rdlo_in(a2_wr[843]),  .coef_in(coef[300]), .rdup_out(a3_wr[587]), .rdlo_out(a3_wr[843]));
			radix2 #(.width(width)) rd_st2_588  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[588]), .rdlo_in(a2_wr[844]),  .coef_in(coef[304]), .rdup_out(a3_wr[588]), .rdlo_out(a3_wr[844]));
			radix2 #(.width(width)) rd_st2_589  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[589]), .rdlo_in(a2_wr[845]),  .coef_in(coef[308]), .rdup_out(a3_wr[589]), .rdlo_out(a3_wr[845]));
			radix2 #(.width(width)) rd_st2_590  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[590]), .rdlo_in(a2_wr[846]),  .coef_in(coef[312]), .rdup_out(a3_wr[590]), .rdlo_out(a3_wr[846]));
			radix2 #(.width(width)) rd_st2_591  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[591]), .rdlo_in(a2_wr[847]),  .coef_in(coef[316]), .rdup_out(a3_wr[591]), .rdlo_out(a3_wr[847]));
			radix2 #(.width(width)) rd_st2_592  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[592]), .rdlo_in(a2_wr[848]),  .coef_in(coef[320]), .rdup_out(a3_wr[592]), .rdlo_out(a3_wr[848]));
			radix2 #(.width(width)) rd_st2_593  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[593]), .rdlo_in(a2_wr[849]),  .coef_in(coef[324]), .rdup_out(a3_wr[593]), .rdlo_out(a3_wr[849]));
			radix2 #(.width(width)) rd_st2_594  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[594]), .rdlo_in(a2_wr[850]),  .coef_in(coef[328]), .rdup_out(a3_wr[594]), .rdlo_out(a3_wr[850]));
			radix2 #(.width(width)) rd_st2_595  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[595]), .rdlo_in(a2_wr[851]),  .coef_in(coef[332]), .rdup_out(a3_wr[595]), .rdlo_out(a3_wr[851]));
			radix2 #(.width(width)) rd_st2_596  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[596]), .rdlo_in(a2_wr[852]),  .coef_in(coef[336]), .rdup_out(a3_wr[596]), .rdlo_out(a3_wr[852]));
			radix2 #(.width(width)) rd_st2_597  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[597]), .rdlo_in(a2_wr[853]),  .coef_in(coef[340]), .rdup_out(a3_wr[597]), .rdlo_out(a3_wr[853]));
			radix2 #(.width(width)) rd_st2_598  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[598]), .rdlo_in(a2_wr[854]),  .coef_in(coef[344]), .rdup_out(a3_wr[598]), .rdlo_out(a3_wr[854]));
			radix2 #(.width(width)) rd_st2_599  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[599]), .rdlo_in(a2_wr[855]),  .coef_in(coef[348]), .rdup_out(a3_wr[599]), .rdlo_out(a3_wr[855]));
			radix2 #(.width(width)) rd_st2_600  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[600]), .rdlo_in(a2_wr[856]),  .coef_in(coef[352]), .rdup_out(a3_wr[600]), .rdlo_out(a3_wr[856]));
			radix2 #(.width(width)) rd_st2_601  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[601]), .rdlo_in(a2_wr[857]),  .coef_in(coef[356]), .rdup_out(a3_wr[601]), .rdlo_out(a3_wr[857]));
			radix2 #(.width(width)) rd_st2_602  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[602]), .rdlo_in(a2_wr[858]),  .coef_in(coef[360]), .rdup_out(a3_wr[602]), .rdlo_out(a3_wr[858]));
			radix2 #(.width(width)) rd_st2_603  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[603]), .rdlo_in(a2_wr[859]),  .coef_in(coef[364]), .rdup_out(a3_wr[603]), .rdlo_out(a3_wr[859]));
			radix2 #(.width(width)) rd_st2_604  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[604]), .rdlo_in(a2_wr[860]),  .coef_in(coef[368]), .rdup_out(a3_wr[604]), .rdlo_out(a3_wr[860]));
			radix2 #(.width(width)) rd_st2_605  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[605]), .rdlo_in(a2_wr[861]),  .coef_in(coef[372]), .rdup_out(a3_wr[605]), .rdlo_out(a3_wr[861]));
			radix2 #(.width(width)) rd_st2_606  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[606]), .rdlo_in(a2_wr[862]),  .coef_in(coef[376]), .rdup_out(a3_wr[606]), .rdlo_out(a3_wr[862]));
			radix2 #(.width(width)) rd_st2_607  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[607]), .rdlo_in(a2_wr[863]),  .coef_in(coef[380]), .rdup_out(a3_wr[607]), .rdlo_out(a3_wr[863]));
			radix2 #(.width(width)) rd_st2_608  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[608]), .rdlo_in(a2_wr[864]),  .coef_in(coef[384]), .rdup_out(a3_wr[608]), .rdlo_out(a3_wr[864]));
			radix2 #(.width(width)) rd_st2_609  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[609]), .rdlo_in(a2_wr[865]),  .coef_in(coef[388]), .rdup_out(a3_wr[609]), .rdlo_out(a3_wr[865]));
			radix2 #(.width(width)) rd_st2_610  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[610]), .rdlo_in(a2_wr[866]),  .coef_in(coef[392]), .rdup_out(a3_wr[610]), .rdlo_out(a3_wr[866]));
			radix2 #(.width(width)) rd_st2_611  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[611]), .rdlo_in(a2_wr[867]),  .coef_in(coef[396]), .rdup_out(a3_wr[611]), .rdlo_out(a3_wr[867]));
			radix2 #(.width(width)) rd_st2_612  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[612]), .rdlo_in(a2_wr[868]),  .coef_in(coef[400]), .rdup_out(a3_wr[612]), .rdlo_out(a3_wr[868]));
			radix2 #(.width(width)) rd_st2_613  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[613]), .rdlo_in(a2_wr[869]),  .coef_in(coef[404]), .rdup_out(a3_wr[613]), .rdlo_out(a3_wr[869]));
			radix2 #(.width(width)) rd_st2_614  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[614]), .rdlo_in(a2_wr[870]),  .coef_in(coef[408]), .rdup_out(a3_wr[614]), .rdlo_out(a3_wr[870]));
			radix2 #(.width(width)) rd_st2_615  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[615]), .rdlo_in(a2_wr[871]),  .coef_in(coef[412]), .rdup_out(a3_wr[615]), .rdlo_out(a3_wr[871]));
			radix2 #(.width(width)) rd_st2_616  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[616]), .rdlo_in(a2_wr[872]),  .coef_in(coef[416]), .rdup_out(a3_wr[616]), .rdlo_out(a3_wr[872]));
			radix2 #(.width(width)) rd_st2_617  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[617]), .rdlo_in(a2_wr[873]),  .coef_in(coef[420]), .rdup_out(a3_wr[617]), .rdlo_out(a3_wr[873]));
			radix2 #(.width(width)) rd_st2_618  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[618]), .rdlo_in(a2_wr[874]),  .coef_in(coef[424]), .rdup_out(a3_wr[618]), .rdlo_out(a3_wr[874]));
			radix2 #(.width(width)) rd_st2_619  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[619]), .rdlo_in(a2_wr[875]),  .coef_in(coef[428]), .rdup_out(a3_wr[619]), .rdlo_out(a3_wr[875]));
			radix2 #(.width(width)) rd_st2_620  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[620]), .rdlo_in(a2_wr[876]),  .coef_in(coef[432]), .rdup_out(a3_wr[620]), .rdlo_out(a3_wr[876]));
			radix2 #(.width(width)) rd_st2_621  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[621]), .rdlo_in(a2_wr[877]),  .coef_in(coef[436]), .rdup_out(a3_wr[621]), .rdlo_out(a3_wr[877]));
			radix2 #(.width(width)) rd_st2_622  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[622]), .rdlo_in(a2_wr[878]),  .coef_in(coef[440]), .rdup_out(a3_wr[622]), .rdlo_out(a3_wr[878]));
			radix2 #(.width(width)) rd_st2_623  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[623]), .rdlo_in(a2_wr[879]),  .coef_in(coef[444]), .rdup_out(a3_wr[623]), .rdlo_out(a3_wr[879]));
			radix2 #(.width(width)) rd_st2_624  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[624]), .rdlo_in(a2_wr[880]),  .coef_in(coef[448]), .rdup_out(a3_wr[624]), .rdlo_out(a3_wr[880]));
			radix2 #(.width(width)) rd_st2_625  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[625]), .rdlo_in(a2_wr[881]),  .coef_in(coef[452]), .rdup_out(a3_wr[625]), .rdlo_out(a3_wr[881]));
			radix2 #(.width(width)) rd_st2_626  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[626]), .rdlo_in(a2_wr[882]),  .coef_in(coef[456]), .rdup_out(a3_wr[626]), .rdlo_out(a3_wr[882]));
			radix2 #(.width(width)) rd_st2_627  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[627]), .rdlo_in(a2_wr[883]),  .coef_in(coef[460]), .rdup_out(a3_wr[627]), .rdlo_out(a3_wr[883]));
			radix2 #(.width(width)) rd_st2_628  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[628]), .rdlo_in(a2_wr[884]),  .coef_in(coef[464]), .rdup_out(a3_wr[628]), .rdlo_out(a3_wr[884]));
			radix2 #(.width(width)) rd_st2_629  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[629]), .rdlo_in(a2_wr[885]),  .coef_in(coef[468]), .rdup_out(a3_wr[629]), .rdlo_out(a3_wr[885]));
			radix2 #(.width(width)) rd_st2_630  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[630]), .rdlo_in(a2_wr[886]),  .coef_in(coef[472]), .rdup_out(a3_wr[630]), .rdlo_out(a3_wr[886]));
			radix2 #(.width(width)) rd_st2_631  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[631]), .rdlo_in(a2_wr[887]),  .coef_in(coef[476]), .rdup_out(a3_wr[631]), .rdlo_out(a3_wr[887]));
			radix2 #(.width(width)) rd_st2_632  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[632]), .rdlo_in(a2_wr[888]),  .coef_in(coef[480]), .rdup_out(a3_wr[632]), .rdlo_out(a3_wr[888]));
			radix2 #(.width(width)) rd_st2_633  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[633]), .rdlo_in(a2_wr[889]),  .coef_in(coef[484]), .rdup_out(a3_wr[633]), .rdlo_out(a3_wr[889]));
			radix2 #(.width(width)) rd_st2_634  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[634]), .rdlo_in(a2_wr[890]),  .coef_in(coef[488]), .rdup_out(a3_wr[634]), .rdlo_out(a3_wr[890]));
			radix2 #(.width(width)) rd_st2_635  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[635]), .rdlo_in(a2_wr[891]),  .coef_in(coef[492]), .rdup_out(a3_wr[635]), .rdlo_out(a3_wr[891]));
			radix2 #(.width(width)) rd_st2_636  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[636]), .rdlo_in(a2_wr[892]),  .coef_in(coef[496]), .rdup_out(a3_wr[636]), .rdlo_out(a3_wr[892]));
			radix2 #(.width(width)) rd_st2_637  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[637]), .rdlo_in(a2_wr[893]),  .coef_in(coef[500]), .rdup_out(a3_wr[637]), .rdlo_out(a3_wr[893]));
			radix2 #(.width(width)) rd_st2_638  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[638]), .rdlo_in(a2_wr[894]),  .coef_in(coef[504]), .rdup_out(a3_wr[638]), .rdlo_out(a3_wr[894]));
			radix2 #(.width(width)) rd_st2_639  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[639]), .rdlo_in(a2_wr[895]),  .coef_in(coef[508]), .rdup_out(a3_wr[639]), .rdlo_out(a3_wr[895]));
			radix2 #(.width(width)) rd_st2_640  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[640]), .rdlo_in(a2_wr[896]),  .coef_in(coef[512]), .rdup_out(a3_wr[640]), .rdlo_out(a3_wr[896]));
			radix2 #(.width(width)) rd_st2_641  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[641]), .rdlo_in(a2_wr[897]),  .coef_in(coef[516]), .rdup_out(a3_wr[641]), .rdlo_out(a3_wr[897]));
			radix2 #(.width(width)) rd_st2_642  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[642]), .rdlo_in(a2_wr[898]),  .coef_in(coef[520]), .rdup_out(a3_wr[642]), .rdlo_out(a3_wr[898]));
			radix2 #(.width(width)) rd_st2_643  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[643]), .rdlo_in(a2_wr[899]),  .coef_in(coef[524]), .rdup_out(a3_wr[643]), .rdlo_out(a3_wr[899]));
			radix2 #(.width(width)) rd_st2_644  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[644]), .rdlo_in(a2_wr[900]),  .coef_in(coef[528]), .rdup_out(a3_wr[644]), .rdlo_out(a3_wr[900]));
			radix2 #(.width(width)) rd_st2_645  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[645]), .rdlo_in(a2_wr[901]),  .coef_in(coef[532]), .rdup_out(a3_wr[645]), .rdlo_out(a3_wr[901]));
			radix2 #(.width(width)) rd_st2_646  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[646]), .rdlo_in(a2_wr[902]),  .coef_in(coef[536]), .rdup_out(a3_wr[646]), .rdlo_out(a3_wr[902]));
			radix2 #(.width(width)) rd_st2_647  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[647]), .rdlo_in(a2_wr[903]),  .coef_in(coef[540]), .rdup_out(a3_wr[647]), .rdlo_out(a3_wr[903]));
			radix2 #(.width(width)) rd_st2_648  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[648]), .rdlo_in(a2_wr[904]),  .coef_in(coef[544]), .rdup_out(a3_wr[648]), .rdlo_out(a3_wr[904]));
			radix2 #(.width(width)) rd_st2_649  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[649]), .rdlo_in(a2_wr[905]),  .coef_in(coef[548]), .rdup_out(a3_wr[649]), .rdlo_out(a3_wr[905]));
			radix2 #(.width(width)) rd_st2_650  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[650]), .rdlo_in(a2_wr[906]),  .coef_in(coef[552]), .rdup_out(a3_wr[650]), .rdlo_out(a3_wr[906]));
			radix2 #(.width(width)) rd_st2_651  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[651]), .rdlo_in(a2_wr[907]),  .coef_in(coef[556]), .rdup_out(a3_wr[651]), .rdlo_out(a3_wr[907]));
			radix2 #(.width(width)) rd_st2_652  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[652]), .rdlo_in(a2_wr[908]),  .coef_in(coef[560]), .rdup_out(a3_wr[652]), .rdlo_out(a3_wr[908]));
			radix2 #(.width(width)) rd_st2_653  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[653]), .rdlo_in(a2_wr[909]),  .coef_in(coef[564]), .rdup_out(a3_wr[653]), .rdlo_out(a3_wr[909]));
			radix2 #(.width(width)) rd_st2_654  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[654]), .rdlo_in(a2_wr[910]),  .coef_in(coef[568]), .rdup_out(a3_wr[654]), .rdlo_out(a3_wr[910]));
			radix2 #(.width(width)) rd_st2_655  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[655]), .rdlo_in(a2_wr[911]),  .coef_in(coef[572]), .rdup_out(a3_wr[655]), .rdlo_out(a3_wr[911]));
			radix2 #(.width(width)) rd_st2_656  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[656]), .rdlo_in(a2_wr[912]),  .coef_in(coef[576]), .rdup_out(a3_wr[656]), .rdlo_out(a3_wr[912]));
			radix2 #(.width(width)) rd_st2_657  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[657]), .rdlo_in(a2_wr[913]),  .coef_in(coef[580]), .rdup_out(a3_wr[657]), .rdlo_out(a3_wr[913]));
			radix2 #(.width(width)) rd_st2_658  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[658]), .rdlo_in(a2_wr[914]),  .coef_in(coef[584]), .rdup_out(a3_wr[658]), .rdlo_out(a3_wr[914]));
			radix2 #(.width(width)) rd_st2_659  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[659]), .rdlo_in(a2_wr[915]),  .coef_in(coef[588]), .rdup_out(a3_wr[659]), .rdlo_out(a3_wr[915]));
			radix2 #(.width(width)) rd_st2_660  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[660]), .rdlo_in(a2_wr[916]),  .coef_in(coef[592]), .rdup_out(a3_wr[660]), .rdlo_out(a3_wr[916]));
			radix2 #(.width(width)) rd_st2_661  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[661]), .rdlo_in(a2_wr[917]),  .coef_in(coef[596]), .rdup_out(a3_wr[661]), .rdlo_out(a3_wr[917]));
			radix2 #(.width(width)) rd_st2_662  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[662]), .rdlo_in(a2_wr[918]),  .coef_in(coef[600]), .rdup_out(a3_wr[662]), .rdlo_out(a3_wr[918]));
			radix2 #(.width(width)) rd_st2_663  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[663]), .rdlo_in(a2_wr[919]),  .coef_in(coef[604]), .rdup_out(a3_wr[663]), .rdlo_out(a3_wr[919]));
			radix2 #(.width(width)) rd_st2_664  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[664]), .rdlo_in(a2_wr[920]),  .coef_in(coef[608]), .rdup_out(a3_wr[664]), .rdlo_out(a3_wr[920]));
			radix2 #(.width(width)) rd_st2_665  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[665]), .rdlo_in(a2_wr[921]),  .coef_in(coef[612]), .rdup_out(a3_wr[665]), .rdlo_out(a3_wr[921]));
			radix2 #(.width(width)) rd_st2_666  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[666]), .rdlo_in(a2_wr[922]),  .coef_in(coef[616]), .rdup_out(a3_wr[666]), .rdlo_out(a3_wr[922]));
			radix2 #(.width(width)) rd_st2_667  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[667]), .rdlo_in(a2_wr[923]),  .coef_in(coef[620]), .rdup_out(a3_wr[667]), .rdlo_out(a3_wr[923]));
			radix2 #(.width(width)) rd_st2_668  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[668]), .rdlo_in(a2_wr[924]),  .coef_in(coef[624]), .rdup_out(a3_wr[668]), .rdlo_out(a3_wr[924]));
			radix2 #(.width(width)) rd_st2_669  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[669]), .rdlo_in(a2_wr[925]),  .coef_in(coef[628]), .rdup_out(a3_wr[669]), .rdlo_out(a3_wr[925]));
			radix2 #(.width(width)) rd_st2_670  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[670]), .rdlo_in(a2_wr[926]),  .coef_in(coef[632]), .rdup_out(a3_wr[670]), .rdlo_out(a3_wr[926]));
			radix2 #(.width(width)) rd_st2_671  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[671]), .rdlo_in(a2_wr[927]),  .coef_in(coef[636]), .rdup_out(a3_wr[671]), .rdlo_out(a3_wr[927]));
			radix2 #(.width(width)) rd_st2_672  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[672]), .rdlo_in(a2_wr[928]),  .coef_in(coef[640]), .rdup_out(a3_wr[672]), .rdlo_out(a3_wr[928]));
			radix2 #(.width(width)) rd_st2_673  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[673]), .rdlo_in(a2_wr[929]),  .coef_in(coef[644]), .rdup_out(a3_wr[673]), .rdlo_out(a3_wr[929]));
			radix2 #(.width(width)) rd_st2_674  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[674]), .rdlo_in(a2_wr[930]),  .coef_in(coef[648]), .rdup_out(a3_wr[674]), .rdlo_out(a3_wr[930]));
			radix2 #(.width(width)) rd_st2_675  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[675]), .rdlo_in(a2_wr[931]),  .coef_in(coef[652]), .rdup_out(a3_wr[675]), .rdlo_out(a3_wr[931]));
			radix2 #(.width(width)) rd_st2_676  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[676]), .rdlo_in(a2_wr[932]),  .coef_in(coef[656]), .rdup_out(a3_wr[676]), .rdlo_out(a3_wr[932]));
			radix2 #(.width(width)) rd_st2_677  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[677]), .rdlo_in(a2_wr[933]),  .coef_in(coef[660]), .rdup_out(a3_wr[677]), .rdlo_out(a3_wr[933]));
			radix2 #(.width(width)) rd_st2_678  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[678]), .rdlo_in(a2_wr[934]),  .coef_in(coef[664]), .rdup_out(a3_wr[678]), .rdlo_out(a3_wr[934]));
			radix2 #(.width(width)) rd_st2_679  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[679]), .rdlo_in(a2_wr[935]),  .coef_in(coef[668]), .rdup_out(a3_wr[679]), .rdlo_out(a3_wr[935]));
			radix2 #(.width(width)) rd_st2_680  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[680]), .rdlo_in(a2_wr[936]),  .coef_in(coef[672]), .rdup_out(a3_wr[680]), .rdlo_out(a3_wr[936]));
			radix2 #(.width(width)) rd_st2_681  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[681]), .rdlo_in(a2_wr[937]),  .coef_in(coef[676]), .rdup_out(a3_wr[681]), .rdlo_out(a3_wr[937]));
			radix2 #(.width(width)) rd_st2_682  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[682]), .rdlo_in(a2_wr[938]),  .coef_in(coef[680]), .rdup_out(a3_wr[682]), .rdlo_out(a3_wr[938]));
			radix2 #(.width(width)) rd_st2_683  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[683]), .rdlo_in(a2_wr[939]),  .coef_in(coef[684]), .rdup_out(a3_wr[683]), .rdlo_out(a3_wr[939]));
			radix2 #(.width(width)) rd_st2_684  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[684]), .rdlo_in(a2_wr[940]),  .coef_in(coef[688]), .rdup_out(a3_wr[684]), .rdlo_out(a3_wr[940]));
			radix2 #(.width(width)) rd_st2_685  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[685]), .rdlo_in(a2_wr[941]),  .coef_in(coef[692]), .rdup_out(a3_wr[685]), .rdlo_out(a3_wr[941]));
			radix2 #(.width(width)) rd_st2_686  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[686]), .rdlo_in(a2_wr[942]),  .coef_in(coef[696]), .rdup_out(a3_wr[686]), .rdlo_out(a3_wr[942]));
			radix2 #(.width(width)) rd_st2_687  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[687]), .rdlo_in(a2_wr[943]),  .coef_in(coef[700]), .rdup_out(a3_wr[687]), .rdlo_out(a3_wr[943]));
			radix2 #(.width(width)) rd_st2_688  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[688]), .rdlo_in(a2_wr[944]),  .coef_in(coef[704]), .rdup_out(a3_wr[688]), .rdlo_out(a3_wr[944]));
			radix2 #(.width(width)) rd_st2_689  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[689]), .rdlo_in(a2_wr[945]),  .coef_in(coef[708]), .rdup_out(a3_wr[689]), .rdlo_out(a3_wr[945]));
			radix2 #(.width(width)) rd_st2_690  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[690]), .rdlo_in(a2_wr[946]),  .coef_in(coef[712]), .rdup_out(a3_wr[690]), .rdlo_out(a3_wr[946]));
			radix2 #(.width(width)) rd_st2_691  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[691]), .rdlo_in(a2_wr[947]),  .coef_in(coef[716]), .rdup_out(a3_wr[691]), .rdlo_out(a3_wr[947]));
			radix2 #(.width(width)) rd_st2_692  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[692]), .rdlo_in(a2_wr[948]),  .coef_in(coef[720]), .rdup_out(a3_wr[692]), .rdlo_out(a3_wr[948]));
			radix2 #(.width(width)) rd_st2_693  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[693]), .rdlo_in(a2_wr[949]),  .coef_in(coef[724]), .rdup_out(a3_wr[693]), .rdlo_out(a3_wr[949]));
			radix2 #(.width(width)) rd_st2_694  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[694]), .rdlo_in(a2_wr[950]),  .coef_in(coef[728]), .rdup_out(a3_wr[694]), .rdlo_out(a3_wr[950]));
			radix2 #(.width(width)) rd_st2_695  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[695]), .rdlo_in(a2_wr[951]),  .coef_in(coef[732]), .rdup_out(a3_wr[695]), .rdlo_out(a3_wr[951]));
			radix2 #(.width(width)) rd_st2_696  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[696]), .rdlo_in(a2_wr[952]),  .coef_in(coef[736]), .rdup_out(a3_wr[696]), .rdlo_out(a3_wr[952]));
			radix2 #(.width(width)) rd_st2_697  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[697]), .rdlo_in(a2_wr[953]),  .coef_in(coef[740]), .rdup_out(a3_wr[697]), .rdlo_out(a3_wr[953]));
			radix2 #(.width(width)) rd_st2_698  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[698]), .rdlo_in(a2_wr[954]),  .coef_in(coef[744]), .rdup_out(a3_wr[698]), .rdlo_out(a3_wr[954]));
			radix2 #(.width(width)) rd_st2_699  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[699]), .rdlo_in(a2_wr[955]),  .coef_in(coef[748]), .rdup_out(a3_wr[699]), .rdlo_out(a3_wr[955]));
			radix2 #(.width(width)) rd_st2_700  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[700]), .rdlo_in(a2_wr[956]),  .coef_in(coef[752]), .rdup_out(a3_wr[700]), .rdlo_out(a3_wr[956]));
			radix2 #(.width(width)) rd_st2_701  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[701]), .rdlo_in(a2_wr[957]),  .coef_in(coef[756]), .rdup_out(a3_wr[701]), .rdlo_out(a3_wr[957]));
			radix2 #(.width(width)) rd_st2_702  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[702]), .rdlo_in(a2_wr[958]),  .coef_in(coef[760]), .rdup_out(a3_wr[702]), .rdlo_out(a3_wr[958]));
			radix2 #(.width(width)) rd_st2_703  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[703]), .rdlo_in(a2_wr[959]),  .coef_in(coef[764]), .rdup_out(a3_wr[703]), .rdlo_out(a3_wr[959]));
			radix2 #(.width(width)) rd_st2_704  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[704]), .rdlo_in(a2_wr[960]),  .coef_in(coef[768]), .rdup_out(a3_wr[704]), .rdlo_out(a3_wr[960]));
			radix2 #(.width(width)) rd_st2_705  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[705]), .rdlo_in(a2_wr[961]),  .coef_in(coef[772]), .rdup_out(a3_wr[705]), .rdlo_out(a3_wr[961]));
			radix2 #(.width(width)) rd_st2_706  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[706]), .rdlo_in(a2_wr[962]),  .coef_in(coef[776]), .rdup_out(a3_wr[706]), .rdlo_out(a3_wr[962]));
			radix2 #(.width(width)) rd_st2_707  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[707]), .rdlo_in(a2_wr[963]),  .coef_in(coef[780]), .rdup_out(a3_wr[707]), .rdlo_out(a3_wr[963]));
			radix2 #(.width(width)) rd_st2_708  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[708]), .rdlo_in(a2_wr[964]),  .coef_in(coef[784]), .rdup_out(a3_wr[708]), .rdlo_out(a3_wr[964]));
			radix2 #(.width(width)) rd_st2_709  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[709]), .rdlo_in(a2_wr[965]),  .coef_in(coef[788]), .rdup_out(a3_wr[709]), .rdlo_out(a3_wr[965]));
			radix2 #(.width(width)) rd_st2_710  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[710]), .rdlo_in(a2_wr[966]),  .coef_in(coef[792]), .rdup_out(a3_wr[710]), .rdlo_out(a3_wr[966]));
			radix2 #(.width(width)) rd_st2_711  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[711]), .rdlo_in(a2_wr[967]),  .coef_in(coef[796]), .rdup_out(a3_wr[711]), .rdlo_out(a3_wr[967]));
			radix2 #(.width(width)) rd_st2_712  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[712]), .rdlo_in(a2_wr[968]),  .coef_in(coef[800]), .rdup_out(a3_wr[712]), .rdlo_out(a3_wr[968]));
			radix2 #(.width(width)) rd_st2_713  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[713]), .rdlo_in(a2_wr[969]),  .coef_in(coef[804]), .rdup_out(a3_wr[713]), .rdlo_out(a3_wr[969]));
			radix2 #(.width(width)) rd_st2_714  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[714]), .rdlo_in(a2_wr[970]),  .coef_in(coef[808]), .rdup_out(a3_wr[714]), .rdlo_out(a3_wr[970]));
			radix2 #(.width(width)) rd_st2_715  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[715]), .rdlo_in(a2_wr[971]),  .coef_in(coef[812]), .rdup_out(a3_wr[715]), .rdlo_out(a3_wr[971]));
			radix2 #(.width(width)) rd_st2_716  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[716]), .rdlo_in(a2_wr[972]),  .coef_in(coef[816]), .rdup_out(a3_wr[716]), .rdlo_out(a3_wr[972]));
			radix2 #(.width(width)) rd_st2_717  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[717]), .rdlo_in(a2_wr[973]),  .coef_in(coef[820]), .rdup_out(a3_wr[717]), .rdlo_out(a3_wr[973]));
			radix2 #(.width(width)) rd_st2_718  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[718]), .rdlo_in(a2_wr[974]),  .coef_in(coef[824]), .rdup_out(a3_wr[718]), .rdlo_out(a3_wr[974]));
			radix2 #(.width(width)) rd_st2_719  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[719]), .rdlo_in(a2_wr[975]),  .coef_in(coef[828]), .rdup_out(a3_wr[719]), .rdlo_out(a3_wr[975]));
			radix2 #(.width(width)) rd_st2_720  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[720]), .rdlo_in(a2_wr[976]),  .coef_in(coef[832]), .rdup_out(a3_wr[720]), .rdlo_out(a3_wr[976]));
			radix2 #(.width(width)) rd_st2_721  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[721]), .rdlo_in(a2_wr[977]),  .coef_in(coef[836]), .rdup_out(a3_wr[721]), .rdlo_out(a3_wr[977]));
			radix2 #(.width(width)) rd_st2_722  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[722]), .rdlo_in(a2_wr[978]),  .coef_in(coef[840]), .rdup_out(a3_wr[722]), .rdlo_out(a3_wr[978]));
			radix2 #(.width(width)) rd_st2_723  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[723]), .rdlo_in(a2_wr[979]),  .coef_in(coef[844]), .rdup_out(a3_wr[723]), .rdlo_out(a3_wr[979]));
			radix2 #(.width(width)) rd_st2_724  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[724]), .rdlo_in(a2_wr[980]),  .coef_in(coef[848]), .rdup_out(a3_wr[724]), .rdlo_out(a3_wr[980]));
			radix2 #(.width(width)) rd_st2_725  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[725]), .rdlo_in(a2_wr[981]),  .coef_in(coef[852]), .rdup_out(a3_wr[725]), .rdlo_out(a3_wr[981]));
			radix2 #(.width(width)) rd_st2_726  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[726]), .rdlo_in(a2_wr[982]),  .coef_in(coef[856]), .rdup_out(a3_wr[726]), .rdlo_out(a3_wr[982]));
			radix2 #(.width(width)) rd_st2_727  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[727]), .rdlo_in(a2_wr[983]),  .coef_in(coef[860]), .rdup_out(a3_wr[727]), .rdlo_out(a3_wr[983]));
			radix2 #(.width(width)) rd_st2_728  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[728]), .rdlo_in(a2_wr[984]),  .coef_in(coef[864]), .rdup_out(a3_wr[728]), .rdlo_out(a3_wr[984]));
			radix2 #(.width(width)) rd_st2_729  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[729]), .rdlo_in(a2_wr[985]),  .coef_in(coef[868]), .rdup_out(a3_wr[729]), .rdlo_out(a3_wr[985]));
			radix2 #(.width(width)) rd_st2_730  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[730]), .rdlo_in(a2_wr[986]),  .coef_in(coef[872]), .rdup_out(a3_wr[730]), .rdlo_out(a3_wr[986]));
			radix2 #(.width(width)) rd_st2_731  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[731]), .rdlo_in(a2_wr[987]),  .coef_in(coef[876]), .rdup_out(a3_wr[731]), .rdlo_out(a3_wr[987]));
			radix2 #(.width(width)) rd_st2_732  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[732]), .rdlo_in(a2_wr[988]),  .coef_in(coef[880]), .rdup_out(a3_wr[732]), .rdlo_out(a3_wr[988]));
			radix2 #(.width(width)) rd_st2_733  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[733]), .rdlo_in(a2_wr[989]),  .coef_in(coef[884]), .rdup_out(a3_wr[733]), .rdlo_out(a3_wr[989]));
			radix2 #(.width(width)) rd_st2_734  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[734]), .rdlo_in(a2_wr[990]),  .coef_in(coef[888]), .rdup_out(a3_wr[734]), .rdlo_out(a3_wr[990]));
			radix2 #(.width(width)) rd_st2_735  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[735]), .rdlo_in(a2_wr[991]),  .coef_in(coef[892]), .rdup_out(a3_wr[735]), .rdlo_out(a3_wr[991]));
			radix2 #(.width(width)) rd_st2_736  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[736]), .rdlo_in(a2_wr[992]),  .coef_in(coef[896]), .rdup_out(a3_wr[736]), .rdlo_out(a3_wr[992]));
			radix2 #(.width(width)) rd_st2_737  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[737]), .rdlo_in(a2_wr[993]),  .coef_in(coef[900]), .rdup_out(a3_wr[737]), .rdlo_out(a3_wr[993]));
			radix2 #(.width(width)) rd_st2_738  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[738]), .rdlo_in(a2_wr[994]),  .coef_in(coef[904]), .rdup_out(a3_wr[738]), .rdlo_out(a3_wr[994]));
			radix2 #(.width(width)) rd_st2_739  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[739]), .rdlo_in(a2_wr[995]),  .coef_in(coef[908]), .rdup_out(a3_wr[739]), .rdlo_out(a3_wr[995]));
			radix2 #(.width(width)) rd_st2_740  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[740]), .rdlo_in(a2_wr[996]),  .coef_in(coef[912]), .rdup_out(a3_wr[740]), .rdlo_out(a3_wr[996]));
			radix2 #(.width(width)) rd_st2_741  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[741]), .rdlo_in(a2_wr[997]),  .coef_in(coef[916]), .rdup_out(a3_wr[741]), .rdlo_out(a3_wr[997]));
			radix2 #(.width(width)) rd_st2_742  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[742]), .rdlo_in(a2_wr[998]),  .coef_in(coef[920]), .rdup_out(a3_wr[742]), .rdlo_out(a3_wr[998]));
			radix2 #(.width(width)) rd_st2_743  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[743]), .rdlo_in(a2_wr[999]),  .coef_in(coef[924]), .rdup_out(a3_wr[743]), .rdlo_out(a3_wr[999]));
			radix2 #(.width(width)) rd_st2_744  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[744]), .rdlo_in(a2_wr[1000]),  .coef_in(coef[928]), .rdup_out(a3_wr[744]), .rdlo_out(a3_wr[1000]));
			radix2 #(.width(width)) rd_st2_745  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[745]), .rdlo_in(a2_wr[1001]),  .coef_in(coef[932]), .rdup_out(a3_wr[745]), .rdlo_out(a3_wr[1001]));
			radix2 #(.width(width)) rd_st2_746  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[746]), .rdlo_in(a2_wr[1002]),  .coef_in(coef[936]), .rdup_out(a3_wr[746]), .rdlo_out(a3_wr[1002]));
			radix2 #(.width(width)) rd_st2_747  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[747]), .rdlo_in(a2_wr[1003]),  .coef_in(coef[940]), .rdup_out(a3_wr[747]), .rdlo_out(a3_wr[1003]));
			radix2 #(.width(width)) rd_st2_748  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[748]), .rdlo_in(a2_wr[1004]),  .coef_in(coef[944]), .rdup_out(a3_wr[748]), .rdlo_out(a3_wr[1004]));
			radix2 #(.width(width)) rd_st2_749  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[749]), .rdlo_in(a2_wr[1005]),  .coef_in(coef[948]), .rdup_out(a3_wr[749]), .rdlo_out(a3_wr[1005]));
			radix2 #(.width(width)) rd_st2_750  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[750]), .rdlo_in(a2_wr[1006]),  .coef_in(coef[952]), .rdup_out(a3_wr[750]), .rdlo_out(a3_wr[1006]));
			radix2 #(.width(width)) rd_st2_751  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[751]), .rdlo_in(a2_wr[1007]),  .coef_in(coef[956]), .rdup_out(a3_wr[751]), .rdlo_out(a3_wr[1007]));
			radix2 #(.width(width)) rd_st2_752  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[752]), .rdlo_in(a2_wr[1008]),  .coef_in(coef[960]), .rdup_out(a3_wr[752]), .rdlo_out(a3_wr[1008]));
			radix2 #(.width(width)) rd_st2_753  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[753]), .rdlo_in(a2_wr[1009]),  .coef_in(coef[964]), .rdup_out(a3_wr[753]), .rdlo_out(a3_wr[1009]));
			radix2 #(.width(width)) rd_st2_754  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[754]), .rdlo_in(a2_wr[1010]),  .coef_in(coef[968]), .rdup_out(a3_wr[754]), .rdlo_out(a3_wr[1010]));
			radix2 #(.width(width)) rd_st2_755  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[755]), .rdlo_in(a2_wr[1011]),  .coef_in(coef[972]), .rdup_out(a3_wr[755]), .rdlo_out(a3_wr[1011]));
			radix2 #(.width(width)) rd_st2_756  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[756]), .rdlo_in(a2_wr[1012]),  .coef_in(coef[976]), .rdup_out(a3_wr[756]), .rdlo_out(a3_wr[1012]));
			radix2 #(.width(width)) rd_st2_757  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[757]), .rdlo_in(a2_wr[1013]),  .coef_in(coef[980]), .rdup_out(a3_wr[757]), .rdlo_out(a3_wr[1013]));
			radix2 #(.width(width)) rd_st2_758  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[758]), .rdlo_in(a2_wr[1014]),  .coef_in(coef[984]), .rdup_out(a3_wr[758]), .rdlo_out(a3_wr[1014]));
			radix2 #(.width(width)) rd_st2_759  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[759]), .rdlo_in(a2_wr[1015]),  .coef_in(coef[988]), .rdup_out(a3_wr[759]), .rdlo_out(a3_wr[1015]));
			radix2 #(.width(width)) rd_st2_760  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[760]), .rdlo_in(a2_wr[1016]),  .coef_in(coef[992]), .rdup_out(a3_wr[760]), .rdlo_out(a3_wr[1016]));
			radix2 #(.width(width)) rd_st2_761  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[761]), .rdlo_in(a2_wr[1017]),  .coef_in(coef[996]), .rdup_out(a3_wr[761]), .rdlo_out(a3_wr[1017]));
			radix2 #(.width(width)) rd_st2_762  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[762]), .rdlo_in(a2_wr[1018]),  .coef_in(coef[1000]), .rdup_out(a3_wr[762]), .rdlo_out(a3_wr[1018]));
			radix2 #(.width(width)) rd_st2_763  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[763]), .rdlo_in(a2_wr[1019]),  .coef_in(coef[1004]), .rdup_out(a3_wr[763]), .rdlo_out(a3_wr[1019]));
			radix2 #(.width(width)) rd_st2_764  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[764]), .rdlo_in(a2_wr[1020]),  .coef_in(coef[1008]), .rdup_out(a3_wr[764]), .rdlo_out(a3_wr[1020]));
			radix2 #(.width(width)) rd_st2_765  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[765]), .rdlo_in(a2_wr[1021]),  .coef_in(coef[1012]), .rdup_out(a3_wr[765]), .rdlo_out(a3_wr[1021]));
			radix2 #(.width(width)) rd_st2_766  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[766]), .rdlo_in(a2_wr[1022]),  .coef_in(coef[1016]), .rdup_out(a3_wr[766]), .rdlo_out(a3_wr[1022]));
			radix2 #(.width(width)) rd_st2_767  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[767]), .rdlo_in(a2_wr[1023]),  .coef_in(coef[1020]), .rdup_out(a3_wr[767]), .rdlo_out(a3_wr[1023]));
			radix2 #(.width(width)) rd_st2_1024  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1024]), .rdlo_in(a2_wr[1280]),  .coef_in(coef[0]), .rdup_out(a3_wr[1024]), .rdlo_out(a3_wr[1280]));
			radix2 #(.width(width)) rd_st2_1025  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1025]), .rdlo_in(a2_wr[1281]),  .coef_in(coef[4]), .rdup_out(a3_wr[1025]), .rdlo_out(a3_wr[1281]));
			radix2 #(.width(width)) rd_st2_1026  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1026]), .rdlo_in(a2_wr[1282]),  .coef_in(coef[8]), .rdup_out(a3_wr[1026]), .rdlo_out(a3_wr[1282]));
			radix2 #(.width(width)) rd_st2_1027  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1027]), .rdlo_in(a2_wr[1283]),  .coef_in(coef[12]), .rdup_out(a3_wr[1027]), .rdlo_out(a3_wr[1283]));
			radix2 #(.width(width)) rd_st2_1028  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1028]), .rdlo_in(a2_wr[1284]),  .coef_in(coef[16]), .rdup_out(a3_wr[1028]), .rdlo_out(a3_wr[1284]));
			radix2 #(.width(width)) rd_st2_1029  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1029]), .rdlo_in(a2_wr[1285]),  .coef_in(coef[20]), .rdup_out(a3_wr[1029]), .rdlo_out(a3_wr[1285]));
			radix2 #(.width(width)) rd_st2_1030  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1030]), .rdlo_in(a2_wr[1286]),  .coef_in(coef[24]), .rdup_out(a3_wr[1030]), .rdlo_out(a3_wr[1286]));
			radix2 #(.width(width)) rd_st2_1031  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1031]), .rdlo_in(a2_wr[1287]),  .coef_in(coef[28]), .rdup_out(a3_wr[1031]), .rdlo_out(a3_wr[1287]));
			radix2 #(.width(width)) rd_st2_1032  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1032]), .rdlo_in(a2_wr[1288]),  .coef_in(coef[32]), .rdup_out(a3_wr[1032]), .rdlo_out(a3_wr[1288]));
			radix2 #(.width(width)) rd_st2_1033  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1033]), .rdlo_in(a2_wr[1289]),  .coef_in(coef[36]), .rdup_out(a3_wr[1033]), .rdlo_out(a3_wr[1289]));
			radix2 #(.width(width)) rd_st2_1034  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1034]), .rdlo_in(a2_wr[1290]),  .coef_in(coef[40]), .rdup_out(a3_wr[1034]), .rdlo_out(a3_wr[1290]));
			radix2 #(.width(width)) rd_st2_1035  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1035]), .rdlo_in(a2_wr[1291]),  .coef_in(coef[44]), .rdup_out(a3_wr[1035]), .rdlo_out(a3_wr[1291]));
			radix2 #(.width(width)) rd_st2_1036  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1036]), .rdlo_in(a2_wr[1292]),  .coef_in(coef[48]), .rdup_out(a3_wr[1036]), .rdlo_out(a3_wr[1292]));
			radix2 #(.width(width)) rd_st2_1037  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1037]), .rdlo_in(a2_wr[1293]),  .coef_in(coef[52]), .rdup_out(a3_wr[1037]), .rdlo_out(a3_wr[1293]));
			radix2 #(.width(width)) rd_st2_1038  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1038]), .rdlo_in(a2_wr[1294]),  .coef_in(coef[56]), .rdup_out(a3_wr[1038]), .rdlo_out(a3_wr[1294]));
			radix2 #(.width(width)) rd_st2_1039  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1039]), .rdlo_in(a2_wr[1295]),  .coef_in(coef[60]), .rdup_out(a3_wr[1039]), .rdlo_out(a3_wr[1295]));
			radix2 #(.width(width)) rd_st2_1040  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1040]), .rdlo_in(a2_wr[1296]),  .coef_in(coef[64]), .rdup_out(a3_wr[1040]), .rdlo_out(a3_wr[1296]));
			radix2 #(.width(width)) rd_st2_1041  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1041]), .rdlo_in(a2_wr[1297]),  .coef_in(coef[68]), .rdup_out(a3_wr[1041]), .rdlo_out(a3_wr[1297]));
			radix2 #(.width(width)) rd_st2_1042  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1042]), .rdlo_in(a2_wr[1298]),  .coef_in(coef[72]), .rdup_out(a3_wr[1042]), .rdlo_out(a3_wr[1298]));
			radix2 #(.width(width)) rd_st2_1043  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1043]), .rdlo_in(a2_wr[1299]),  .coef_in(coef[76]), .rdup_out(a3_wr[1043]), .rdlo_out(a3_wr[1299]));
			radix2 #(.width(width)) rd_st2_1044  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1044]), .rdlo_in(a2_wr[1300]),  .coef_in(coef[80]), .rdup_out(a3_wr[1044]), .rdlo_out(a3_wr[1300]));
			radix2 #(.width(width)) rd_st2_1045  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1045]), .rdlo_in(a2_wr[1301]),  .coef_in(coef[84]), .rdup_out(a3_wr[1045]), .rdlo_out(a3_wr[1301]));
			radix2 #(.width(width)) rd_st2_1046  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1046]), .rdlo_in(a2_wr[1302]),  .coef_in(coef[88]), .rdup_out(a3_wr[1046]), .rdlo_out(a3_wr[1302]));
			radix2 #(.width(width)) rd_st2_1047  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1047]), .rdlo_in(a2_wr[1303]),  .coef_in(coef[92]), .rdup_out(a3_wr[1047]), .rdlo_out(a3_wr[1303]));
			radix2 #(.width(width)) rd_st2_1048  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1048]), .rdlo_in(a2_wr[1304]),  .coef_in(coef[96]), .rdup_out(a3_wr[1048]), .rdlo_out(a3_wr[1304]));
			radix2 #(.width(width)) rd_st2_1049  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1049]), .rdlo_in(a2_wr[1305]),  .coef_in(coef[100]), .rdup_out(a3_wr[1049]), .rdlo_out(a3_wr[1305]));
			radix2 #(.width(width)) rd_st2_1050  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1050]), .rdlo_in(a2_wr[1306]),  .coef_in(coef[104]), .rdup_out(a3_wr[1050]), .rdlo_out(a3_wr[1306]));
			radix2 #(.width(width)) rd_st2_1051  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1051]), .rdlo_in(a2_wr[1307]),  .coef_in(coef[108]), .rdup_out(a3_wr[1051]), .rdlo_out(a3_wr[1307]));
			radix2 #(.width(width)) rd_st2_1052  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1052]), .rdlo_in(a2_wr[1308]),  .coef_in(coef[112]), .rdup_out(a3_wr[1052]), .rdlo_out(a3_wr[1308]));
			radix2 #(.width(width)) rd_st2_1053  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1053]), .rdlo_in(a2_wr[1309]),  .coef_in(coef[116]), .rdup_out(a3_wr[1053]), .rdlo_out(a3_wr[1309]));
			radix2 #(.width(width)) rd_st2_1054  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1054]), .rdlo_in(a2_wr[1310]),  .coef_in(coef[120]), .rdup_out(a3_wr[1054]), .rdlo_out(a3_wr[1310]));
			radix2 #(.width(width)) rd_st2_1055  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1055]), .rdlo_in(a2_wr[1311]),  .coef_in(coef[124]), .rdup_out(a3_wr[1055]), .rdlo_out(a3_wr[1311]));
			radix2 #(.width(width)) rd_st2_1056  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1056]), .rdlo_in(a2_wr[1312]),  .coef_in(coef[128]), .rdup_out(a3_wr[1056]), .rdlo_out(a3_wr[1312]));
			radix2 #(.width(width)) rd_st2_1057  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1057]), .rdlo_in(a2_wr[1313]),  .coef_in(coef[132]), .rdup_out(a3_wr[1057]), .rdlo_out(a3_wr[1313]));
			radix2 #(.width(width)) rd_st2_1058  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1058]), .rdlo_in(a2_wr[1314]),  .coef_in(coef[136]), .rdup_out(a3_wr[1058]), .rdlo_out(a3_wr[1314]));
			radix2 #(.width(width)) rd_st2_1059  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1059]), .rdlo_in(a2_wr[1315]),  .coef_in(coef[140]), .rdup_out(a3_wr[1059]), .rdlo_out(a3_wr[1315]));
			radix2 #(.width(width)) rd_st2_1060  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1060]), .rdlo_in(a2_wr[1316]),  .coef_in(coef[144]), .rdup_out(a3_wr[1060]), .rdlo_out(a3_wr[1316]));
			radix2 #(.width(width)) rd_st2_1061  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1061]), .rdlo_in(a2_wr[1317]),  .coef_in(coef[148]), .rdup_out(a3_wr[1061]), .rdlo_out(a3_wr[1317]));
			radix2 #(.width(width)) rd_st2_1062  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1062]), .rdlo_in(a2_wr[1318]),  .coef_in(coef[152]), .rdup_out(a3_wr[1062]), .rdlo_out(a3_wr[1318]));
			radix2 #(.width(width)) rd_st2_1063  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1063]), .rdlo_in(a2_wr[1319]),  .coef_in(coef[156]), .rdup_out(a3_wr[1063]), .rdlo_out(a3_wr[1319]));
			radix2 #(.width(width)) rd_st2_1064  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1064]), .rdlo_in(a2_wr[1320]),  .coef_in(coef[160]), .rdup_out(a3_wr[1064]), .rdlo_out(a3_wr[1320]));
			radix2 #(.width(width)) rd_st2_1065  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1065]), .rdlo_in(a2_wr[1321]),  .coef_in(coef[164]), .rdup_out(a3_wr[1065]), .rdlo_out(a3_wr[1321]));
			radix2 #(.width(width)) rd_st2_1066  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1066]), .rdlo_in(a2_wr[1322]),  .coef_in(coef[168]), .rdup_out(a3_wr[1066]), .rdlo_out(a3_wr[1322]));
			radix2 #(.width(width)) rd_st2_1067  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1067]), .rdlo_in(a2_wr[1323]),  .coef_in(coef[172]), .rdup_out(a3_wr[1067]), .rdlo_out(a3_wr[1323]));
			radix2 #(.width(width)) rd_st2_1068  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1068]), .rdlo_in(a2_wr[1324]),  .coef_in(coef[176]), .rdup_out(a3_wr[1068]), .rdlo_out(a3_wr[1324]));
			radix2 #(.width(width)) rd_st2_1069  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1069]), .rdlo_in(a2_wr[1325]),  .coef_in(coef[180]), .rdup_out(a3_wr[1069]), .rdlo_out(a3_wr[1325]));
			radix2 #(.width(width)) rd_st2_1070  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1070]), .rdlo_in(a2_wr[1326]),  .coef_in(coef[184]), .rdup_out(a3_wr[1070]), .rdlo_out(a3_wr[1326]));
			radix2 #(.width(width)) rd_st2_1071  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1071]), .rdlo_in(a2_wr[1327]),  .coef_in(coef[188]), .rdup_out(a3_wr[1071]), .rdlo_out(a3_wr[1327]));
			radix2 #(.width(width)) rd_st2_1072  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1072]), .rdlo_in(a2_wr[1328]),  .coef_in(coef[192]), .rdup_out(a3_wr[1072]), .rdlo_out(a3_wr[1328]));
			radix2 #(.width(width)) rd_st2_1073  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1073]), .rdlo_in(a2_wr[1329]),  .coef_in(coef[196]), .rdup_out(a3_wr[1073]), .rdlo_out(a3_wr[1329]));
			radix2 #(.width(width)) rd_st2_1074  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1074]), .rdlo_in(a2_wr[1330]),  .coef_in(coef[200]), .rdup_out(a3_wr[1074]), .rdlo_out(a3_wr[1330]));
			radix2 #(.width(width)) rd_st2_1075  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1075]), .rdlo_in(a2_wr[1331]),  .coef_in(coef[204]), .rdup_out(a3_wr[1075]), .rdlo_out(a3_wr[1331]));
			radix2 #(.width(width)) rd_st2_1076  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1076]), .rdlo_in(a2_wr[1332]),  .coef_in(coef[208]), .rdup_out(a3_wr[1076]), .rdlo_out(a3_wr[1332]));
			radix2 #(.width(width)) rd_st2_1077  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1077]), .rdlo_in(a2_wr[1333]),  .coef_in(coef[212]), .rdup_out(a3_wr[1077]), .rdlo_out(a3_wr[1333]));
			radix2 #(.width(width)) rd_st2_1078  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1078]), .rdlo_in(a2_wr[1334]),  .coef_in(coef[216]), .rdup_out(a3_wr[1078]), .rdlo_out(a3_wr[1334]));
			radix2 #(.width(width)) rd_st2_1079  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1079]), .rdlo_in(a2_wr[1335]),  .coef_in(coef[220]), .rdup_out(a3_wr[1079]), .rdlo_out(a3_wr[1335]));
			radix2 #(.width(width)) rd_st2_1080  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1080]), .rdlo_in(a2_wr[1336]),  .coef_in(coef[224]), .rdup_out(a3_wr[1080]), .rdlo_out(a3_wr[1336]));
			radix2 #(.width(width)) rd_st2_1081  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1081]), .rdlo_in(a2_wr[1337]),  .coef_in(coef[228]), .rdup_out(a3_wr[1081]), .rdlo_out(a3_wr[1337]));
			radix2 #(.width(width)) rd_st2_1082  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1082]), .rdlo_in(a2_wr[1338]),  .coef_in(coef[232]), .rdup_out(a3_wr[1082]), .rdlo_out(a3_wr[1338]));
			radix2 #(.width(width)) rd_st2_1083  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1083]), .rdlo_in(a2_wr[1339]),  .coef_in(coef[236]), .rdup_out(a3_wr[1083]), .rdlo_out(a3_wr[1339]));
			radix2 #(.width(width)) rd_st2_1084  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1084]), .rdlo_in(a2_wr[1340]),  .coef_in(coef[240]), .rdup_out(a3_wr[1084]), .rdlo_out(a3_wr[1340]));
			radix2 #(.width(width)) rd_st2_1085  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1085]), .rdlo_in(a2_wr[1341]),  .coef_in(coef[244]), .rdup_out(a3_wr[1085]), .rdlo_out(a3_wr[1341]));
			radix2 #(.width(width)) rd_st2_1086  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1086]), .rdlo_in(a2_wr[1342]),  .coef_in(coef[248]), .rdup_out(a3_wr[1086]), .rdlo_out(a3_wr[1342]));
			radix2 #(.width(width)) rd_st2_1087  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1087]), .rdlo_in(a2_wr[1343]),  .coef_in(coef[252]), .rdup_out(a3_wr[1087]), .rdlo_out(a3_wr[1343]));
			radix2 #(.width(width)) rd_st2_1088  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1088]), .rdlo_in(a2_wr[1344]),  .coef_in(coef[256]), .rdup_out(a3_wr[1088]), .rdlo_out(a3_wr[1344]));
			radix2 #(.width(width)) rd_st2_1089  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1089]), .rdlo_in(a2_wr[1345]),  .coef_in(coef[260]), .rdup_out(a3_wr[1089]), .rdlo_out(a3_wr[1345]));
			radix2 #(.width(width)) rd_st2_1090  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1090]), .rdlo_in(a2_wr[1346]),  .coef_in(coef[264]), .rdup_out(a3_wr[1090]), .rdlo_out(a3_wr[1346]));
			radix2 #(.width(width)) rd_st2_1091  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1091]), .rdlo_in(a2_wr[1347]),  .coef_in(coef[268]), .rdup_out(a3_wr[1091]), .rdlo_out(a3_wr[1347]));
			radix2 #(.width(width)) rd_st2_1092  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1092]), .rdlo_in(a2_wr[1348]),  .coef_in(coef[272]), .rdup_out(a3_wr[1092]), .rdlo_out(a3_wr[1348]));
			radix2 #(.width(width)) rd_st2_1093  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1093]), .rdlo_in(a2_wr[1349]),  .coef_in(coef[276]), .rdup_out(a3_wr[1093]), .rdlo_out(a3_wr[1349]));
			radix2 #(.width(width)) rd_st2_1094  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1094]), .rdlo_in(a2_wr[1350]),  .coef_in(coef[280]), .rdup_out(a3_wr[1094]), .rdlo_out(a3_wr[1350]));
			radix2 #(.width(width)) rd_st2_1095  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1095]), .rdlo_in(a2_wr[1351]),  .coef_in(coef[284]), .rdup_out(a3_wr[1095]), .rdlo_out(a3_wr[1351]));
			radix2 #(.width(width)) rd_st2_1096  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1096]), .rdlo_in(a2_wr[1352]),  .coef_in(coef[288]), .rdup_out(a3_wr[1096]), .rdlo_out(a3_wr[1352]));
			radix2 #(.width(width)) rd_st2_1097  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1097]), .rdlo_in(a2_wr[1353]),  .coef_in(coef[292]), .rdup_out(a3_wr[1097]), .rdlo_out(a3_wr[1353]));
			radix2 #(.width(width)) rd_st2_1098  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1098]), .rdlo_in(a2_wr[1354]),  .coef_in(coef[296]), .rdup_out(a3_wr[1098]), .rdlo_out(a3_wr[1354]));
			radix2 #(.width(width)) rd_st2_1099  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1099]), .rdlo_in(a2_wr[1355]),  .coef_in(coef[300]), .rdup_out(a3_wr[1099]), .rdlo_out(a3_wr[1355]));
			radix2 #(.width(width)) rd_st2_1100  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1100]), .rdlo_in(a2_wr[1356]),  .coef_in(coef[304]), .rdup_out(a3_wr[1100]), .rdlo_out(a3_wr[1356]));
			radix2 #(.width(width)) rd_st2_1101  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1101]), .rdlo_in(a2_wr[1357]),  .coef_in(coef[308]), .rdup_out(a3_wr[1101]), .rdlo_out(a3_wr[1357]));
			radix2 #(.width(width)) rd_st2_1102  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1102]), .rdlo_in(a2_wr[1358]),  .coef_in(coef[312]), .rdup_out(a3_wr[1102]), .rdlo_out(a3_wr[1358]));
			radix2 #(.width(width)) rd_st2_1103  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1103]), .rdlo_in(a2_wr[1359]),  .coef_in(coef[316]), .rdup_out(a3_wr[1103]), .rdlo_out(a3_wr[1359]));
			radix2 #(.width(width)) rd_st2_1104  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1104]), .rdlo_in(a2_wr[1360]),  .coef_in(coef[320]), .rdup_out(a3_wr[1104]), .rdlo_out(a3_wr[1360]));
			radix2 #(.width(width)) rd_st2_1105  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1105]), .rdlo_in(a2_wr[1361]),  .coef_in(coef[324]), .rdup_out(a3_wr[1105]), .rdlo_out(a3_wr[1361]));
			radix2 #(.width(width)) rd_st2_1106  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1106]), .rdlo_in(a2_wr[1362]),  .coef_in(coef[328]), .rdup_out(a3_wr[1106]), .rdlo_out(a3_wr[1362]));
			radix2 #(.width(width)) rd_st2_1107  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1107]), .rdlo_in(a2_wr[1363]),  .coef_in(coef[332]), .rdup_out(a3_wr[1107]), .rdlo_out(a3_wr[1363]));
			radix2 #(.width(width)) rd_st2_1108  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1108]), .rdlo_in(a2_wr[1364]),  .coef_in(coef[336]), .rdup_out(a3_wr[1108]), .rdlo_out(a3_wr[1364]));
			radix2 #(.width(width)) rd_st2_1109  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1109]), .rdlo_in(a2_wr[1365]),  .coef_in(coef[340]), .rdup_out(a3_wr[1109]), .rdlo_out(a3_wr[1365]));
			radix2 #(.width(width)) rd_st2_1110  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1110]), .rdlo_in(a2_wr[1366]),  .coef_in(coef[344]), .rdup_out(a3_wr[1110]), .rdlo_out(a3_wr[1366]));
			radix2 #(.width(width)) rd_st2_1111  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1111]), .rdlo_in(a2_wr[1367]),  .coef_in(coef[348]), .rdup_out(a3_wr[1111]), .rdlo_out(a3_wr[1367]));
			radix2 #(.width(width)) rd_st2_1112  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1112]), .rdlo_in(a2_wr[1368]),  .coef_in(coef[352]), .rdup_out(a3_wr[1112]), .rdlo_out(a3_wr[1368]));
			radix2 #(.width(width)) rd_st2_1113  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1113]), .rdlo_in(a2_wr[1369]),  .coef_in(coef[356]), .rdup_out(a3_wr[1113]), .rdlo_out(a3_wr[1369]));
			radix2 #(.width(width)) rd_st2_1114  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1114]), .rdlo_in(a2_wr[1370]),  .coef_in(coef[360]), .rdup_out(a3_wr[1114]), .rdlo_out(a3_wr[1370]));
			radix2 #(.width(width)) rd_st2_1115  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1115]), .rdlo_in(a2_wr[1371]),  .coef_in(coef[364]), .rdup_out(a3_wr[1115]), .rdlo_out(a3_wr[1371]));
			radix2 #(.width(width)) rd_st2_1116  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1116]), .rdlo_in(a2_wr[1372]),  .coef_in(coef[368]), .rdup_out(a3_wr[1116]), .rdlo_out(a3_wr[1372]));
			radix2 #(.width(width)) rd_st2_1117  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1117]), .rdlo_in(a2_wr[1373]),  .coef_in(coef[372]), .rdup_out(a3_wr[1117]), .rdlo_out(a3_wr[1373]));
			radix2 #(.width(width)) rd_st2_1118  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1118]), .rdlo_in(a2_wr[1374]),  .coef_in(coef[376]), .rdup_out(a3_wr[1118]), .rdlo_out(a3_wr[1374]));
			radix2 #(.width(width)) rd_st2_1119  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1119]), .rdlo_in(a2_wr[1375]),  .coef_in(coef[380]), .rdup_out(a3_wr[1119]), .rdlo_out(a3_wr[1375]));
			radix2 #(.width(width)) rd_st2_1120  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1120]), .rdlo_in(a2_wr[1376]),  .coef_in(coef[384]), .rdup_out(a3_wr[1120]), .rdlo_out(a3_wr[1376]));
			radix2 #(.width(width)) rd_st2_1121  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1121]), .rdlo_in(a2_wr[1377]),  .coef_in(coef[388]), .rdup_out(a3_wr[1121]), .rdlo_out(a3_wr[1377]));
			radix2 #(.width(width)) rd_st2_1122  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1122]), .rdlo_in(a2_wr[1378]),  .coef_in(coef[392]), .rdup_out(a3_wr[1122]), .rdlo_out(a3_wr[1378]));
			radix2 #(.width(width)) rd_st2_1123  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1123]), .rdlo_in(a2_wr[1379]),  .coef_in(coef[396]), .rdup_out(a3_wr[1123]), .rdlo_out(a3_wr[1379]));
			radix2 #(.width(width)) rd_st2_1124  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1124]), .rdlo_in(a2_wr[1380]),  .coef_in(coef[400]), .rdup_out(a3_wr[1124]), .rdlo_out(a3_wr[1380]));
			radix2 #(.width(width)) rd_st2_1125  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1125]), .rdlo_in(a2_wr[1381]),  .coef_in(coef[404]), .rdup_out(a3_wr[1125]), .rdlo_out(a3_wr[1381]));
			radix2 #(.width(width)) rd_st2_1126  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1126]), .rdlo_in(a2_wr[1382]),  .coef_in(coef[408]), .rdup_out(a3_wr[1126]), .rdlo_out(a3_wr[1382]));
			radix2 #(.width(width)) rd_st2_1127  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1127]), .rdlo_in(a2_wr[1383]),  .coef_in(coef[412]), .rdup_out(a3_wr[1127]), .rdlo_out(a3_wr[1383]));
			radix2 #(.width(width)) rd_st2_1128  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1128]), .rdlo_in(a2_wr[1384]),  .coef_in(coef[416]), .rdup_out(a3_wr[1128]), .rdlo_out(a3_wr[1384]));
			radix2 #(.width(width)) rd_st2_1129  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1129]), .rdlo_in(a2_wr[1385]),  .coef_in(coef[420]), .rdup_out(a3_wr[1129]), .rdlo_out(a3_wr[1385]));
			radix2 #(.width(width)) rd_st2_1130  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1130]), .rdlo_in(a2_wr[1386]),  .coef_in(coef[424]), .rdup_out(a3_wr[1130]), .rdlo_out(a3_wr[1386]));
			radix2 #(.width(width)) rd_st2_1131  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1131]), .rdlo_in(a2_wr[1387]),  .coef_in(coef[428]), .rdup_out(a3_wr[1131]), .rdlo_out(a3_wr[1387]));
			radix2 #(.width(width)) rd_st2_1132  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1132]), .rdlo_in(a2_wr[1388]),  .coef_in(coef[432]), .rdup_out(a3_wr[1132]), .rdlo_out(a3_wr[1388]));
			radix2 #(.width(width)) rd_st2_1133  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1133]), .rdlo_in(a2_wr[1389]),  .coef_in(coef[436]), .rdup_out(a3_wr[1133]), .rdlo_out(a3_wr[1389]));
			radix2 #(.width(width)) rd_st2_1134  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1134]), .rdlo_in(a2_wr[1390]),  .coef_in(coef[440]), .rdup_out(a3_wr[1134]), .rdlo_out(a3_wr[1390]));
			radix2 #(.width(width)) rd_st2_1135  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1135]), .rdlo_in(a2_wr[1391]),  .coef_in(coef[444]), .rdup_out(a3_wr[1135]), .rdlo_out(a3_wr[1391]));
			radix2 #(.width(width)) rd_st2_1136  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1136]), .rdlo_in(a2_wr[1392]),  .coef_in(coef[448]), .rdup_out(a3_wr[1136]), .rdlo_out(a3_wr[1392]));
			radix2 #(.width(width)) rd_st2_1137  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1137]), .rdlo_in(a2_wr[1393]),  .coef_in(coef[452]), .rdup_out(a3_wr[1137]), .rdlo_out(a3_wr[1393]));
			radix2 #(.width(width)) rd_st2_1138  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1138]), .rdlo_in(a2_wr[1394]),  .coef_in(coef[456]), .rdup_out(a3_wr[1138]), .rdlo_out(a3_wr[1394]));
			radix2 #(.width(width)) rd_st2_1139  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1139]), .rdlo_in(a2_wr[1395]),  .coef_in(coef[460]), .rdup_out(a3_wr[1139]), .rdlo_out(a3_wr[1395]));
			radix2 #(.width(width)) rd_st2_1140  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1140]), .rdlo_in(a2_wr[1396]),  .coef_in(coef[464]), .rdup_out(a3_wr[1140]), .rdlo_out(a3_wr[1396]));
			radix2 #(.width(width)) rd_st2_1141  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1141]), .rdlo_in(a2_wr[1397]),  .coef_in(coef[468]), .rdup_out(a3_wr[1141]), .rdlo_out(a3_wr[1397]));
			radix2 #(.width(width)) rd_st2_1142  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1142]), .rdlo_in(a2_wr[1398]),  .coef_in(coef[472]), .rdup_out(a3_wr[1142]), .rdlo_out(a3_wr[1398]));
			radix2 #(.width(width)) rd_st2_1143  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1143]), .rdlo_in(a2_wr[1399]),  .coef_in(coef[476]), .rdup_out(a3_wr[1143]), .rdlo_out(a3_wr[1399]));
			radix2 #(.width(width)) rd_st2_1144  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1144]), .rdlo_in(a2_wr[1400]),  .coef_in(coef[480]), .rdup_out(a3_wr[1144]), .rdlo_out(a3_wr[1400]));
			radix2 #(.width(width)) rd_st2_1145  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1145]), .rdlo_in(a2_wr[1401]),  .coef_in(coef[484]), .rdup_out(a3_wr[1145]), .rdlo_out(a3_wr[1401]));
			radix2 #(.width(width)) rd_st2_1146  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1146]), .rdlo_in(a2_wr[1402]),  .coef_in(coef[488]), .rdup_out(a3_wr[1146]), .rdlo_out(a3_wr[1402]));
			radix2 #(.width(width)) rd_st2_1147  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1147]), .rdlo_in(a2_wr[1403]),  .coef_in(coef[492]), .rdup_out(a3_wr[1147]), .rdlo_out(a3_wr[1403]));
			radix2 #(.width(width)) rd_st2_1148  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1148]), .rdlo_in(a2_wr[1404]),  .coef_in(coef[496]), .rdup_out(a3_wr[1148]), .rdlo_out(a3_wr[1404]));
			radix2 #(.width(width)) rd_st2_1149  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1149]), .rdlo_in(a2_wr[1405]),  .coef_in(coef[500]), .rdup_out(a3_wr[1149]), .rdlo_out(a3_wr[1405]));
			radix2 #(.width(width)) rd_st2_1150  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1150]), .rdlo_in(a2_wr[1406]),  .coef_in(coef[504]), .rdup_out(a3_wr[1150]), .rdlo_out(a3_wr[1406]));
			radix2 #(.width(width)) rd_st2_1151  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1151]), .rdlo_in(a2_wr[1407]),  .coef_in(coef[508]), .rdup_out(a3_wr[1151]), .rdlo_out(a3_wr[1407]));
			radix2 #(.width(width)) rd_st2_1152  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1152]), .rdlo_in(a2_wr[1408]),  .coef_in(coef[512]), .rdup_out(a3_wr[1152]), .rdlo_out(a3_wr[1408]));
			radix2 #(.width(width)) rd_st2_1153  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1153]), .rdlo_in(a2_wr[1409]),  .coef_in(coef[516]), .rdup_out(a3_wr[1153]), .rdlo_out(a3_wr[1409]));
			radix2 #(.width(width)) rd_st2_1154  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1154]), .rdlo_in(a2_wr[1410]),  .coef_in(coef[520]), .rdup_out(a3_wr[1154]), .rdlo_out(a3_wr[1410]));
			radix2 #(.width(width)) rd_st2_1155  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1155]), .rdlo_in(a2_wr[1411]),  .coef_in(coef[524]), .rdup_out(a3_wr[1155]), .rdlo_out(a3_wr[1411]));
			radix2 #(.width(width)) rd_st2_1156  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1156]), .rdlo_in(a2_wr[1412]),  .coef_in(coef[528]), .rdup_out(a3_wr[1156]), .rdlo_out(a3_wr[1412]));
			radix2 #(.width(width)) rd_st2_1157  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1157]), .rdlo_in(a2_wr[1413]),  .coef_in(coef[532]), .rdup_out(a3_wr[1157]), .rdlo_out(a3_wr[1413]));
			radix2 #(.width(width)) rd_st2_1158  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1158]), .rdlo_in(a2_wr[1414]),  .coef_in(coef[536]), .rdup_out(a3_wr[1158]), .rdlo_out(a3_wr[1414]));
			radix2 #(.width(width)) rd_st2_1159  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1159]), .rdlo_in(a2_wr[1415]),  .coef_in(coef[540]), .rdup_out(a3_wr[1159]), .rdlo_out(a3_wr[1415]));
			radix2 #(.width(width)) rd_st2_1160  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1160]), .rdlo_in(a2_wr[1416]),  .coef_in(coef[544]), .rdup_out(a3_wr[1160]), .rdlo_out(a3_wr[1416]));
			radix2 #(.width(width)) rd_st2_1161  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1161]), .rdlo_in(a2_wr[1417]),  .coef_in(coef[548]), .rdup_out(a3_wr[1161]), .rdlo_out(a3_wr[1417]));
			radix2 #(.width(width)) rd_st2_1162  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1162]), .rdlo_in(a2_wr[1418]),  .coef_in(coef[552]), .rdup_out(a3_wr[1162]), .rdlo_out(a3_wr[1418]));
			radix2 #(.width(width)) rd_st2_1163  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1163]), .rdlo_in(a2_wr[1419]),  .coef_in(coef[556]), .rdup_out(a3_wr[1163]), .rdlo_out(a3_wr[1419]));
			radix2 #(.width(width)) rd_st2_1164  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1164]), .rdlo_in(a2_wr[1420]),  .coef_in(coef[560]), .rdup_out(a3_wr[1164]), .rdlo_out(a3_wr[1420]));
			radix2 #(.width(width)) rd_st2_1165  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1165]), .rdlo_in(a2_wr[1421]),  .coef_in(coef[564]), .rdup_out(a3_wr[1165]), .rdlo_out(a3_wr[1421]));
			radix2 #(.width(width)) rd_st2_1166  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1166]), .rdlo_in(a2_wr[1422]),  .coef_in(coef[568]), .rdup_out(a3_wr[1166]), .rdlo_out(a3_wr[1422]));
			radix2 #(.width(width)) rd_st2_1167  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1167]), .rdlo_in(a2_wr[1423]),  .coef_in(coef[572]), .rdup_out(a3_wr[1167]), .rdlo_out(a3_wr[1423]));
			radix2 #(.width(width)) rd_st2_1168  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1168]), .rdlo_in(a2_wr[1424]),  .coef_in(coef[576]), .rdup_out(a3_wr[1168]), .rdlo_out(a3_wr[1424]));
			radix2 #(.width(width)) rd_st2_1169  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1169]), .rdlo_in(a2_wr[1425]),  .coef_in(coef[580]), .rdup_out(a3_wr[1169]), .rdlo_out(a3_wr[1425]));
			radix2 #(.width(width)) rd_st2_1170  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1170]), .rdlo_in(a2_wr[1426]),  .coef_in(coef[584]), .rdup_out(a3_wr[1170]), .rdlo_out(a3_wr[1426]));
			radix2 #(.width(width)) rd_st2_1171  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1171]), .rdlo_in(a2_wr[1427]),  .coef_in(coef[588]), .rdup_out(a3_wr[1171]), .rdlo_out(a3_wr[1427]));
			radix2 #(.width(width)) rd_st2_1172  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1172]), .rdlo_in(a2_wr[1428]),  .coef_in(coef[592]), .rdup_out(a3_wr[1172]), .rdlo_out(a3_wr[1428]));
			radix2 #(.width(width)) rd_st2_1173  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1173]), .rdlo_in(a2_wr[1429]),  .coef_in(coef[596]), .rdup_out(a3_wr[1173]), .rdlo_out(a3_wr[1429]));
			radix2 #(.width(width)) rd_st2_1174  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1174]), .rdlo_in(a2_wr[1430]),  .coef_in(coef[600]), .rdup_out(a3_wr[1174]), .rdlo_out(a3_wr[1430]));
			radix2 #(.width(width)) rd_st2_1175  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1175]), .rdlo_in(a2_wr[1431]),  .coef_in(coef[604]), .rdup_out(a3_wr[1175]), .rdlo_out(a3_wr[1431]));
			radix2 #(.width(width)) rd_st2_1176  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1176]), .rdlo_in(a2_wr[1432]),  .coef_in(coef[608]), .rdup_out(a3_wr[1176]), .rdlo_out(a3_wr[1432]));
			radix2 #(.width(width)) rd_st2_1177  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1177]), .rdlo_in(a2_wr[1433]),  .coef_in(coef[612]), .rdup_out(a3_wr[1177]), .rdlo_out(a3_wr[1433]));
			radix2 #(.width(width)) rd_st2_1178  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1178]), .rdlo_in(a2_wr[1434]),  .coef_in(coef[616]), .rdup_out(a3_wr[1178]), .rdlo_out(a3_wr[1434]));
			radix2 #(.width(width)) rd_st2_1179  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1179]), .rdlo_in(a2_wr[1435]),  .coef_in(coef[620]), .rdup_out(a3_wr[1179]), .rdlo_out(a3_wr[1435]));
			radix2 #(.width(width)) rd_st2_1180  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1180]), .rdlo_in(a2_wr[1436]),  .coef_in(coef[624]), .rdup_out(a3_wr[1180]), .rdlo_out(a3_wr[1436]));
			radix2 #(.width(width)) rd_st2_1181  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1181]), .rdlo_in(a2_wr[1437]),  .coef_in(coef[628]), .rdup_out(a3_wr[1181]), .rdlo_out(a3_wr[1437]));
			radix2 #(.width(width)) rd_st2_1182  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1182]), .rdlo_in(a2_wr[1438]),  .coef_in(coef[632]), .rdup_out(a3_wr[1182]), .rdlo_out(a3_wr[1438]));
			radix2 #(.width(width)) rd_st2_1183  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1183]), .rdlo_in(a2_wr[1439]),  .coef_in(coef[636]), .rdup_out(a3_wr[1183]), .rdlo_out(a3_wr[1439]));
			radix2 #(.width(width)) rd_st2_1184  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1184]), .rdlo_in(a2_wr[1440]),  .coef_in(coef[640]), .rdup_out(a3_wr[1184]), .rdlo_out(a3_wr[1440]));
			radix2 #(.width(width)) rd_st2_1185  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1185]), .rdlo_in(a2_wr[1441]),  .coef_in(coef[644]), .rdup_out(a3_wr[1185]), .rdlo_out(a3_wr[1441]));
			radix2 #(.width(width)) rd_st2_1186  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1186]), .rdlo_in(a2_wr[1442]),  .coef_in(coef[648]), .rdup_out(a3_wr[1186]), .rdlo_out(a3_wr[1442]));
			radix2 #(.width(width)) rd_st2_1187  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1187]), .rdlo_in(a2_wr[1443]),  .coef_in(coef[652]), .rdup_out(a3_wr[1187]), .rdlo_out(a3_wr[1443]));
			radix2 #(.width(width)) rd_st2_1188  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1188]), .rdlo_in(a2_wr[1444]),  .coef_in(coef[656]), .rdup_out(a3_wr[1188]), .rdlo_out(a3_wr[1444]));
			radix2 #(.width(width)) rd_st2_1189  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1189]), .rdlo_in(a2_wr[1445]),  .coef_in(coef[660]), .rdup_out(a3_wr[1189]), .rdlo_out(a3_wr[1445]));
			radix2 #(.width(width)) rd_st2_1190  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1190]), .rdlo_in(a2_wr[1446]),  .coef_in(coef[664]), .rdup_out(a3_wr[1190]), .rdlo_out(a3_wr[1446]));
			radix2 #(.width(width)) rd_st2_1191  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1191]), .rdlo_in(a2_wr[1447]),  .coef_in(coef[668]), .rdup_out(a3_wr[1191]), .rdlo_out(a3_wr[1447]));
			radix2 #(.width(width)) rd_st2_1192  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1192]), .rdlo_in(a2_wr[1448]),  .coef_in(coef[672]), .rdup_out(a3_wr[1192]), .rdlo_out(a3_wr[1448]));
			radix2 #(.width(width)) rd_st2_1193  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1193]), .rdlo_in(a2_wr[1449]),  .coef_in(coef[676]), .rdup_out(a3_wr[1193]), .rdlo_out(a3_wr[1449]));
			radix2 #(.width(width)) rd_st2_1194  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1194]), .rdlo_in(a2_wr[1450]),  .coef_in(coef[680]), .rdup_out(a3_wr[1194]), .rdlo_out(a3_wr[1450]));
			radix2 #(.width(width)) rd_st2_1195  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1195]), .rdlo_in(a2_wr[1451]),  .coef_in(coef[684]), .rdup_out(a3_wr[1195]), .rdlo_out(a3_wr[1451]));
			radix2 #(.width(width)) rd_st2_1196  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1196]), .rdlo_in(a2_wr[1452]),  .coef_in(coef[688]), .rdup_out(a3_wr[1196]), .rdlo_out(a3_wr[1452]));
			radix2 #(.width(width)) rd_st2_1197  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1197]), .rdlo_in(a2_wr[1453]),  .coef_in(coef[692]), .rdup_out(a3_wr[1197]), .rdlo_out(a3_wr[1453]));
			radix2 #(.width(width)) rd_st2_1198  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1198]), .rdlo_in(a2_wr[1454]),  .coef_in(coef[696]), .rdup_out(a3_wr[1198]), .rdlo_out(a3_wr[1454]));
			radix2 #(.width(width)) rd_st2_1199  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1199]), .rdlo_in(a2_wr[1455]),  .coef_in(coef[700]), .rdup_out(a3_wr[1199]), .rdlo_out(a3_wr[1455]));
			radix2 #(.width(width)) rd_st2_1200  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1200]), .rdlo_in(a2_wr[1456]),  .coef_in(coef[704]), .rdup_out(a3_wr[1200]), .rdlo_out(a3_wr[1456]));
			radix2 #(.width(width)) rd_st2_1201  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1201]), .rdlo_in(a2_wr[1457]),  .coef_in(coef[708]), .rdup_out(a3_wr[1201]), .rdlo_out(a3_wr[1457]));
			radix2 #(.width(width)) rd_st2_1202  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1202]), .rdlo_in(a2_wr[1458]),  .coef_in(coef[712]), .rdup_out(a3_wr[1202]), .rdlo_out(a3_wr[1458]));
			radix2 #(.width(width)) rd_st2_1203  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1203]), .rdlo_in(a2_wr[1459]),  .coef_in(coef[716]), .rdup_out(a3_wr[1203]), .rdlo_out(a3_wr[1459]));
			radix2 #(.width(width)) rd_st2_1204  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1204]), .rdlo_in(a2_wr[1460]),  .coef_in(coef[720]), .rdup_out(a3_wr[1204]), .rdlo_out(a3_wr[1460]));
			radix2 #(.width(width)) rd_st2_1205  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1205]), .rdlo_in(a2_wr[1461]),  .coef_in(coef[724]), .rdup_out(a3_wr[1205]), .rdlo_out(a3_wr[1461]));
			radix2 #(.width(width)) rd_st2_1206  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1206]), .rdlo_in(a2_wr[1462]),  .coef_in(coef[728]), .rdup_out(a3_wr[1206]), .rdlo_out(a3_wr[1462]));
			radix2 #(.width(width)) rd_st2_1207  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1207]), .rdlo_in(a2_wr[1463]),  .coef_in(coef[732]), .rdup_out(a3_wr[1207]), .rdlo_out(a3_wr[1463]));
			radix2 #(.width(width)) rd_st2_1208  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1208]), .rdlo_in(a2_wr[1464]),  .coef_in(coef[736]), .rdup_out(a3_wr[1208]), .rdlo_out(a3_wr[1464]));
			radix2 #(.width(width)) rd_st2_1209  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1209]), .rdlo_in(a2_wr[1465]),  .coef_in(coef[740]), .rdup_out(a3_wr[1209]), .rdlo_out(a3_wr[1465]));
			radix2 #(.width(width)) rd_st2_1210  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1210]), .rdlo_in(a2_wr[1466]),  .coef_in(coef[744]), .rdup_out(a3_wr[1210]), .rdlo_out(a3_wr[1466]));
			radix2 #(.width(width)) rd_st2_1211  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1211]), .rdlo_in(a2_wr[1467]),  .coef_in(coef[748]), .rdup_out(a3_wr[1211]), .rdlo_out(a3_wr[1467]));
			radix2 #(.width(width)) rd_st2_1212  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1212]), .rdlo_in(a2_wr[1468]),  .coef_in(coef[752]), .rdup_out(a3_wr[1212]), .rdlo_out(a3_wr[1468]));
			radix2 #(.width(width)) rd_st2_1213  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1213]), .rdlo_in(a2_wr[1469]),  .coef_in(coef[756]), .rdup_out(a3_wr[1213]), .rdlo_out(a3_wr[1469]));
			radix2 #(.width(width)) rd_st2_1214  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1214]), .rdlo_in(a2_wr[1470]),  .coef_in(coef[760]), .rdup_out(a3_wr[1214]), .rdlo_out(a3_wr[1470]));
			radix2 #(.width(width)) rd_st2_1215  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1215]), .rdlo_in(a2_wr[1471]),  .coef_in(coef[764]), .rdup_out(a3_wr[1215]), .rdlo_out(a3_wr[1471]));
			radix2 #(.width(width)) rd_st2_1216  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1216]), .rdlo_in(a2_wr[1472]),  .coef_in(coef[768]), .rdup_out(a3_wr[1216]), .rdlo_out(a3_wr[1472]));
			radix2 #(.width(width)) rd_st2_1217  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1217]), .rdlo_in(a2_wr[1473]),  .coef_in(coef[772]), .rdup_out(a3_wr[1217]), .rdlo_out(a3_wr[1473]));
			radix2 #(.width(width)) rd_st2_1218  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1218]), .rdlo_in(a2_wr[1474]),  .coef_in(coef[776]), .rdup_out(a3_wr[1218]), .rdlo_out(a3_wr[1474]));
			radix2 #(.width(width)) rd_st2_1219  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1219]), .rdlo_in(a2_wr[1475]),  .coef_in(coef[780]), .rdup_out(a3_wr[1219]), .rdlo_out(a3_wr[1475]));
			radix2 #(.width(width)) rd_st2_1220  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1220]), .rdlo_in(a2_wr[1476]),  .coef_in(coef[784]), .rdup_out(a3_wr[1220]), .rdlo_out(a3_wr[1476]));
			radix2 #(.width(width)) rd_st2_1221  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1221]), .rdlo_in(a2_wr[1477]),  .coef_in(coef[788]), .rdup_out(a3_wr[1221]), .rdlo_out(a3_wr[1477]));
			radix2 #(.width(width)) rd_st2_1222  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1222]), .rdlo_in(a2_wr[1478]),  .coef_in(coef[792]), .rdup_out(a3_wr[1222]), .rdlo_out(a3_wr[1478]));
			radix2 #(.width(width)) rd_st2_1223  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1223]), .rdlo_in(a2_wr[1479]),  .coef_in(coef[796]), .rdup_out(a3_wr[1223]), .rdlo_out(a3_wr[1479]));
			radix2 #(.width(width)) rd_st2_1224  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1224]), .rdlo_in(a2_wr[1480]),  .coef_in(coef[800]), .rdup_out(a3_wr[1224]), .rdlo_out(a3_wr[1480]));
			radix2 #(.width(width)) rd_st2_1225  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1225]), .rdlo_in(a2_wr[1481]),  .coef_in(coef[804]), .rdup_out(a3_wr[1225]), .rdlo_out(a3_wr[1481]));
			radix2 #(.width(width)) rd_st2_1226  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1226]), .rdlo_in(a2_wr[1482]),  .coef_in(coef[808]), .rdup_out(a3_wr[1226]), .rdlo_out(a3_wr[1482]));
			radix2 #(.width(width)) rd_st2_1227  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1227]), .rdlo_in(a2_wr[1483]),  .coef_in(coef[812]), .rdup_out(a3_wr[1227]), .rdlo_out(a3_wr[1483]));
			radix2 #(.width(width)) rd_st2_1228  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1228]), .rdlo_in(a2_wr[1484]),  .coef_in(coef[816]), .rdup_out(a3_wr[1228]), .rdlo_out(a3_wr[1484]));
			radix2 #(.width(width)) rd_st2_1229  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1229]), .rdlo_in(a2_wr[1485]),  .coef_in(coef[820]), .rdup_out(a3_wr[1229]), .rdlo_out(a3_wr[1485]));
			radix2 #(.width(width)) rd_st2_1230  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1230]), .rdlo_in(a2_wr[1486]),  .coef_in(coef[824]), .rdup_out(a3_wr[1230]), .rdlo_out(a3_wr[1486]));
			radix2 #(.width(width)) rd_st2_1231  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1231]), .rdlo_in(a2_wr[1487]),  .coef_in(coef[828]), .rdup_out(a3_wr[1231]), .rdlo_out(a3_wr[1487]));
			radix2 #(.width(width)) rd_st2_1232  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1232]), .rdlo_in(a2_wr[1488]),  .coef_in(coef[832]), .rdup_out(a3_wr[1232]), .rdlo_out(a3_wr[1488]));
			radix2 #(.width(width)) rd_st2_1233  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1233]), .rdlo_in(a2_wr[1489]),  .coef_in(coef[836]), .rdup_out(a3_wr[1233]), .rdlo_out(a3_wr[1489]));
			radix2 #(.width(width)) rd_st2_1234  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1234]), .rdlo_in(a2_wr[1490]),  .coef_in(coef[840]), .rdup_out(a3_wr[1234]), .rdlo_out(a3_wr[1490]));
			radix2 #(.width(width)) rd_st2_1235  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1235]), .rdlo_in(a2_wr[1491]),  .coef_in(coef[844]), .rdup_out(a3_wr[1235]), .rdlo_out(a3_wr[1491]));
			radix2 #(.width(width)) rd_st2_1236  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1236]), .rdlo_in(a2_wr[1492]),  .coef_in(coef[848]), .rdup_out(a3_wr[1236]), .rdlo_out(a3_wr[1492]));
			radix2 #(.width(width)) rd_st2_1237  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1237]), .rdlo_in(a2_wr[1493]),  .coef_in(coef[852]), .rdup_out(a3_wr[1237]), .rdlo_out(a3_wr[1493]));
			radix2 #(.width(width)) rd_st2_1238  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1238]), .rdlo_in(a2_wr[1494]),  .coef_in(coef[856]), .rdup_out(a3_wr[1238]), .rdlo_out(a3_wr[1494]));
			radix2 #(.width(width)) rd_st2_1239  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1239]), .rdlo_in(a2_wr[1495]),  .coef_in(coef[860]), .rdup_out(a3_wr[1239]), .rdlo_out(a3_wr[1495]));
			radix2 #(.width(width)) rd_st2_1240  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1240]), .rdlo_in(a2_wr[1496]),  .coef_in(coef[864]), .rdup_out(a3_wr[1240]), .rdlo_out(a3_wr[1496]));
			radix2 #(.width(width)) rd_st2_1241  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1241]), .rdlo_in(a2_wr[1497]),  .coef_in(coef[868]), .rdup_out(a3_wr[1241]), .rdlo_out(a3_wr[1497]));
			radix2 #(.width(width)) rd_st2_1242  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1242]), .rdlo_in(a2_wr[1498]),  .coef_in(coef[872]), .rdup_out(a3_wr[1242]), .rdlo_out(a3_wr[1498]));
			radix2 #(.width(width)) rd_st2_1243  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1243]), .rdlo_in(a2_wr[1499]),  .coef_in(coef[876]), .rdup_out(a3_wr[1243]), .rdlo_out(a3_wr[1499]));
			radix2 #(.width(width)) rd_st2_1244  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1244]), .rdlo_in(a2_wr[1500]),  .coef_in(coef[880]), .rdup_out(a3_wr[1244]), .rdlo_out(a3_wr[1500]));
			radix2 #(.width(width)) rd_st2_1245  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1245]), .rdlo_in(a2_wr[1501]),  .coef_in(coef[884]), .rdup_out(a3_wr[1245]), .rdlo_out(a3_wr[1501]));
			radix2 #(.width(width)) rd_st2_1246  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1246]), .rdlo_in(a2_wr[1502]),  .coef_in(coef[888]), .rdup_out(a3_wr[1246]), .rdlo_out(a3_wr[1502]));
			radix2 #(.width(width)) rd_st2_1247  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1247]), .rdlo_in(a2_wr[1503]),  .coef_in(coef[892]), .rdup_out(a3_wr[1247]), .rdlo_out(a3_wr[1503]));
			radix2 #(.width(width)) rd_st2_1248  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1248]), .rdlo_in(a2_wr[1504]),  .coef_in(coef[896]), .rdup_out(a3_wr[1248]), .rdlo_out(a3_wr[1504]));
			radix2 #(.width(width)) rd_st2_1249  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1249]), .rdlo_in(a2_wr[1505]),  .coef_in(coef[900]), .rdup_out(a3_wr[1249]), .rdlo_out(a3_wr[1505]));
			radix2 #(.width(width)) rd_st2_1250  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1250]), .rdlo_in(a2_wr[1506]),  .coef_in(coef[904]), .rdup_out(a3_wr[1250]), .rdlo_out(a3_wr[1506]));
			radix2 #(.width(width)) rd_st2_1251  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1251]), .rdlo_in(a2_wr[1507]),  .coef_in(coef[908]), .rdup_out(a3_wr[1251]), .rdlo_out(a3_wr[1507]));
			radix2 #(.width(width)) rd_st2_1252  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1252]), .rdlo_in(a2_wr[1508]),  .coef_in(coef[912]), .rdup_out(a3_wr[1252]), .rdlo_out(a3_wr[1508]));
			radix2 #(.width(width)) rd_st2_1253  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1253]), .rdlo_in(a2_wr[1509]),  .coef_in(coef[916]), .rdup_out(a3_wr[1253]), .rdlo_out(a3_wr[1509]));
			radix2 #(.width(width)) rd_st2_1254  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1254]), .rdlo_in(a2_wr[1510]),  .coef_in(coef[920]), .rdup_out(a3_wr[1254]), .rdlo_out(a3_wr[1510]));
			radix2 #(.width(width)) rd_st2_1255  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1255]), .rdlo_in(a2_wr[1511]),  .coef_in(coef[924]), .rdup_out(a3_wr[1255]), .rdlo_out(a3_wr[1511]));
			radix2 #(.width(width)) rd_st2_1256  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1256]), .rdlo_in(a2_wr[1512]),  .coef_in(coef[928]), .rdup_out(a3_wr[1256]), .rdlo_out(a3_wr[1512]));
			radix2 #(.width(width)) rd_st2_1257  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1257]), .rdlo_in(a2_wr[1513]),  .coef_in(coef[932]), .rdup_out(a3_wr[1257]), .rdlo_out(a3_wr[1513]));
			radix2 #(.width(width)) rd_st2_1258  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1258]), .rdlo_in(a2_wr[1514]),  .coef_in(coef[936]), .rdup_out(a3_wr[1258]), .rdlo_out(a3_wr[1514]));
			radix2 #(.width(width)) rd_st2_1259  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1259]), .rdlo_in(a2_wr[1515]),  .coef_in(coef[940]), .rdup_out(a3_wr[1259]), .rdlo_out(a3_wr[1515]));
			radix2 #(.width(width)) rd_st2_1260  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1260]), .rdlo_in(a2_wr[1516]),  .coef_in(coef[944]), .rdup_out(a3_wr[1260]), .rdlo_out(a3_wr[1516]));
			radix2 #(.width(width)) rd_st2_1261  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1261]), .rdlo_in(a2_wr[1517]),  .coef_in(coef[948]), .rdup_out(a3_wr[1261]), .rdlo_out(a3_wr[1517]));
			radix2 #(.width(width)) rd_st2_1262  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1262]), .rdlo_in(a2_wr[1518]),  .coef_in(coef[952]), .rdup_out(a3_wr[1262]), .rdlo_out(a3_wr[1518]));
			radix2 #(.width(width)) rd_st2_1263  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1263]), .rdlo_in(a2_wr[1519]),  .coef_in(coef[956]), .rdup_out(a3_wr[1263]), .rdlo_out(a3_wr[1519]));
			radix2 #(.width(width)) rd_st2_1264  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1264]), .rdlo_in(a2_wr[1520]),  .coef_in(coef[960]), .rdup_out(a3_wr[1264]), .rdlo_out(a3_wr[1520]));
			radix2 #(.width(width)) rd_st2_1265  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1265]), .rdlo_in(a2_wr[1521]),  .coef_in(coef[964]), .rdup_out(a3_wr[1265]), .rdlo_out(a3_wr[1521]));
			radix2 #(.width(width)) rd_st2_1266  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1266]), .rdlo_in(a2_wr[1522]),  .coef_in(coef[968]), .rdup_out(a3_wr[1266]), .rdlo_out(a3_wr[1522]));
			radix2 #(.width(width)) rd_st2_1267  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1267]), .rdlo_in(a2_wr[1523]),  .coef_in(coef[972]), .rdup_out(a3_wr[1267]), .rdlo_out(a3_wr[1523]));
			radix2 #(.width(width)) rd_st2_1268  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1268]), .rdlo_in(a2_wr[1524]),  .coef_in(coef[976]), .rdup_out(a3_wr[1268]), .rdlo_out(a3_wr[1524]));
			radix2 #(.width(width)) rd_st2_1269  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1269]), .rdlo_in(a2_wr[1525]),  .coef_in(coef[980]), .rdup_out(a3_wr[1269]), .rdlo_out(a3_wr[1525]));
			radix2 #(.width(width)) rd_st2_1270  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1270]), .rdlo_in(a2_wr[1526]),  .coef_in(coef[984]), .rdup_out(a3_wr[1270]), .rdlo_out(a3_wr[1526]));
			radix2 #(.width(width)) rd_st2_1271  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1271]), .rdlo_in(a2_wr[1527]),  .coef_in(coef[988]), .rdup_out(a3_wr[1271]), .rdlo_out(a3_wr[1527]));
			radix2 #(.width(width)) rd_st2_1272  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1272]), .rdlo_in(a2_wr[1528]),  .coef_in(coef[992]), .rdup_out(a3_wr[1272]), .rdlo_out(a3_wr[1528]));
			radix2 #(.width(width)) rd_st2_1273  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1273]), .rdlo_in(a2_wr[1529]),  .coef_in(coef[996]), .rdup_out(a3_wr[1273]), .rdlo_out(a3_wr[1529]));
			radix2 #(.width(width)) rd_st2_1274  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1274]), .rdlo_in(a2_wr[1530]),  .coef_in(coef[1000]), .rdup_out(a3_wr[1274]), .rdlo_out(a3_wr[1530]));
			radix2 #(.width(width)) rd_st2_1275  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1275]), .rdlo_in(a2_wr[1531]),  .coef_in(coef[1004]), .rdup_out(a3_wr[1275]), .rdlo_out(a3_wr[1531]));
			radix2 #(.width(width)) rd_st2_1276  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1276]), .rdlo_in(a2_wr[1532]),  .coef_in(coef[1008]), .rdup_out(a3_wr[1276]), .rdlo_out(a3_wr[1532]));
			radix2 #(.width(width)) rd_st2_1277  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1277]), .rdlo_in(a2_wr[1533]),  .coef_in(coef[1012]), .rdup_out(a3_wr[1277]), .rdlo_out(a3_wr[1533]));
			radix2 #(.width(width)) rd_st2_1278  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1278]), .rdlo_in(a2_wr[1534]),  .coef_in(coef[1016]), .rdup_out(a3_wr[1278]), .rdlo_out(a3_wr[1534]));
			radix2 #(.width(width)) rd_st2_1279  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1279]), .rdlo_in(a2_wr[1535]),  .coef_in(coef[1020]), .rdup_out(a3_wr[1279]), .rdlo_out(a3_wr[1535]));
			radix2 #(.width(width)) rd_st2_1536  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1536]), .rdlo_in(a2_wr[1792]),  .coef_in(coef[0]), .rdup_out(a3_wr[1536]), .rdlo_out(a3_wr[1792]));
			radix2 #(.width(width)) rd_st2_1537  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1537]), .rdlo_in(a2_wr[1793]),  .coef_in(coef[4]), .rdup_out(a3_wr[1537]), .rdlo_out(a3_wr[1793]));
			radix2 #(.width(width)) rd_st2_1538  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1538]), .rdlo_in(a2_wr[1794]),  .coef_in(coef[8]), .rdup_out(a3_wr[1538]), .rdlo_out(a3_wr[1794]));
			radix2 #(.width(width)) rd_st2_1539  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1539]), .rdlo_in(a2_wr[1795]),  .coef_in(coef[12]), .rdup_out(a3_wr[1539]), .rdlo_out(a3_wr[1795]));
			radix2 #(.width(width)) rd_st2_1540  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1540]), .rdlo_in(a2_wr[1796]),  .coef_in(coef[16]), .rdup_out(a3_wr[1540]), .rdlo_out(a3_wr[1796]));
			radix2 #(.width(width)) rd_st2_1541  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1541]), .rdlo_in(a2_wr[1797]),  .coef_in(coef[20]), .rdup_out(a3_wr[1541]), .rdlo_out(a3_wr[1797]));
			radix2 #(.width(width)) rd_st2_1542  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1542]), .rdlo_in(a2_wr[1798]),  .coef_in(coef[24]), .rdup_out(a3_wr[1542]), .rdlo_out(a3_wr[1798]));
			radix2 #(.width(width)) rd_st2_1543  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1543]), .rdlo_in(a2_wr[1799]),  .coef_in(coef[28]), .rdup_out(a3_wr[1543]), .rdlo_out(a3_wr[1799]));
			radix2 #(.width(width)) rd_st2_1544  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1544]), .rdlo_in(a2_wr[1800]),  .coef_in(coef[32]), .rdup_out(a3_wr[1544]), .rdlo_out(a3_wr[1800]));
			radix2 #(.width(width)) rd_st2_1545  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1545]), .rdlo_in(a2_wr[1801]),  .coef_in(coef[36]), .rdup_out(a3_wr[1545]), .rdlo_out(a3_wr[1801]));
			radix2 #(.width(width)) rd_st2_1546  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1546]), .rdlo_in(a2_wr[1802]),  .coef_in(coef[40]), .rdup_out(a3_wr[1546]), .rdlo_out(a3_wr[1802]));
			radix2 #(.width(width)) rd_st2_1547  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1547]), .rdlo_in(a2_wr[1803]),  .coef_in(coef[44]), .rdup_out(a3_wr[1547]), .rdlo_out(a3_wr[1803]));
			radix2 #(.width(width)) rd_st2_1548  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1548]), .rdlo_in(a2_wr[1804]),  .coef_in(coef[48]), .rdup_out(a3_wr[1548]), .rdlo_out(a3_wr[1804]));
			radix2 #(.width(width)) rd_st2_1549  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1549]), .rdlo_in(a2_wr[1805]),  .coef_in(coef[52]), .rdup_out(a3_wr[1549]), .rdlo_out(a3_wr[1805]));
			radix2 #(.width(width)) rd_st2_1550  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1550]), .rdlo_in(a2_wr[1806]),  .coef_in(coef[56]), .rdup_out(a3_wr[1550]), .rdlo_out(a3_wr[1806]));
			radix2 #(.width(width)) rd_st2_1551  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1551]), .rdlo_in(a2_wr[1807]),  .coef_in(coef[60]), .rdup_out(a3_wr[1551]), .rdlo_out(a3_wr[1807]));
			radix2 #(.width(width)) rd_st2_1552  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1552]), .rdlo_in(a2_wr[1808]),  .coef_in(coef[64]), .rdup_out(a3_wr[1552]), .rdlo_out(a3_wr[1808]));
			radix2 #(.width(width)) rd_st2_1553  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1553]), .rdlo_in(a2_wr[1809]),  .coef_in(coef[68]), .rdup_out(a3_wr[1553]), .rdlo_out(a3_wr[1809]));
			radix2 #(.width(width)) rd_st2_1554  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1554]), .rdlo_in(a2_wr[1810]),  .coef_in(coef[72]), .rdup_out(a3_wr[1554]), .rdlo_out(a3_wr[1810]));
			radix2 #(.width(width)) rd_st2_1555  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1555]), .rdlo_in(a2_wr[1811]),  .coef_in(coef[76]), .rdup_out(a3_wr[1555]), .rdlo_out(a3_wr[1811]));
			radix2 #(.width(width)) rd_st2_1556  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1556]), .rdlo_in(a2_wr[1812]),  .coef_in(coef[80]), .rdup_out(a3_wr[1556]), .rdlo_out(a3_wr[1812]));
			radix2 #(.width(width)) rd_st2_1557  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1557]), .rdlo_in(a2_wr[1813]),  .coef_in(coef[84]), .rdup_out(a3_wr[1557]), .rdlo_out(a3_wr[1813]));
			radix2 #(.width(width)) rd_st2_1558  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1558]), .rdlo_in(a2_wr[1814]),  .coef_in(coef[88]), .rdup_out(a3_wr[1558]), .rdlo_out(a3_wr[1814]));
			radix2 #(.width(width)) rd_st2_1559  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1559]), .rdlo_in(a2_wr[1815]),  .coef_in(coef[92]), .rdup_out(a3_wr[1559]), .rdlo_out(a3_wr[1815]));
			radix2 #(.width(width)) rd_st2_1560  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1560]), .rdlo_in(a2_wr[1816]),  .coef_in(coef[96]), .rdup_out(a3_wr[1560]), .rdlo_out(a3_wr[1816]));
			radix2 #(.width(width)) rd_st2_1561  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1561]), .rdlo_in(a2_wr[1817]),  .coef_in(coef[100]), .rdup_out(a3_wr[1561]), .rdlo_out(a3_wr[1817]));
			radix2 #(.width(width)) rd_st2_1562  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1562]), .rdlo_in(a2_wr[1818]),  .coef_in(coef[104]), .rdup_out(a3_wr[1562]), .rdlo_out(a3_wr[1818]));
			radix2 #(.width(width)) rd_st2_1563  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1563]), .rdlo_in(a2_wr[1819]),  .coef_in(coef[108]), .rdup_out(a3_wr[1563]), .rdlo_out(a3_wr[1819]));
			radix2 #(.width(width)) rd_st2_1564  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1564]), .rdlo_in(a2_wr[1820]),  .coef_in(coef[112]), .rdup_out(a3_wr[1564]), .rdlo_out(a3_wr[1820]));
			radix2 #(.width(width)) rd_st2_1565  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1565]), .rdlo_in(a2_wr[1821]),  .coef_in(coef[116]), .rdup_out(a3_wr[1565]), .rdlo_out(a3_wr[1821]));
			radix2 #(.width(width)) rd_st2_1566  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1566]), .rdlo_in(a2_wr[1822]),  .coef_in(coef[120]), .rdup_out(a3_wr[1566]), .rdlo_out(a3_wr[1822]));
			radix2 #(.width(width)) rd_st2_1567  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1567]), .rdlo_in(a2_wr[1823]),  .coef_in(coef[124]), .rdup_out(a3_wr[1567]), .rdlo_out(a3_wr[1823]));
			radix2 #(.width(width)) rd_st2_1568  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1568]), .rdlo_in(a2_wr[1824]),  .coef_in(coef[128]), .rdup_out(a3_wr[1568]), .rdlo_out(a3_wr[1824]));
			radix2 #(.width(width)) rd_st2_1569  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1569]), .rdlo_in(a2_wr[1825]),  .coef_in(coef[132]), .rdup_out(a3_wr[1569]), .rdlo_out(a3_wr[1825]));
			radix2 #(.width(width)) rd_st2_1570  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1570]), .rdlo_in(a2_wr[1826]),  .coef_in(coef[136]), .rdup_out(a3_wr[1570]), .rdlo_out(a3_wr[1826]));
			radix2 #(.width(width)) rd_st2_1571  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1571]), .rdlo_in(a2_wr[1827]),  .coef_in(coef[140]), .rdup_out(a3_wr[1571]), .rdlo_out(a3_wr[1827]));
			radix2 #(.width(width)) rd_st2_1572  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1572]), .rdlo_in(a2_wr[1828]),  .coef_in(coef[144]), .rdup_out(a3_wr[1572]), .rdlo_out(a3_wr[1828]));
			radix2 #(.width(width)) rd_st2_1573  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1573]), .rdlo_in(a2_wr[1829]),  .coef_in(coef[148]), .rdup_out(a3_wr[1573]), .rdlo_out(a3_wr[1829]));
			radix2 #(.width(width)) rd_st2_1574  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1574]), .rdlo_in(a2_wr[1830]),  .coef_in(coef[152]), .rdup_out(a3_wr[1574]), .rdlo_out(a3_wr[1830]));
			radix2 #(.width(width)) rd_st2_1575  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1575]), .rdlo_in(a2_wr[1831]),  .coef_in(coef[156]), .rdup_out(a3_wr[1575]), .rdlo_out(a3_wr[1831]));
			radix2 #(.width(width)) rd_st2_1576  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1576]), .rdlo_in(a2_wr[1832]),  .coef_in(coef[160]), .rdup_out(a3_wr[1576]), .rdlo_out(a3_wr[1832]));
			radix2 #(.width(width)) rd_st2_1577  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1577]), .rdlo_in(a2_wr[1833]),  .coef_in(coef[164]), .rdup_out(a3_wr[1577]), .rdlo_out(a3_wr[1833]));
			radix2 #(.width(width)) rd_st2_1578  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1578]), .rdlo_in(a2_wr[1834]),  .coef_in(coef[168]), .rdup_out(a3_wr[1578]), .rdlo_out(a3_wr[1834]));
			radix2 #(.width(width)) rd_st2_1579  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1579]), .rdlo_in(a2_wr[1835]),  .coef_in(coef[172]), .rdup_out(a3_wr[1579]), .rdlo_out(a3_wr[1835]));
			radix2 #(.width(width)) rd_st2_1580  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1580]), .rdlo_in(a2_wr[1836]),  .coef_in(coef[176]), .rdup_out(a3_wr[1580]), .rdlo_out(a3_wr[1836]));
			radix2 #(.width(width)) rd_st2_1581  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1581]), .rdlo_in(a2_wr[1837]),  .coef_in(coef[180]), .rdup_out(a3_wr[1581]), .rdlo_out(a3_wr[1837]));
			radix2 #(.width(width)) rd_st2_1582  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1582]), .rdlo_in(a2_wr[1838]),  .coef_in(coef[184]), .rdup_out(a3_wr[1582]), .rdlo_out(a3_wr[1838]));
			radix2 #(.width(width)) rd_st2_1583  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1583]), .rdlo_in(a2_wr[1839]),  .coef_in(coef[188]), .rdup_out(a3_wr[1583]), .rdlo_out(a3_wr[1839]));
			radix2 #(.width(width)) rd_st2_1584  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1584]), .rdlo_in(a2_wr[1840]),  .coef_in(coef[192]), .rdup_out(a3_wr[1584]), .rdlo_out(a3_wr[1840]));
			radix2 #(.width(width)) rd_st2_1585  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1585]), .rdlo_in(a2_wr[1841]),  .coef_in(coef[196]), .rdup_out(a3_wr[1585]), .rdlo_out(a3_wr[1841]));
			radix2 #(.width(width)) rd_st2_1586  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1586]), .rdlo_in(a2_wr[1842]),  .coef_in(coef[200]), .rdup_out(a3_wr[1586]), .rdlo_out(a3_wr[1842]));
			radix2 #(.width(width)) rd_st2_1587  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1587]), .rdlo_in(a2_wr[1843]),  .coef_in(coef[204]), .rdup_out(a3_wr[1587]), .rdlo_out(a3_wr[1843]));
			radix2 #(.width(width)) rd_st2_1588  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1588]), .rdlo_in(a2_wr[1844]),  .coef_in(coef[208]), .rdup_out(a3_wr[1588]), .rdlo_out(a3_wr[1844]));
			radix2 #(.width(width)) rd_st2_1589  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1589]), .rdlo_in(a2_wr[1845]),  .coef_in(coef[212]), .rdup_out(a3_wr[1589]), .rdlo_out(a3_wr[1845]));
			radix2 #(.width(width)) rd_st2_1590  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1590]), .rdlo_in(a2_wr[1846]),  .coef_in(coef[216]), .rdup_out(a3_wr[1590]), .rdlo_out(a3_wr[1846]));
			radix2 #(.width(width)) rd_st2_1591  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1591]), .rdlo_in(a2_wr[1847]),  .coef_in(coef[220]), .rdup_out(a3_wr[1591]), .rdlo_out(a3_wr[1847]));
			radix2 #(.width(width)) rd_st2_1592  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1592]), .rdlo_in(a2_wr[1848]),  .coef_in(coef[224]), .rdup_out(a3_wr[1592]), .rdlo_out(a3_wr[1848]));
			radix2 #(.width(width)) rd_st2_1593  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1593]), .rdlo_in(a2_wr[1849]),  .coef_in(coef[228]), .rdup_out(a3_wr[1593]), .rdlo_out(a3_wr[1849]));
			radix2 #(.width(width)) rd_st2_1594  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1594]), .rdlo_in(a2_wr[1850]),  .coef_in(coef[232]), .rdup_out(a3_wr[1594]), .rdlo_out(a3_wr[1850]));
			radix2 #(.width(width)) rd_st2_1595  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1595]), .rdlo_in(a2_wr[1851]),  .coef_in(coef[236]), .rdup_out(a3_wr[1595]), .rdlo_out(a3_wr[1851]));
			radix2 #(.width(width)) rd_st2_1596  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1596]), .rdlo_in(a2_wr[1852]),  .coef_in(coef[240]), .rdup_out(a3_wr[1596]), .rdlo_out(a3_wr[1852]));
			radix2 #(.width(width)) rd_st2_1597  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1597]), .rdlo_in(a2_wr[1853]),  .coef_in(coef[244]), .rdup_out(a3_wr[1597]), .rdlo_out(a3_wr[1853]));
			radix2 #(.width(width)) rd_st2_1598  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1598]), .rdlo_in(a2_wr[1854]),  .coef_in(coef[248]), .rdup_out(a3_wr[1598]), .rdlo_out(a3_wr[1854]));
			radix2 #(.width(width)) rd_st2_1599  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1599]), .rdlo_in(a2_wr[1855]),  .coef_in(coef[252]), .rdup_out(a3_wr[1599]), .rdlo_out(a3_wr[1855]));
			radix2 #(.width(width)) rd_st2_1600  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1600]), .rdlo_in(a2_wr[1856]),  .coef_in(coef[256]), .rdup_out(a3_wr[1600]), .rdlo_out(a3_wr[1856]));
			radix2 #(.width(width)) rd_st2_1601  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1601]), .rdlo_in(a2_wr[1857]),  .coef_in(coef[260]), .rdup_out(a3_wr[1601]), .rdlo_out(a3_wr[1857]));
			radix2 #(.width(width)) rd_st2_1602  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1602]), .rdlo_in(a2_wr[1858]),  .coef_in(coef[264]), .rdup_out(a3_wr[1602]), .rdlo_out(a3_wr[1858]));
			radix2 #(.width(width)) rd_st2_1603  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1603]), .rdlo_in(a2_wr[1859]),  .coef_in(coef[268]), .rdup_out(a3_wr[1603]), .rdlo_out(a3_wr[1859]));
			radix2 #(.width(width)) rd_st2_1604  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1604]), .rdlo_in(a2_wr[1860]),  .coef_in(coef[272]), .rdup_out(a3_wr[1604]), .rdlo_out(a3_wr[1860]));
			radix2 #(.width(width)) rd_st2_1605  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1605]), .rdlo_in(a2_wr[1861]),  .coef_in(coef[276]), .rdup_out(a3_wr[1605]), .rdlo_out(a3_wr[1861]));
			radix2 #(.width(width)) rd_st2_1606  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1606]), .rdlo_in(a2_wr[1862]),  .coef_in(coef[280]), .rdup_out(a3_wr[1606]), .rdlo_out(a3_wr[1862]));
			radix2 #(.width(width)) rd_st2_1607  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1607]), .rdlo_in(a2_wr[1863]),  .coef_in(coef[284]), .rdup_out(a3_wr[1607]), .rdlo_out(a3_wr[1863]));
			radix2 #(.width(width)) rd_st2_1608  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1608]), .rdlo_in(a2_wr[1864]),  .coef_in(coef[288]), .rdup_out(a3_wr[1608]), .rdlo_out(a3_wr[1864]));
			radix2 #(.width(width)) rd_st2_1609  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1609]), .rdlo_in(a2_wr[1865]),  .coef_in(coef[292]), .rdup_out(a3_wr[1609]), .rdlo_out(a3_wr[1865]));
			radix2 #(.width(width)) rd_st2_1610  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1610]), .rdlo_in(a2_wr[1866]),  .coef_in(coef[296]), .rdup_out(a3_wr[1610]), .rdlo_out(a3_wr[1866]));
			radix2 #(.width(width)) rd_st2_1611  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1611]), .rdlo_in(a2_wr[1867]),  .coef_in(coef[300]), .rdup_out(a3_wr[1611]), .rdlo_out(a3_wr[1867]));
			radix2 #(.width(width)) rd_st2_1612  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1612]), .rdlo_in(a2_wr[1868]),  .coef_in(coef[304]), .rdup_out(a3_wr[1612]), .rdlo_out(a3_wr[1868]));
			radix2 #(.width(width)) rd_st2_1613  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1613]), .rdlo_in(a2_wr[1869]),  .coef_in(coef[308]), .rdup_out(a3_wr[1613]), .rdlo_out(a3_wr[1869]));
			radix2 #(.width(width)) rd_st2_1614  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1614]), .rdlo_in(a2_wr[1870]),  .coef_in(coef[312]), .rdup_out(a3_wr[1614]), .rdlo_out(a3_wr[1870]));
			radix2 #(.width(width)) rd_st2_1615  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1615]), .rdlo_in(a2_wr[1871]),  .coef_in(coef[316]), .rdup_out(a3_wr[1615]), .rdlo_out(a3_wr[1871]));
			radix2 #(.width(width)) rd_st2_1616  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1616]), .rdlo_in(a2_wr[1872]),  .coef_in(coef[320]), .rdup_out(a3_wr[1616]), .rdlo_out(a3_wr[1872]));
			radix2 #(.width(width)) rd_st2_1617  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1617]), .rdlo_in(a2_wr[1873]),  .coef_in(coef[324]), .rdup_out(a3_wr[1617]), .rdlo_out(a3_wr[1873]));
			radix2 #(.width(width)) rd_st2_1618  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1618]), .rdlo_in(a2_wr[1874]),  .coef_in(coef[328]), .rdup_out(a3_wr[1618]), .rdlo_out(a3_wr[1874]));
			radix2 #(.width(width)) rd_st2_1619  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1619]), .rdlo_in(a2_wr[1875]),  .coef_in(coef[332]), .rdup_out(a3_wr[1619]), .rdlo_out(a3_wr[1875]));
			radix2 #(.width(width)) rd_st2_1620  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1620]), .rdlo_in(a2_wr[1876]),  .coef_in(coef[336]), .rdup_out(a3_wr[1620]), .rdlo_out(a3_wr[1876]));
			radix2 #(.width(width)) rd_st2_1621  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1621]), .rdlo_in(a2_wr[1877]),  .coef_in(coef[340]), .rdup_out(a3_wr[1621]), .rdlo_out(a3_wr[1877]));
			radix2 #(.width(width)) rd_st2_1622  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1622]), .rdlo_in(a2_wr[1878]),  .coef_in(coef[344]), .rdup_out(a3_wr[1622]), .rdlo_out(a3_wr[1878]));
			radix2 #(.width(width)) rd_st2_1623  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1623]), .rdlo_in(a2_wr[1879]),  .coef_in(coef[348]), .rdup_out(a3_wr[1623]), .rdlo_out(a3_wr[1879]));
			radix2 #(.width(width)) rd_st2_1624  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1624]), .rdlo_in(a2_wr[1880]),  .coef_in(coef[352]), .rdup_out(a3_wr[1624]), .rdlo_out(a3_wr[1880]));
			radix2 #(.width(width)) rd_st2_1625  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1625]), .rdlo_in(a2_wr[1881]),  .coef_in(coef[356]), .rdup_out(a3_wr[1625]), .rdlo_out(a3_wr[1881]));
			radix2 #(.width(width)) rd_st2_1626  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1626]), .rdlo_in(a2_wr[1882]),  .coef_in(coef[360]), .rdup_out(a3_wr[1626]), .rdlo_out(a3_wr[1882]));
			radix2 #(.width(width)) rd_st2_1627  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1627]), .rdlo_in(a2_wr[1883]),  .coef_in(coef[364]), .rdup_out(a3_wr[1627]), .rdlo_out(a3_wr[1883]));
			radix2 #(.width(width)) rd_st2_1628  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1628]), .rdlo_in(a2_wr[1884]),  .coef_in(coef[368]), .rdup_out(a3_wr[1628]), .rdlo_out(a3_wr[1884]));
			radix2 #(.width(width)) rd_st2_1629  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1629]), .rdlo_in(a2_wr[1885]),  .coef_in(coef[372]), .rdup_out(a3_wr[1629]), .rdlo_out(a3_wr[1885]));
			radix2 #(.width(width)) rd_st2_1630  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1630]), .rdlo_in(a2_wr[1886]),  .coef_in(coef[376]), .rdup_out(a3_wr[1630]), .rdlo_out(a3_wr[1886]));
			radix2 #(.width(width)) rd_st2_1631  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1631]), .rdlo_in(a2_wr[1887]),  .coef_in(coef[380]), .rdup_out(a3_wr[1631]), .rdlo_out(a3_wr[1887]));
			radix2 #(.width(width)) rd_st2_1632  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1632]), .rdlo_in(a2_wr[1888]),  .coef_in(coef[384]), .rdup_out(a3_wr[1632]), .rdlo_out(a3_wr[1888]));
			radix2 #(.width(width)) rd_st2_1633  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1633]), .rdlo_in(a2_wr[1889]),  .coef_in(coef[388]), .rdup_out(a3_wr[1633]), .rdlo_out(a3_wr[1889]));
			radix2 #(.width(width)) rd_st2_1634  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1634]), .rdlo_in(a2_wr[1890]),  .coef_in(coef[392]), .rdup_out(a3_wr[1634]), .rdlo_out(a3_wr[1890]));
			radix2 #(.width(width)) rd_st2_1635  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1635]), .rdlo_in(a2_wr[1891]),  .coef_in(coef[396]), .rdup_out(a3_wr[1635]), .rdlo_out(a3_wr[1891]));
			radix2 #(.width(width)) rd_st2_1636  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1636]), .rdlo_in(a2_wr[1892]),  .coef_in(coef[400]), .rdup_out(a3_wr[1636]), .rdlo_out(a3_wr[1892]));
			radix2 #(.width(width)) rd_st2_1637  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1637]), .rdlo_in(a2_wr[1893]),  .coef_in(coef[404]), .rdup_out(a3_wr[1637]), .rdlo_out(a3_wr[1893]));
			radix2 #(.width(width)) rd_st2_1638  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1638]), .rdlo_in(a2_wr[1894]),  .coef_in(coef[408]), .rdup_out(a3_wr[1638]), .rdlo_out(a3_wr[1894]));
			radix2 #(.width(width)) rd_st2_1639  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1639]), .rdlo_in(a2_wr[1895]),  .coef_in(coef[412]), .rdup_out(a3_wr[1639]), .rdlo_out(a3_wr[1895]));
			radix2 #(.width(width)) rd_st2_1640  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1640]), .rdlo_in(a2_wr[1896]),  .coef_in(coef[416]), .rdup_out(a3_wr[1640]), .rdlo_out(a3_wr[1896]));
			radix2 #(.width(width)) rd_st2_1641  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1641]), .rdlo_in(a2_wr[1897]),  .coef_in(coef[420]), .rdup_out(a3_wr[1641]), .rdlo_out(a3_wr[1897]));
			radix2 #(.width(width)) rd_st2_1642  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1642]), .rdlo_in(a2_wr[1898]),  .coef_in(coef[424]), .rdup_out(a3_wr[1642]), .rdlo_out(a3_wr[1898]));
			radix2 #(.width(width)) rd_st2_1643  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1643]), .rdlo_in(a2_wr[1899]),  .coef_in(coef[428]), .rdup_out(a3_wr[1643]), .rdlo_out(a3_wr[1899]));
			radix2 #(.width(width)) rd_st2_1644  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1644]), .rdlo_in(a2_wr[1900]),  .coef_in(coef[432]), .rdup_out(a3_wr[1644]), .rdlo_out(a3_wr[1900]));
			radix2 #(.width(width)) rd_st2_1645  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1645]), .rdlo_in(a2_wr[1901]),  .coef_in(coef[436]), .rdup_out(a3_wr[1645]), .rdlo_out(a3_wr[1901]));
			radix2 #(.width(width)) rd_st2_1646  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1646]), .rdlo_in(a2_wr[1902]),  .coef_in(coef[440]), .rdup_out(a3_wr[1646]), .rdlo_out(a3_wr[1902]));
			radix2 #(.width(width)) rd_st2_1647  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1647]), .rdlo_in(a2_wr[1903]),  .coef_in(coef[444]), .rdup_out(a3_wr[1647]), .rdlo_out(a3_wr[1903]));
			radix2 #(.width(width)) rd_st2_1648  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1648]), .rdlo_in(a2_wr[1904]),  .coef_in(coef[448]), .rdup_out(a3_wr[1648]), .rdlo_out(a3_wr[1904]));
			radix2 #(.width(width)) rd_st2_1649  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1649]), .rdlo_in(a2_wr[1905]),  .coef_in(coef[452]), .rdup_out(a3_wr[1649]), .rdlo_out(a3_wr[1905]));
			radix2 #(.width(width)) rd_st2_1650  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1650]), .rdlo_in(a2_wr[1906]),  .coef_in(coef[456]), .rdup_out(a3_wr[1650]), .rdlo_out(a3_wr[1906]));
			radix2 #(.width(width)) rd_st2_1651  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1651]), .rdlo_in(a2_wr[1907]),  .coef_in(coef[460]), .rdup_out(a3_wr[1651]), .rdlo_out(a3_wr[1907]));
			radix2 #(.width(width)) rd_st2_1652  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1652]), .rdlo_in(a2_wr[1908]),  .coef_in(coef[464]), .rdup_out(a3_wr[1652]), .rdlo_out(a3_wr[1908]));
			radix2 #(.width(width)) rd_st2_1653  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1653]), .rdlo_in(a2_wr[1909]),  .coef_in(coef[468]), .rdup_out(a3_wr[1653]), .rdlo_out(a3_wr[1909]));
			radix2 #(.width(width)) rd_st2_1654  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1654]), .rdlo_in(a2_wr[1910]),  .coef_in(coef[472]), .rdup_out(a3_wr[1654]), .rdlo_out(a3_wr[1910]));
			radix2 #(.width(width)) rd_st2_1655  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1655]), .rdlo_in(a2_wr[1911]),  .coef_in(coef[476]), .rdup_out(a3_wr[1655]), .rdlo_out(a3_wr[1911]));
			radix2 #(.width(width)) rd_st2_1656  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1656]), .rdlo_in(a2_wr[1912]),  .coef_in(coef[480]), .rdup_out(a3_wr[1656]), .rdlo_out(a3_wr[1912]));
			radix2 #(.width(width)) rd_st2_1657  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1657]), .rdlo_in(a2_wr[1913]),  .coef_in(coef[484]), .rdup_out(a3_wr[1657]), .rdlo_out(a3_wr[1913]));
			radix2 #(.width(width)) rd_st2_1658  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1658]), .rdlo_in(a2_wr[1914]),  .coef_in(coef[488]), .rdup_out(a3_wr[1658]), .rdlo_out(a3_wr[1914]));
			radix2 #(.width(width)) rd_st2_1659  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1659]), .rdlo_in(a2_wr[1915]),  .coef_in(coef[492]), .rdup_out(a3_wr[1659]), .rdlo_out(a3_wr[1915]));
			radix2 #(.width(width)) rd_st2_1660  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1660]), .rdlo_in(a2_wr[1916]),  .coef_in(coef[496]), .rdup_out(a3_wr[1660]), .rdlo_out(a3_wr[1916]));
			radix2 #(.width(width)) rd_st2_1661  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1661]), .rdlo_in(a2_wr[1917]),  .coef_in(coef[500]), .rdup_out(a3_wr[1661]), .rdlo_out(a3_wr[1917]));
			radix2 #(.width(width)) rd_st2_1662  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1662]), .rdlo_in(a2_wr[1918]),  .coef_in(coef[504]), .rdup_out(a3_wr[1662]), .rdlo_out(a3_wr[1918]));
			radix2 #(.width(width)) rd_st2_1663  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1663]), .rdlo_in(a2_wr[1919]),  .coef_in(coef[508]), .rdup_out(a3_wr[1663]), .rdlo_out(a3_wr[1919]));
			radix2 #(.width(width)) rd_st2_1664  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1664]), .rdlo_in(a2_wr[1920]),  .coef_in(coef[512]), .rdup_out(a3_wr[1664]), .rdlo_out(a3_wr[1920]));
			radix2 #(.width(width)) rd_st2_1665  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1665]), .rdlo_in(a2_wr[1921]),  .coef_in(coef[516]), .rdup_out(a3_wr[1665]), .rdlo_out(a3_wr[1921]));
			radix2 #(.width(width)) rd_st2_1666  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1666]), .rdlo_in(a2_wr[1922]),  .coef_in(coef[520]), .rdup_out(a3_wr[1666]), .rdlo_out(a3_wr[1922]));
			radix2 #(.width(width)) rd_st2_1667  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1667]), .rdlo_in(a2_wr[1923]),  .coef_in(coef[524]), .rdup_out(a3_wr[1667]), .rdlo_out(a3_wr[1923]));
			radix2 #(.width(width)) rd_st2_1668  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1668]), .rdlo_in(a2_wr[1924]),  .coef_in(coef[528]), .rdup_out(a3_wr[1668]), .rdlo_out(a3_wr[1924]));
			radix2 #(.width(width)) rd_st2_1669  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1669]), .rdlo_in(a2_wr[1925]),  .coef_in(coef[532]), .rdup_out(a3_wr[1669]), .rdlo_out(a3_wr[1925]));
			radix2 #(.width(width)) rd_st2_1670  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1670]), .rdlo_in(a2_wr[1926]),  .coef_in(coef[536]), .rdup_out(a3_wr[1670]), .rdlo_out(a3_wr[1926]));
			radix2 #(.width(width)) rd_st2_1671  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1671]), .rdlo_in(a2_wr[1927]),  .coef_in(coef[540]), .rdup_out(a3_wr[1671]), .rdlo_out(a3_wr[1927]));
			radix2 #(.width(width)) rd_st2_1672  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1672]), .rdlo_in(a2_wr[1928]),  .coef_in(coef[544]), .rdup_out(a3_wr[1672]), .rdlo_out(a3_wr[1928]));
			radix2 #(.width(width)) rd_st2_1673  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1673]), .rdlo_in(a2_wr[1929]),  .coef_in(coef[548]), .rdup_out(a3_wr[1673]), .rdlo_out(a3_wr[1929]));
			radix2 #(.width(width)) rd_st2_1674  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1674]), .rdlo_in(a2_wr[1930]),  .coef_in(coef[552]), .rdup_out(a3_wr[1674]), .rdlo_out(a3_wr[1930]));
			radix2 #(.width(width)) rd_st2_1675  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1675]), .rdlo_in(a2_wr[1931]),  .coef_in(coef[556]), .rdup_out(a3_wr[1675]), .rdlo_out(a3_wr[1931]));
			radix2 #(.width(width)) rd_st2_1676  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1676]), .rdlo_in(a2_wr[1932]),  .coef_in(coef[560]), .rdup_out(a3_wr[1676]), .rdlo_out(a3_wr[1932]));
			radix2 #(.width(width)) rd_st2_1677  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1677]), .rdlo_in(a2_wr[1933]),  .coef_in(coef[564]), .rdup_out(a3_wr[1677]), .rdlo_out(a3_wr[1933]));
			radix2 #(.width(width)) rd_st2_1678  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1678]), .rdlo_in(a2_wr[1934]),  .coef_in(coef[568]), .rdup_out(a3_wr[1678]), .rdlo_out(a3_wr[1934]));
			radix2 #(.width(width)) rd_st2_1679  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1679]), .rdlo_in(a2_wr[1935]),  .coef_in(coef[572]), .rdup_out(a3_wr[1679]), .rdlo_out(a3_wr[1935]));
			radix2 #(.width(width)) rd_st2_1680  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1680]), .rdlo_in(a2_wr[1936]),  .coef_in(coef[576]), .rdup_out(a3_wr[1680]), .rdlo_out(a3_wr[1936]));
			radix2 #(.width(width)) rd_st2_1681  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1681]), .rdlo_in(a2_wr[1937]),  .coef_in(coef[580]), .rdup_out(a3_wr[1681]), .rdlo_out(a3_wr[1937]));
			radix2 #(.width(width)) rd_st2_1682  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1682]), .rdlo_in(a2_wr[1938]),  .coef_in(coef[584]), .rdup_out(a3_wr[1682]), .rdlo_out(a3_wr[1938]));
			radix2 #(.width(width)) rd_st2_1683  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1683]), .rdlo_in(a2_wr[1939]),  .coef_in(coef[588]), .rdup_out(a3_wr[1683]), .rdlo_out(a3_wr[1939]));
			radix2 #(.width(width)) rd_st2_1684  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1684]), .rdlo_in(a2_wr[1940]),  .coef_in(coef[592]), .rdup_out(a3_wr[1684]), .rdlo_out(a3_wr[1940]));
			radix2 #(.width(width)) rd_st2_1685  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1685]), .rdlo_in(a2_wr[1941]),  .coef_in(coef[596]), .rdup_out(a3_wr[1685]), .rdlo_out(a3_wr[1941]));
			radix2 #(.width(width)) rd_st2_1686  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1686]), .rdlo_in(a2_wr[1942]),  .coef_in(coef[600]), .rdup_out(a3_wr[1686]), .rdlo_out(a3_wr[1942]));
			radix2 #(.width(width)) rd_st2_1687  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1687]), .rdlo_in(a2_wr[1943]),  .coef_in(coef[604]), .rdup_out(a3_wr[1687]), .rdlo_out(a3_wr[1943]));
			radix2 #(.width(width)) rd_st2_1688  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1688]), .rdlo_in(a2_wr[1944]),  .coef_in(coef[608]), .rdup_out(a3_wr[1688]), .rdlo_out(a3_wr[1944]));
			radix2 #(.width(width)) rd_st2_1689  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1689]), .rdlo_in(a2_wr[1945]),  .coef_in(coef[612]), .rdup_out(a3_wr[1689]), .rdlo_out(a3_wr[1945]));
			radix2 #(.width(width)) rd_st2_1690  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1690]), .rdlo_in(a2_wr[1946]),  .coef_in(coef[616]), .rdup_out(a3_wr[1690]), .rdlo_out(a3_wr[1946]));
			radix2 #(.width(width)) rd_st2_1691  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1691]), .rdlo_in(a2_wr[1947]),  .coef_in(coef[620]), .rdup_out(a3_wr[1691]), .rdlo_out(a3_wr[1947]));
			radix2 #(.width(width)) rd_st2_1692  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1692]), .rdlo_in(a2_wr[1948]),  .coef_in(coef[624]), .rdup_out(a3_wr[1692]), .rdlo_out(a3_wr[1948]));
			radix2 #(.width(width)) rd_st2_1693  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1693]), .rdlo_in(a2_wr[1949]),  .coef_in(coef[628]), .rdup_out(a3_wr[1693]), .rdlo_out(a3_wr[1949]));
			radix2 #(.width(width)) rd_st2_1694  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1694]), .rdlo_in(a2_wr[1950]),  .coef_in(coef[632]), .rdup_out(a3_wr[1694]), .rdlo_out(a3_wr[1950]));
			radix2 #(.width(width)) rd_st2_1695  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1695]), .rdlo_in(a2_wr[1951]),  .coef_in(coef[636]), .rdup_out(a3_wr[1695]), .rdlo_out(a3_wr[1951]));
			radix2 #(.width(width)) rd_st2_1696  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1696]), .rdlo_in(a2_wr[1952]),  .coef_in(coef[640]), .rdup_out(a3_wr[1696]), .rdlo_out(a3_wr[1952]));
			radix2 #(.width(width)) rd_st2_1697  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1697]), .rdlo_in(a2_wr[1953]),  .coef_in(coef[644]), .rdup_out(a3_wr[1697]), .rdlo_out(a3_wr[1953]));
			radix2 #(.width(width)) rd_st2_1698  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1698]), .rdlo_in(a2_wr[1954]),  .coef_in(coef[648]), .rdup_out(a3_wr[1698]), .rdlo_out(a3_wr[1954]));
			radix2 #(.width(width)) rd_st2_1699  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1699]), .rdlo_in(a2_wr[1955]),  .coef_in(coef[652]), .rdup_out(a3_wr[1699]), .rdlo_out(a3_wr[1955]));
			radix2 #(.width(width)) rd_st2_1700  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1700]), .rdlo_in(a2_wr[1956]),  .coef_in(coef[656]), .rdup_out(a3_wr[1700]), .rdlo_out(a3_wr[1956]));
			radix2 #(.width(width)) rd_st2_1701  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1701]), .rdlo_in(a2_wr[1957]),  .coef_in(coef[660]), .rdup_out(a3_wr[1701]), .rdlo_out(a3_wr[1957]));
			radix2 #(.width(width)) rd_st2_1702  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1702]), .rdlo_in(a2_wr[1958]),  .coef_in(coef[664]), .rdup_out(a3_wr[1702]), .rdlo_out(a3_wr[1958]));
			radix2 #(.width(width)) rd_st2_1703  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1703]), .rdlo_in(a2_wr[1959]),  .coef_in(coef[668]), .rdup_out(a3_wr[1703]), .rdlo_out(a3_wr[1959]));
			radix2 #(.width(width)) rd_st2_1704  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1704]), .rdlo_in(a2_wr[1960]),  .coef_in(coef[672]), .rdup_out(a3_wr[1704]), .rdlo_out(a3_wr[1960]));
			radix2 #(.width(width)) rd_st2_1705  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1705]), .rdlo_in(a2_wr[1961]),  .coef_in(coef[676]), .rdup_out(a3_wr[1705]), .rdlo_out(a3_wr[1961]));
			radix2 #(.width(width)) rd_st2_1706  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1706]), .rdlo_in(a2_wr[1962]),  .coef_in(coef[680]), .rdup_out(a3_wr[1706]), .rdlo_out(a3_wr[1962]));
			radix2 #(.width(width)) rd_st2_1707  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1707]), .rdlo_in(a2_wr[1963]),  .coef_in(coef[684]), .rdup_out(a3_wr[1707]), .rdlo_out(a3_wr[1963]));
			radix2 #(.width(width)) rd_st2_1708  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1708]), .rdlo_in(a2_wr[1964]),  .coef_in(coef[688]), .rdup_out(a3_wr[1708]), .rdlo_out(a3_wr[1964]));
			radix2 #(.width(width)) rd_st2_1709  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1709]), .rdlo_in(a2_wr[1965]),  .coef_in(coef[692]), .rdup_out(a3_wr[1709]), .rdlo_out(a3_wr[1965]));
			radix2 #(.width(width)) rd_st2_1710  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1710]), .rdlo_in(a2_wr[1966]),  .coef_in(coef[696]), .rdup_out(a3_wr[1710]), .rdlo_out(a3_wr[1966]));
			radix2 #(.width(width)) rd_st2_1711  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1711]), .rdlo_in(a2_wr[1967]),  .coef_in(coef[700]), .rdup_out(a3_wr[1711]), .rdlo_out(a3_wr[1967]));
			radix2 #(.width(width)) rd_st2_1712  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1712]), .rdlo_in(a2_wr[1968]),  .coef_in(coef[704]), .rdup_out(a3_wr[1712]), .rdlo_out(a3_wr[1968]));
			radix2 #(.width(width)) rd_st2_1713  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1713]), .rdlo_in(a2_wr[1969]),  .coef_in(coef[708]), .rdup_out(a3_wr[1713]), .rdlo_out(a3_wr[1969]));
			radix2 #(.width(width)) rd_st2_1714  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1714]), .rdlo_in(a2_wr[1970]),  .coef_in(coef[712]), .rdup_out(a3_wr[1714]), .rdlo_out(a3_wr[1970]));
			radix2 #(.width(width)) rd_st2_1715  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1715]), .rdlo_in(a2_wr[1971]),  .coef_in(coef[716]), .rdup_out(a3_wr[1715]), .rdlo_out(a3_wr[1971]));
			radix2 #(.width(width)) rd_st2_1716  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1716]), .rdlo_in(a2_wr[1972]),  .coef_in(coef[720]), .rdup_out(a3_wr[1716]), .rdlo_out(a3_wr[1972]));
			radix2 #(.width(width)) rd_st2_1717  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1717]), .rdlo_in(a2_wr[1973]),  .coef_in(coef[724]), .rdup_out(a3_wr[1717]), .rdlo_out(a3_wr[1973]));
			radix2 #(.width(width)) rd_st2_1718  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1718]), .rdlo_in(a2_wr[1974]),  .coef_in(coef[728]), .rdup_out(a3_wr[1718]), .rdlo_out(a3_wr[1974]));
			radix2 #(.width(width)) rd_st2_1719  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1719]), .rdlo_in(a2_wr[1975]),  .coef_in(coef[732]), .rdup_out(a3_wr[1719]), .rdlo_out(a3_wr[1975]));
			radix2 #(.width(width)) rd_st2_1720  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1720]), .rdlo_in(a2_wr[1976]),  .coef_in(coef[736]), .rdup_out(a3_wr[1720]), .rdlo_out(a3_wr[1976]));
			radix2 #(.width(width)) rd_st2_1721  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1721]), .rdlo_in(a2_wr[1977]),  .coef_in(coef[740]), .rdup_out(a3_wr[1721]), .rdlo_out(a3_wr[1977]));
			radix2 #(.width(width)) rd_st2_1722  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1722]), .rdlo_in(a2_wr[1978]),  .coef_in(coef[744]), .rdup_out(a3_wr[1722]), .rdlo_out(a3_wr[1978]));
			radix2 #(.width(width)) rd_st2_1723  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1723]), .rdlo_in(a2_wr[1979]),  .coef_in(coef[748]), .rdup_out(a3_wr[1723]), .rdlo_out(a3_wr[1979]));
			radix2 #(.width(width)) rd_st2_1724  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1724]), .rdlo_in(a2_wr[1980]),  .coef_in(coef[752]), .rdup_out(a3_wr[1724]), .rdlo_out(a3_wr[1980]));
			radix2 #(.width(width)) rd_st2_1725  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1725]), .rdlo_in(a2_wr[1981]),  .coef_in(coef[756]), .rdup_out(a3_wr[1725]), .rdlo_out(a3_wr[1981]));
			radix2 #(.width(width)) rd_st2_1726  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1726]), .rdlo_in(a2_wr[1982]),  .coef_in(coef[760]), .rdup_out(a3_wr[1726]), .rdlo_out(a3_wr[1982]));
			radix2 #(.width(width)) rd_st2_1727  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1727]), .rdlo_in(a2_wr[1983]),  .coef_in(coef[764]), .rdup_out(a3_wr[1727]), .rdlo_out(a3_wr[1983]));
			radix2 #(.width(width)) rd_st2_1728  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1728]), .rdlo_in(a2_wr[1984]),  .coef_in(coef[768]), .rdup_out(a3_wr[1728]), .rdlo_out(a3_wr[1984]));
			radix2 #(.width(width)) rd_st2_1729  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1729]), .rdlo_in(a2_wr[1985]),  .coef_in(coef[772]), .rdup_out(a3_wr[1729]), .rdlo_out(a3_wr[1985]));
			radix2 #(.width(width)) rd_st2_1730  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1730]), .rdlo_in(a2_wr[1986]),  .coef_in(coef[776]), .rdup_out(a3_wr[1730]), .rdlo_out(a3_wr[1986]));
			radix2 #(.width(width)) rd_st2_1731  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1731]), .rdlo_in(a2_wr[1987]),  .coef_in(coef[780]), .rdup_out(a3_wr[1731]), .rdlo_out(a3_wr[1987]));
			radix2 #(.width(width)) rd_st2_1732  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1732]), .rdlo_in(a2_wr[1988]),  .coef_in(coef[784]), .rdup_out(a3_wr[1732]), .rdlo_out(a3_wr[1988]));
			radix2 #(.width(width)) rd_st2_1733  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1733]), .rdlo_in(a2_wr[1989]),  .coef_in(coef[788]), .rdup_out(a3_wr[1733]), .rdlo_out(a3_wr[1989]));
			radix2 #(.width(width)) rd_st2_1734  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1734]), .rdlo_in(a2_wr[1990]),  .coef_in(coef[792]), .rdup_out(a3_wr[1734]), .rdlo_out(a3_wr[1990]));
			radix2 #(.width(width)) rd_st2_1735  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1735]), .rdlo_in(a2_wr[1991]),  .coef_in(coef[796]), .rdup_out(a3_wr[1735]), .rdlo_out(a3_wr[1991]));
			radix2 #(.width(width)) rd_st2_1736  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1736]), .rdlo_in(a2_wr[1992]),  .coef_in(coef[800]), .rdup_out(a3_wr[1736]), .rdlo_out(a3_wr[1992]));
			radix2 #(.width(width)) rd_st2_1737  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1737]), .rdlo_in(a2_wr[1993]),  .coef_in(coef[804]), .rdup_out(a3_wr[1737]), .rdlo_out(a3_wr[1993]));
			radix2 #(.width(width)) rd_st2_1738  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1738]), .rdlo_in(a2_wr[1994]),  .coef_in(coef[808]), .rdup_out(a3_wr[1738]), .rdlo_out(a3_wr[1994]));
			radix2 #(.width(width)) rd_st2_1739  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1739]), .rdlo_in(a2_wr[1995]),  .coef_in(coef[812]), .rdup_out(a3_wr[1739]), .rdlo_out(a3_wr[1995]));
			radix2 #(.width(width)) rd_st2_1740  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1740]), .rdlo_in(a2_wr[1996]),  .coef_in(coef[816]), .rdup_out(a3_wr[1740]), .rdlo_out(a3_wr[1996]));
			radix2 #(.width(width)) rd_st2_1741  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1741]), .rdlo_in(a2_wr[1997]),  .coef_in(coef[820]), .rdup_out(a3_wr[1741]), .rdlo_out(a3_wr[1997]));
			radix2 #(.width(width)) rd_st2_1742  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1742]), .rdlo_in(a2_wr[1998]),  .coef_in(coef[824]), .rdup_out(a3_wr[1742]), .rdlo_out(a3_wr[1998]));
			radix2 #(.width(width)) rd_st2_1743  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1743]), .rdlo_in(a2_wr[1999]),  .coef_in(coef[828]), .rdup_out(a3_wr[1743]), .rdlo_out(a3_wr[1999]));
			radix2 #(.width(width)) rd_st2_1744  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1744]), .rdlo_in(a2_wr[2000]),  .coef_in(coef[832]), .rdup_out(a3_wr[1744]), .rdlo_out(a3_wr[2000]));
			radix2 #(.width(width)) rd_st2_1745  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1745]), .rdlo_in(a2_wr[2001]),  .coef_in(coef[836]), .rdup_out(a3_wr[1745]), .rdlo_out(a3_wr[2001]));
			radix2 #(.width(width)) rd_st2_1746  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1746]), .rdlo_in(a2_wr[2002]),  .coef_in(coef[840]), .rdup_out(a3_wr[1746]), .rdlo_out(a3_wr[2002]));
			radix2 #(.width(width)) rd_st2_1747  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1747]), .rdlo_in(a2_wr[2003]),  .coef_in(coef[844]), .rdup_out(a3_wr[1747]), .rdlo_out(a3_wr[2003]));
			radix2 #(.width(width)) rd_st2_1748  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1748]), .rdlo_in(a2_wr[2004]),  .coef_in(coef[848]), .rdup_out(a3_wr[1748]), .rdlo_out(a3_wr[2004]));
			radix2 #(.width(width)) rd_st2_1749  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1749]), .rdlo_in(a2_wr[2005]),  .coef_in(coef[852]), .rdup_out(a3_wr[1749]), .rdlo_out(a3_wr[2005]));
			radix2 #(.width(width)) rd_st2_1750  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1750]), .rdlo_in(a2_wr[2006]),  .coef_in(coef[856]), .rdup_out(a3_wr[1750]), .rdlo_out(a3_wr[2006]));
			radix2 #(.width(width)) rd_st2_1751  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1751]), .rdlo_in(a2_wr[2007]),  .coef_in(coef[860]), .rdup_out(a3_wr[1751]), .rdlo_out(a3_wr[2007]));
			radix2 #(.width(width)) rd_st2_1752  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1752]), .rdlo_in(a2_wr[2008]),  .coef_in(coef[864]), .rdup_out(a3_wr[1752]), .rdlo_out(a3_wr[2008]));
			radix2 #(.width(width)) rd_st2_1753  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1753]), .rdlo_in(a2_wr[2009]),  .coef_in(coef[868]), .rdup_out(a3_wr[1753]), .rdlo_out(a3_wr[2009]));
			radix2 #(.width(width)) rd_st2_1754  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1754]), .rdlo_in(a2_wr[2010]),  .coef_in(coef[872]), .rdup_out(a3_wr[1754]), .rdlo_out(a3_wr[2010]));
			radix2 #(.width(width)) rd_st2_1755  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1755]), .rdlo_in(a2_wr[2011]),  .coef_in(coef[876]), .rdup_out(a3_wr[1755]), .rdlo_out(a3_wr[2011]));
			radix2 #(.width(width)) rd_st2_1756  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1756]), .rdlo_in(a2_wr[2012]),  .coef_in(coef[880]), .rdup_out(a3_wr[1756]), .rdlo_out(a3_wr[2012]));
			radix2 #(.width(width)) rd_st2_1757  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1757]), .rdlo_in(a2_wr[2013]),  .coef_in(coef[884]), .rdup_out(a3_wr[1757]), .rdlo_out(a3_wr[2013]));
			radix2 #(.width(width)) rd_st2_1758  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1758]), .rdlo_in(a2_wr[2014]),  .coef_in(coef[888]), .rdup_out(a3_wr[1758]), .rdlo_out(a3_wr[2014]));
			radix2 #(.width(width)) rd_st2_1759  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1759]), .rdlo_in(a2_wr[2015]),  .coef_in(coef[892]), .rdup_out(a3_wr[1759]), .rdlo_out(a3_wr[2015]));
			radix2 #(.width(width)) rd_st2_1760  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1760]), .rdlo_in(a2_wr[2016]),  .coef_in(coef[896]), .rdup_out(a3_wr[1760]), .rdlo_out(a3_wr[2016]));
			radix2 #(.width(width)) rd_st2_1761  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1761]), .rdlo_in(a2_wr[2017]),  .coef_in(coef[900]), .rdup_out(a3_wr[1761]), .rdlo_out(a3_wr[2017]));
			radix2 #(.width(width)) rd_st2_1762  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1762]), .rdlo_in(a2_wr[2018]),  .coef_in(coef[904]), .rdup_out(a3_wr[1762]), .rdlo_out(a3_wr[2018]));
			radix2 #(.width(width)) rd_st2_1763  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1763]), .rdlo_in(a2_wr[2019]),  .coef_in(coef[908]), .rdup_out(a3_wr[1763]), .rdlo_out(a3_wr[2019]));
			radix2 #(.width(width)) rd_st2_1764  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1764]), .rdlo_in(a2_wr[2020]),  .coef_in(coef[912]), .rdup_out(a3_wr[1764]), .rdlo_out(a3_wr[2020]));
			radix2 #(.width(width)) rd_st2_1765  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1765]), .rdlo_in(a2_wr[2021]),  .coef_in(coef[916]), .rdup_out(a3_wr[1765]), .rdlo_out(a3_wr[2021]));
			radix2 #(.width(width)) rd_st2_1766  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1766]), .rdlo_in(a2_wr[2022]),  .coef_in(coef[920]), .rdup_out(a3_wr[1766]), .rdlo_out(a3_wr[2022]));
			radix2 #(.width(width)) rd_st2_1767  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1767]), .rdlo_in(a2_wr[2023]),  .coef_in(coef[924]), .rdup_out(a3_wr[1767]), .rdlo_out(a3_wr[2023]));
			radix2 #(.width(width)) rd_st2_1768  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1768]), .rdlo_in(a2_wr[2024]),  .coef_in(coef[928]), .rdup_out(a3_wr[1768]), .rdlo_out(a3_wr[2024]));
			radix2 #(.width(width)) rd_st2_1769  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1769]), .rdlo_in(a2_wr[2025]),  .coef_in(coef[932]), .rdup_out(a3_wr[1769]), .rdlo_out(a3_wr[2025]));
			radix2 #(.width(width)) rd_st2_1770  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1770]), .rdlo_in(a2_wr[2026]),  .coef_in(coef[936]), .rdup_out(a3_wr[1770]), .rdlo_out(a3_wr[2026]));
			radix2 #(.width(width)) rd_st2_1771  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1771]), .rdlo_in(a2_wr[2027]),  .coef_in(coef[940]), .rdup_out(a3_wr[1771]), .rdlo_out(a3_wr[2027]));
			radix2 #(.width(width)) rd_st2_1772  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1772]), .rdlo_in(a2_wr[2028]),  .coef_in(coef[944]), .rdup_out(a3_wr[1772]), .rdlo_out(a3_wr[2028]));
			radix2 #(.width(width)) rd_st2_1773  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1773]), .rdlo_in(a2_wr[2029]),  .coef_in(coef[948]), .rdup_out(a3_wr[1773]), .rdlo_out(a3_wr[2029]));
			radix2 #(.width(width)) rd_st2_1774  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1774]), .rdlo_in(a2_wr[2030]),  .coef_in(coef[952]), .rdup_out(a3_wr[1774]), .rdlo_out(a3_wr[2030]));
			radix2 #(.width(width)) rd_st2_1775  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1775]), .rdlo_in(a2_wr[2031]),  .coef_in(coef[956]), .rdup_out(a3_wr[1775]), .rdlo_out(a3_wr[2031]));
			radix2 #(.width(width)) rd_st2_1776  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1776]), .rdlo_in(a2_wr[2032]),  .coef_in(coef[960]), .rdup_out(a3_wr[1776]), .rdlo_out(a3_wr[2032]));
			radix2 #(.width(width)) rd_st2_1777  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1777]), .rdlo_in(a2_wr[2033]),  .coef_in(coef[964]), .rdup_out(a3_wr[1777]), .rdlo_out(a3_wr[2033]));
			radix2 #(.width(width)) rd_st2_1778  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1778]), .rdlo_in(a2_wr[2034]),  .coef_in(coef[968]), .rdup_out(a3_wr[1778]), .rdlo_out(a3_wr[2034]));
			radix2 #(.width(width)) rd_st2_1779  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1779]), .rdlo_in(a2_wr[2035]),  .coef_in(coef[972]), .rdup_out(a3_wr[1779]), .rdlo_out(a3_wr[2035]));
			radix2 #(.width(width)) rd_st2_1780  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1780]), .rdlo_in(a2_wr[2036]),  .coef_in(coef[976]), .rdup_out(a3_wr[1780]), .rdlo_out(a3_wr[2036]));
			radix2 #(.width(width)) rd_st2_1781  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1781]), .rdlo_in(a2_wr[2037]),  .coef_in(coef[980]), .rdup_out(a3_wr[1781]), .rdlo_out(a3_wr[2037]));
			radix2 #(.width(width)) rd_st2_1782  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1782]), .rdlo_in(a2_wr[2038]),  .coef_in(coef[984]), .rdup_out(a3_wr[1782]), .rdlo_out(a3_wr[2038]));
			radix2 #(.width(width)) rd_st2_1783  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1783]), .rdlo_in(a2_wr[2039]),  .coef_in(coef[988]), .rdup_out(a3_wr[1783]), .rdlo_out(a3_wr[2039]));
			radix2 #(.width(width)) rd_st2_1784  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1784]), .rdlo_in(a2_wr[2040]),  .coef_in(coef[992]), .rdup_out(a3_wr[1784]), .rdlo_out(a3_wr[2040]));
			radix2 #(.width(width)) rd_st2_1785  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1785]), .rdlo_in(a2_wr[2041]),  .coef_in(coef[996]), .rdup_out(a3_wr[1785]), .rdlo_out(a3_wr[2041]));
			radix2 #(.width(width)) rd_st2_1786  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1786]), .rdlo_in(a2_wr[2042]),  .coef_in(coef[1000]), .rdup_out(a3_wr[1786]), .rdlo_out(a3_wr[2042]));
			radix2 #(.width(width)) rd_st2_1787  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1787]), .rdlo_in(a2_wr[2043]),  .coef_in(coef[1004]), .rdup_out(a3_wr[1787]), .rdlo_out(a3_wr[2043]));
			radix2 #(.width(width)) rd_st2_1788  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1788]), .rdlo_in(a2_wr[2044]),  .coef_in(coef[1008]), .rdup_out(a3_wr[1788]), .rdlo_out(a3_wr[2044]));
			radix2 #(.width(width)) rd_st2_1789  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1789]), .rdlo_in(a2_wr[2045]),  .coef_in(coef[1012]), .rdup_out(a3_wr[1789]), .rdlo_out(a3_wr[2045]));
			radix2 #(.width(width)) rd_st2_1790  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1790]), .rdlo_in(a2_wr[2046]),  .coef_in(coef[1016]), .rdup_out(a3_wr[1790]), .rdlo_out(a3_wr[2046]));
			radix2 #(.width(width)) rd_st2_1791  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a2_wr[1791]), .rdlo_in(a2_wr[2047]),  .coef_in(coef[1020]), .rdup_out(a3_wr[1791]), .rdlo_out(a3_wr[2047]));

		//--- radix stage 3
			radix2 #(.width(width)) rd_st3_0   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[0]), .rdlo_in(a3_wr[128]),  .coef_in(coef[0]), .rdup_out(a4_wr[0]), .rdlo_out(a4_wr[128]));
			radix2 #(.width(width)) rd_st3_1   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1]), .rdlo_in(a3_wr[129]),  .coef_in(coef[8]), .rdup_out(a4_wr[1]), .rdlo_out(a4_wr[129]));
			radix2 #(.width(width)) rd_st3_2   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[2]), .rdlo_in(a3_wr[130]),  .coef_in(coef[16]), .rdup_out(a4_wr[2]), .rdlo_out(a4_wr[130]));
			radix2 #(.width(width)) rd_st3_3   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[3]), .rdlo_in(a3_wr[131]),  .coef_in(coef[24]), .rdup_out(a4_wr[3]), .rdlo_out(a4_wr[131]));
			radix2 #(.width(width)) rd_st3_4   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[4]), .rdlo_in(a3_wr[132]),  .coef_in(coef[32]), .rdup_out(a4_wr[4]), .rdlo_out(a4_wr[132]));
			radix2 #(.width(width)) rd_st3_5   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[5]), .rdlo_in(a3_wr[133]),  .coef_in(coef[40]), .rdup_out(a4_wr[5]), .rdlo_out(a4_wr[133]));
			radix2 #(.width(width)) rd_st3_6   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[6]), .rdlo_in(a3_wr[134]),  .coef_in(coef[48]), .rdup_out(a4_wr[6]), .rdlo_out(a4_wr[134]));
			radix2 #(.width(width)) rd_st3_7   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[7]), .rdlo_in(a3_wr[135]),  .coef_in(coef[56]), .rdup_out(a4_wr[7]), .rdlo_out(a4_wr[135]));
			radix2 #(.width(width)) rd_st3_8   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[8]), .rdlo_in(a3_wr[136]),  .coef_in(coef[64]), .rdup_out(a4_wr[8]), .rdlo_out(a4_wr[136]));
			radix2 #(.width(width)) rd_st3_9   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[9]), .rdlo_in(a3_wr[137]),  .coef_in(coef[72]), .rdup_out(a4_wr[9]), .rdlo_out(a4_wr[137]));
			radix2 #(.width(width)) rd_st3_10  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[10]), .rdlo_in(a3_wr[138]),  .coef_in(coef[80]), .rdup_out(a4_wr[10]), .rdlo_out(a4_wr[138]));
			radix2 #(.width(width)) rd_st3_11  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[11]), .rdlo_in(a3_wr[139]),  .coef_in(coef[88]), .rdup_out(a4_wr[11]), .rdlo_out(a4_wr[139]));
			radix2 #(.width(width)) rd_st3_12  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[12]), .rdlo_in(a3_wr[140]),  .coef_in(coef[96]), .rdup_out(a4_wr[12]), .rdlo_out(a4_wr[140]));
			radix2 #(.width(width)) rd_st3_13  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[13]), .rdlo_in(a3_wr[141]),  .coef_in(coef[104]), .rdup_out(a4_wr[13]), .rdlo_out(a4_wr[141]));
			radix2 #(.width(width)) rd_st3_14  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[14]), .rdlo_in(a3_wr[142]),  .coef_in(coef[112]), .rdup_out(a4_wr[14]), .rdlo_out(a4_wr[142]));
			radix2 #(.width(width)) rd_st3_15  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[15]), .rdlo_in(a3_wr[143]),  .coef_in(coef[120]), .rdup_out(a4_wr[15]), .rdlo_out(a4_wr[143]));
			radix2 #(.width(width)) rd_st3_16  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[16]), .rdlo_in(a3_wr[144]),  .coef_in(coef[128]), .rdup_out(a4_wr[16]), .rdlo_out(a4_wr[144]));
			radix2 #(.width(width)) rd_st3_17  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[17]), .rdlo_in(a3_wr[145]),  .coef_in(coef[136]), .rdup_out(a4_wr[17]), .rdlo_out(a4_wr[145]));
			radix2 #(.width(width)) rd_st3_18  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[18]), .rdlo_in(a3_wr[146]),  .coef_in(coef[144]), .rdup_out(a4_wr[18]), .rdlo_out(a4_wr[146]));
			radix2 #(.width(width)) rd_st3_19  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[19]), .rdlo_in(a3_wr[147]),  .coef_in(coef[152]), .rdup_out(a4_wr[19]), .rdlo_out(a4_wr[147]));
			radix2 #(.width(width)) rd_st3_20  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[20]), .rdlo_in(a3_wr[148]),  .coef_in(coef[160]), .rdup_out(a4_wr[20]), .rdlo_out(a4_wr[148]));
			radix2 #(.width(width)) rd_st3_21  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[21]), .rdlo_in(a3_wr[149]),  .coef_in(coef[168]), .rdup_out(a4_wr[21]), .rdlo_out(a4_wr[149]));
			radix2 #(.width(width)) rd_st3_22  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[22]), .rdlo_in(a3_wr[150]),  .coef_in(coef[176]), .rdup_out(a4_wr[22]), .rdlo_out(a4_wr[150]));
			radix2 #(.width(width)) rd_st3_23  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[23]), .rdlo_in(a3_wr[151]),  .coef_in(coef[184]), .rdup_out(a4_wr[23]), .rdlo_out(a4_wr[151]));
			radix2 #(.width(width)) rd_st3_24  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[24]), .rdlo_in(a3_wr[152]),  .coef_in(coef[192]), .rdup_out(a4_wr[24]), .rdlo_out(a4_wr[152]));
			radix2 #(.width(width)) rd_st3_25  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[25]), .rdlo_in(a3_wr[153]),  .coef_in(coef[200]), .rdup_out(a4_wr[25]), .rdlo_out(a4_wr[153]));
			radix2 #(.width(width)) rd_st3_26  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[26]), .rdlo_in(a3_wr[154]),  .coef_in(coef[208]), .rdup_out(a4_wr[26]), .rdlo_out(a4_wr[154]));
			radix2 #(.width(width)) rd_st3_27  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[27]), .rdlo_in(a3_wr[155]),  .coef_in(coef[216]), .rdup_out(a4_wr[27]), .rdlo_out(a4_wr[155]));
			radix2 #(.width(width)) rd_st3_28  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[28]), .rdlo_in(a3_wr[156]),  .coef_in(coef[224]), .rdup_out(a4_wr[28]), .rdlo_out(a4_wr[156]));
			radix2 #(.width(width)) rd_st3_29  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[29]), .rdlo_in(a3_wr[157]),  .coef_in(coef[232]), .rdup_out(a4_wr[29]), .rdlo_out(a4_wr[157]));
			radix2 #(.width(width)) rd_st3_30  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[30]), .rdlo_in(a3_wr[158]),  .coef_in(coef[240]), .rdup_out(a4_wr[30]), .rdlo_out(a4_wr[158]));
			radix2 #(.width(width)) rd_st3_31  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[31]), .rdlo_in(a3_wr[159]),  .coef_in(coef[248]), .rdup_out(a4_wr[31]), .rdlo_out(a4_wr[159]));
			radix2 #(.width(width)) rd_st3_32  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[32]), .rdlo_in(a3_wr[160]),  .coef_in(coef[256]), .rdup_out(a4_wr[32]), .rdlo_out(a4_wr[160]));
			radix2 #(.width(width)) rd_st3_33  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[33]), .rdlo_in(a3_wr[161]),  .coef_in(coef[264]), .rdup_out(a4_wr[33]), .rdlo_out(a4_wr[161]));
			radix2 #(.width(width)) rd_st3_34  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[34]), .rdlo_in(a3_wr[162]),  .coef_in(coef[272]), .rdup_out(a4_wr[34]), .rdlo_out(a4_wr[162]));
			radix2 #(.width(width)) rd_st3_35  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[35]), .rdlo_in(a3_wr[163]),  .coef_in(coef[280]), .rdup_out(a4_wr[35]), .rdlo_out(a4_wr[163]));
			radix2 #(.width(width)) rd_st3_36  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[36]), .rdlo_in(a3_wr[164]),  .coef_in(coef[288]), .rdup_out(a4_wr[36]), .rdlo_out(a4_wr[164]));
			radix2 #(.width(width)) rd_st3_37  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[37]), .rdlo_in(a3_wr[165]),  .coef_in(coef[296]), .rdup_out(a4_wr[37]), .rdlo_out(a4_wr[165]));
			radix2 #(.width(width)) rd_st3_38  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[38]), .rdlo_in(a3_wr[166]),  .coef_in(coef[304]), .rdup_out(a4_wr[38]), .rdlo_out(a4_wr[166]));
			radix2 #(.width(width)) rd_st3_39  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[39]), .rdlo_in(a3_wr[167]),  .coef_in(coef[312]), .rdup_out(a4_wr[39]), .rdlo_out(a4_wr[167]));
			radix2 #(.width(width)) rd_st3_40  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[40]), .rdlo_in(a3_wr[168]),  .coef_in(coef[320]), .rdup_out(a4_wr[40]), .rdlo_out(a4_wr[168]));
			radix2 #(.width(width)) rd_st3_41  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[41]), .rdlo_in(a3_wr[169]),  .coef_in(coef[328]), .rdup_out(a4_wr[41]), .rdlo_out(a4_wr[169]));
			radix2 #(.width(width)) rd_st3_42  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[42]), .rdlo_in(a3_wr[170]),  .coef_in(coef[336]), .rdup_out(a4_wr[42]), .rdlo_out(a4_wr[170]));
			radix2 #(.width(width)) rd_st3_43  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[43]), .rdlo_in(a3_wr[171]),  .coef_in(coef[344]), .rdup_out(a4_wr[43]), .rdlo_out(a4_wr[171]));
			radix2 #(.width(width)) rd_st3_44  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[44]), .rdlo_in(a3_wr[172]),  .coef_in(coef[352]), .rdup_out(a4_wr[44]), .rdlo_out(a4_wr[172]));
			radix2 #(.width(width)) rd_st3_45  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[45]), .rdlo_in(a3_wr[173]),  .coef_in(coef[360]), .rdup_out(a4_wr[45]), .rdlo_out(a4_wr[173]));
			radix2 #(.width(width)) rd_st3_46  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[46]), .rdlo_in(a3_wr[174]),  .coef_in(coef[368]), .rdup_out(a4_wr[46]), .rdlo_out(a4_wr[174]));
			radix2 #(.width(width)) rd_st3_47  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[47]), .rdlo_in(a3_wr[175]),  .coef_in(coef[376]), .rdup_out(a4_wr[47]), .rdlo_out(a4_wr[175]));
			radix2 #(.width(width)) rd_st3_48  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[48]), .rdlo_in(a3_wr[176]),  .coef_in(coef[384]), .rdup_out(a4_wr[48]), .rdlo_out(a4_wr[176]));
			radix2 #(.width(width)) rd_st3_49  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[49]), .rdlo_in(a3_wr[177]),  .coef_in(coef[392]), .rdup_out(a4_wr[49]), .rdlo_out(a4_wr[177]));
			radix2 #(.width(width)) rd_st3_50  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[50]), .rdlo_in(a3_wr[178]),  .coef_in(coef[400]), .rdup_out(a4_wr[50]), .rdlo_out(a4_wr[178]));
			radix2 #(.width(width)) rd_st3_51  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[51]), .rdlo_in(a3_wr[179]),  .coef_in(coef[408]), .rdup_out(a4_wr[51]), .rdlo_out(a4_wr[179]));
			radix2 #(.width(width)) rd_st3_52  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[52]), .rdlo_in(a3_wr[180]),  .coef_in(coef[416]), .rdup_out(a4_wr[52]), .rdlo_out(a4_wr[180]));
			radix2 #(.width(width)) rd_st3_53  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[53]), .rdlo_in(a3_wr[181]),  .coef_in(coef[424]), .rdup_out(a4_wr[53]), .rdlo_out(a4_wr[181]));
			radix2 #(.width(width)) rd_st3_54  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[54]), .rdlo_in(a3_wr[182]),  .coef_in(coef[432]), .rdup_out(a4_wr[54]), .rdlo_out(a4_wr[182]));
			radix2 #(.width(width)) rd_st3_55  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[55]), .rdlo_in(a3_wr[183]),  .coef_in(coef[440]), .rdup_out(a4_wr[55]), .rdlo_out(a4_wr[183]));
			radix2 #(.width(width)) rd_st3_56  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[56]), .rdlo_in(a3_wr[184]),  .coef_in(coef[448]), .rdup_out(a4_wr[56]), .rdlo_out(a4_wr[184]));
			radix2 #(.width(width)) rd_st3_57  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[57]), .rdlo_in(a3_wr[185]),  .coef_in(coef[456]), .rdup_out(a4_wr[57]), .rdlo_out(a4_wr[185]));
			radix2 #(.width(width)) rd_st3_58  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[58]), .rdlo_in(a3_wr[186]),  .coef_in(coef[464]), .rdup_out(a4_wr[58]), .rdlo_out(a4_wr[186]));
			radix2 #(.width(width)) rd_st3_59  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[59]), .rdlo_in(a3_wr[187]),  .coef_in(coef[472]), .rdup_out(a4_wr[59]), .rdlo_out(a4_wr[187]));
			radix2 #(.width(width)) rd_st3_60  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[60]), .rdlo_in(a3_wr[188]),  .coef_in(coef[480]), .rdup_out(a4_wr[60]), .rdlo_out(a4_wr[188]));
			radix2 #(.width(width)) rd_st3_61  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[61]), .rdlo_in(a3_wr[189]),  .coef_in(coef[488]), .rdup_out(a4_wr[61]), .rdlo_out(a4_wr[189]));
			radix2 #(.width(width)) rd_st3_62  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[62]), .rdlo_in(a3_wr[190]),  .coef_in(coef[496]), .rdup_out(a4_wr[62]), .rdlo_out(a4_wr[190]));
			radix2 #(.width(width)) rd_st3_63  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[63]), .rdlo_in(a3_wr[191]),  .coef_in(coef[504]), .rdup_out(a4_wr[63]), .rdlo_out(a4_wr[191]));
			radix2 #(.width(width)) rd_st3_64  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[64]), .rdlo_in(a3_wr[192]),  .coef_in(coef[512]), .rdup_out(a4_wr[64]), .rdlo_out(a4_wr[192]));
			radix2 #(.width(width)) rd_st3_65  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[65]), .rdlo_in(a3_wr[193]),  .coef_in(coef[520]), .rdup_out(a4_wr[65]), .rdlo_out(a4_wr[193]));
			radix2 #(.width(width)) rd_st3_66  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[66]), .rdlo_in(a3_wr[194]),  .coef_in(coef[528]), .rdup_out(a4_wr[66]), .rdlo_out(a4_wr[194]));
			radix2 #(.width(width)) rd_st3_67  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[67]), .rdlo_in(a3_wr[195]),  .coef_in(coef[536]), .rdup_out(a4_wr[67]), .rdlo_out(a4_wr[195]));
			radix2 #(.width(width)) rd_st3_68  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[68]), .rdlo_in(a3_wr[196]),  .coef_in(coef[544]), .rdup_out(a4_wr[68]), .rdlo_out(a4_wr[196]));
			radix2 #(.width(width)) rd_st3_69  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[69]), .rdlo_in(a3_wr[197]),  .coef_in(coef[552]), .rdup_out(a4_wr[69]), .rdlo_out(a4_wr[197]));
			radix2 #(.width(width)) rd_st3_70  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[70]), .rdlo_in(a3_wr[198]),  .coef_in(coef[560]), .rdup_out(a4_wr[70]), .rdlo_out(a4_wr[198]));
			radix2 #(.width(width)) rd_st3_71  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[71]), .rdlo_in(a3_wr[199]),  .coef_in(coef[568]), .rdup_out(a4_wr[71]), .rdlo_out(a4_wr[199]));
			radix2 #(.width(width)) rd_st3_72  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[72]), .rdlo_in(a3_wr[200]),  .coef_in(coef[576]), .rdup_out(a4_wr[72]), .rdlo_out(a4_wr[200]));
			radix2 #(.width(width)) rd_st3_73  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[73]), .rdlo_in(a3_wr[201]),  .coef_in(coef[584]), .rdup_out(a4_wr[73]), .rdlo_out(a4_wr[201]));
			radix2 #(.width(width)) rd_st3_74  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[74]), .rdlo_in(a3_wr[202]),  .coef_in(coef[592]), .rdup_out(a4_wr[74]), .rdlo_out(a4_wr[202]));
			radix2 #(.width(width)) rd_st3_75  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[75]), .rdlo_in(a3_wr[203]),  .coef_in(coef[600]), .rdup_out(a4_wr[75]), .rdlo_out(a4_wr[203]));
			radix2 #(.width(width)) rd_st3_76  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[76]), .rdlo_in(a3_wr[204]),  .coef_in(coef[608]), .rdup_out(a4_wr[76]), .rdlo_out(a4_wr[204]));
			radix2 #(.width(width)) rd_st3_77  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[77]), .rdlo_in(a3_wr[205]),  .coef_in(coef[616]), .rdup_out(a4_wr[77]), .rdlo_out(a4_wr[205]));
			radix2 #(.width(width)) rd_st3_78  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[78]), .rdlo_in(a3_wr[206]),  .coef_in(coef[624]), .rdup_out(a4_wr[78]), .rdlo_out(a4_wr[206]));
			radix2 #(.width(width)) rd_st3_79  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[79]), .rdlo_in(a3_wr[207]),  .coef_in(coef[632]), .rdup_out(a4_wr[79]), .rdlo_out(a4_wr[207]));
			radix2 #(.width(width)) rd_st3_80  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[80]), .rdlo_in(a3_wr[208]),  .coef_in(coef[640]), .rdup_out(a4_wr[80]), .rdlo_out(a4_wr[208]));
			radix2 #(.width(width)) rd_st3_81  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[81]), .rdlo_in(a3_wr[209]),  .coef_in(coef[648]), .rdup_out(a4_wr[81]), .rdlo_out(a4_wr[209]));
			radix2 #(.width(width)) rd_st3_82  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[82]), .rdlo_in(a3_wr[210]),  .coef_in(coef[656]), .rdup_out(a4_wr[82]), .rdlo_out(a4_wr[210]));
			radix2 #(.width(width)) rd_st3_83  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[83]), .rdlo_in(a3_wr[211]),  .coef_in(coef[664]), .rdup_out(a4_wr[83]), .rdlo_out(a4_wr[211]));
			radix2 #(.width(width)) rd_st3_84  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[84]), .rdlo_in(a3_wr[212]),  .coef_in(coef[672]), .rdup_out(a4_wr[84]), .rdlo_out(a4_wr[212]));
			radix2 #(.width(width)) rd_st3_85  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[85]), .rdlo_in(a3_wr[213]),  .coef_in(coef[680]), .rdup_out(a4_wr[85]), .rdlo_out(a4_wr[213]));
			radix2 #(.width(width)) rd_st3_86  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[86]), .rdlo_in(a3_wr[214]),  .coef_in(coef[688]), .rdup_out(a4_wr[86]), .rdlo_out(a4_wr[214]));
			radix2 #(.width(width)) rd_st3_87  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[87]), .rdlo_in(a3_wr[215]),  .coef_in(coef[696]), .rdup_out(a4_wr[87]), .rdlo_out(a4_wr[215]));
			radix2 #(.width(width)) rd_st3_88  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[88]), .rdlo_in(a3_wr[216]),  .coef_in(coef[704]), .rdup_out(a4_wr[88]), .rdlo_out(a4_wr[216]));
			radix2 #(.width(width)) rd_st3_89  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[89]), .rdlo_in(a3_wr[217]),  .coef_in(coef[712]), .rdup_out(a4_wr[89]), .rdlo_out(a4_wr[217]));
			radix2 #(.width(width)) rd_st3_90  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[90]), .rdlo_in(a3_wr[218]),  .coef_in(coef[720]), .rdup_out(a4_wr[90]), .rdlo_out(a4_wr[218]));
			radix2 #(.width(width)) rd_st3_91  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[91]), .rdlo_in(a3_wr[219]),  .coef_in(coef[728]), .rdup_out(a4_wr[91]), .rdlo_out(a4_wr[219]));
			radix2 #(.width(width)) rd_st3_92  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[92]), .rdlo_in(a3_wr[220]),  .coef_in(coef[736]), .rdup_out(a4_wr[92]), .rdlo_out(a4_wr[220]));
			radix2 #(.width(width)) rd_st3_93  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[93]), .rdlo_in(a3_wr[221]),  .coef_in(coef[744]), .rdup_out(a4_wr[93]), .rdlo_out(a4_wr[221]));
			radix2 #(.width(width)) rd_st3_94  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[94]), .rdlo_in(a3_wr[222]),  .coef_in(coef[752]), .rdup_out(a4_wr[94]), .rdlo_out(a4_wr[222]));
			radix2 #(.width(width)) rd_st3_95  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[95]), .rdlo_in(a3_wr[223]),  .coef_in(coef[760]), .rdup_out(a4_wr[95]), .rdlo_out(a4_wr[223]));
			radix2 #(.width(width)) rd_st3_96  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[96]), .rdlo_in(a3_wr[224]),  .coef_in(coef[768]), .rdup_out(a4_wr[96]), .rdlo_out(a4_wr[224]));
			radix2 #(.width(width)) rd_st3_97  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[97]), .rdlo_in(a3_wr[225]),  .coef_in(coef[776]), .rdup_out(a4_wr[97]), .rdlo_out(a4_wr[225]));
			radix2 #(.width(width)) rd_st3_98  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[98]), .rdlo_in(a3_wr[226]),  .coef_in(coef[784]), .rdup_out(a4_wr[98]), .rdlo_out(a4_wr[226]));
			radix2 #(.width(width)) rd_st3_99  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[99]), .rdlo_in(a3_wr[227]),  .coef_in(coef[792]), .rdup_out(a4_wr[99]), .rdlo_out(a4_wr[227]));
			radix2 #(.width(width)) rd_st3_100  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[100]), .rdlo_in(a3_wr[228]),  .coef_in(coef[800]), .rdup_out(a4_wr[100]), .rdlo_out(a4_wr[228]));
			radix2 #(.width(width)) rd_st3_101  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[101]), .rdlo_in(a3_wr[229]),  .coef_in(coef[808]), .rdup_out(a4_wr[101]), .rdlo_out(a4_wr[229]));
			radix2 #(.width(width)) rd_st3_102  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[102]), .rdlo_in(a3_wr[230]),  .coef_in(coef[816]), .rdup_out(a4_wr[102]), .rdlo_out(a4_wr[230]));
			radix2 #(.width(width)) rd_st3_103  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[103]), .rdlo_in(a3_wr[231]),  .coef_in(coef[824]), .rdup_out(a4_wr[103]), .rdlo_out(a4_wr[231]));
			radix2 #(.width(width)) rd_st3_104  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[104]), .rdlo_in(a3_wr[232]),  .coef_in(coef[832]), .rdup_out(a4_wr[104]), .rdlo_out(a4_wr[232]));
			radix2 #(.width(width)) rd_st3_105  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[105]), .rdlo_in(a3_wr[233]),  .coef_in(coef[840]), .rdup_out(a4_wr[105]), .rdlo_out(a4_wr[233]));
			radix2 #(.width(width)) rd_st3_106  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[106]), .rdlo_in(a3_wr[234]),  .coef_in(coef[848]), .rdup_out(a4_wr[106]), .rdlo_out(a4_wr[234]));
			radix2 #(.width(width)) rd_st3_107  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[107]), .rdlo_in(a3_wr[235]),  .coef_in(coef[856]), .rdup_out(a4_wr[107]), .rdlo_out(a4_wr[235]));
			radix2 #(.width(width)) rd_st3_108  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[108]), .rdlo_in(a3_wr[236]),  .coef_in(coef[864]), .rdup_out(a4_wr[108]), .rdlo_out(a4_wr[236]));
			radix2 #(.width(width)) rd_st3_109  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[109]), .rdlo_in(a3_wr[237]),  .coef_in(coef[872]), .rdup_out(a4_wr[109]), .rdlo_out(a4_wr[237]));
			radix2 #(.width(width)) rd_st3_110  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[110]), .rdlo_in(a3_wr[238]),  .coef_in(coef[880]), .rdup_out(a4_wr[110]), .rdlo_out(a4_wr[238]));
			radix2 #(.width(width)) rd_st3_111  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[111]), .rdlo_in(a3_wr[239]),  .coef_in(coef[888]), .rdup_out(a4_wr[111]), .rdlo_out(a4_wr[239]));
			radix2 #(.width(width)) rd_st3_112  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[112]), .rdlo_in(a3_wr[240]),  .coef_in(coef[896]), .rdup_out(a4_wr[112]), .rdlo_out(a4_wr[240]));
			radix2 #(.width(width)) rd_st3_113  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[113]), .rdlo_in(a3_wr[241]),  .coef_in(coef[904]), .rdup_out(a4_wr[113]), .rdlo_out(a4_wr[241]));
			radix2 #(.width(width)) rd_st3_114  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[114]), .rdlo_in(a3_wr[242]),  .coef_in(coef[912]), .rdup_out(a4_wr[114]), .rdlo_out(a4_wr[242]));
			radix2 #(.width(width)) rd_st3_115  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[115]), .rdlo_in(a3_wr[243]),  .coef_in(coef[920]), .rdup_out(a4_wr[115]), .rdlo_out(a4_wr[243]));
			radix2 #(.width(width)) rd_st3_116  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[116]), .rdlo_in(a3_wr[244]),  .coef_in(coef[928]), .rdup_out(a4_wr[116]), .rdlo_out(a4_wr[244]));
			radix2 #(.width(width)) rd_st3_117  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[117]), .rdlo_in(a3_wr[245]),  .coef_in(coef[936]), .rdup_out(a4_wr[117]), .rdlo_out(a4_wr[245]));
			radix2 #(.width(width)) rd_st3_118  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[118]), .rdlo_in(a3_wr[246]),  .coef_in(coef[944]), .rdup_out(a4_wr[118]), .rdlo_out(a4_wr[246]));
			radix2 #(.width(width)) rd_st3_119  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[119]), .rdlo_in(a3_wr[247]),  .coef_in(coef[952]), .rdup_out(a4_wr[119]), .rdlo_out(a4_wr[247]));
			radix2 #(.width(width)) rd_st3_120  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[120]), .rdlo_in(a3_wr[248]),  .coef_in(coef[960]), .rdup_out(a4_wr[120]), .rdlo_out(a4_wr[248]));
			radix2 #(.width(width)) rd_st3_121  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[121]), .rdlo_in(a3_wr[249]),  .coef_in(coef[968]), .rdup_out(a4_wr[121]), .rdlo_out(a4_wr[249]));
			radix2 #(.width(width)) rd_st3_122  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[122]), .rdlo_in(a3_wr[250]),  .coef_in(coef[976]), .rdup_out(a4_wr[122]), .rdlo_out(a4_wr[250]));
			radix2 #(.width(width)) rd_st3_123  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[123]), .rdlo_in(a3_wr[251]),  .coef_in(coef[984]), .rdup_out(a4_wr[123]), .rdlo_out(a4_wr[251]));
			radix2 #(.width(width)) rd_st3_124  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[124]), .rdlo_in(a3_wr[252]),  .coef_in(coef[992]), .rdup_out(a4_wr[124]), .rdlo_out(a4_wr[252]));
			radix2 #(.width(width)) rd_st3_125  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[125]), .rdlo_in(a3_wr[253]),  .coef_in(coef[1000]), .rdup_out(a4_wr[125]), .rdlo_out(a4_wr[253]));
			radix2 #(.width(width)) rd_st3_126  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[126]), .rdlo_in(a3_wr[254]),  .coef_in(coef[1008]), .rdup_out(a4_wr[126]), .rdlo_out(a4_wr[254]));
			radix2 #(.width(width)) rd_st3_127  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[127]), .rdlo_in(a3_wr[255]),  .coef_in(coef[1016]), .rdup_out(a4_wr[127]), .rdlo_out(a4_wr[255]));
			radix2 #(.width(width)) rd_st3_256  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[256]), .rdlo_in(a3_wr[384]),  .coef_in(coef[0]), .rdup_out(a4_wr[256]), .rdlo_out(a4_wr[384]));
			radix2 #(.width(width)) rd_st3_257  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[257]), .rdlo_in(a3_wr[385]),  .coef_in(coef[8]), .rdup_out(a4_wr[257]), .rdlo_out(a4_wr[385]));
			radix2 #(.width(width)) rd_st3_258  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[258]), .rdlo_in(a3_wr[386]),  .coef_in(coef[16]), .rdup_out(a4_wr[258]), .rdlo_out(a4_wr[386]));
			radix2 #(.width(width)) rd_st3_259  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[259]), .rdlo_in(a3_wr[387]),  .coef_in(coef[24]), .rdup_out(a4_wr[259]), .rdlo_out(a4_wr[387]));
			radix2 #(.width(width)) rd_st3_260  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[260]), .rdlo_in(a3_wr[388]),  .coef_in(coef[32]), .rdup_out(a4_wr[260]), .rdlo_out(a4_wr[388]));
			radix2 #(.width(width)) rd_st3_261  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[261]), .rdlo_in(a3_wr[389]),  .coef_in(coef[40]), .rdup_out(a4_wr[261]), .rdlo_out(a4_wr[389]));
			radix2 #(.width(width)) rd_st3_262  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[262]), .rdlo_in(a3_wr[390]),  .coef_in(coef[48]), .rdup_out(a4_wr[262]), .rdlo_out(a4_wr[390]));
			radix2 #(.width(width)) rd_st3_263  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[263]), .rdlo_in(a3_wr[391]),  .coef_in(coef[56]), .rdup_out(a4_wr[263]), .rdlo_out(a4_wr[391]));
			radix2 #(.width(width)) rd_st3_264  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[264]), .rdlo_in(a3_wr[392]),  .coef_in(coef[64]), .rdup_out(a4_wr[264]), .rdlo_out(a4_wr[392]));
			radix2 #(.width(width)) rd_st3_265  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[265]), .rdlo_in(a3_wr[393]),  .coef_in(coef[72]), .rdup_out(a4_wr[265]), .rdlo_out(a4_wr[393]));
			radix2 #(.width(width)) rd_st3_266  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[266]), .rdlo_in(a3_wr[394]),  .coef_in(coef[80]), .rdup_out(a4_wr[266]), .rdlo_out(a4_wr[394]));
			radix2 #(.width(width)) rd_st3_267  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[267]), .rdlo_in(a3_wr[395]),  .coef_in(coef[88]), .rdup_out(a4_wr[267]), .rdlo_out(a4_wr[395]));
			radix2 #(.width(width)) rd_st3_268  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[268]), .rdlo_in(a3_wr[396]),  .coef_in(coef[96]), .rdup_out(a4_wr[268]), .rdlo_out(a4_wr[396]));
			radix2 #(.width(width)) rd_st3_269  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[269]), .rdlo_in(a3_wr[397]),  .coef_in(coef[104]), .rdup_out(a4_wr[269]), .rdlo_out(a4_wr[397]));
			radix2 #(.width(width)) rd_st3_270  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[270]), .rdlo_in(a3_wr[398]),  .coef_in(coef[112]), .rdup_out(a4_wr[270]), .rdlo_out(a4_wr[398]));
			radix2 #(.width(width)) rd_st3_271  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[271]), .rdlo_in(a3_wr[399]),  .coef_in(coef[120]), .rdup_out(a4_wr[271]), .rdlo_out(a4_wr[399]));
			radix2 #(.width(width)) rd_st3_272  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[272]), .rdlo_in(a3_wr[400]),  .coef_in(coef[128]), .rdup_out(a4_wr[272]), .rdlo_out(a4_wr[400]));
			radix2 #(.width(width)) rd_st3_273  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[273]), .rdlo_in(a3_wr[401]),  .coef_in(coef[136]), .rdup_out(a4_wr[273]), .rdlo_out(a4_wr[401]));
			radix2 #(.width(width)) rd_st3_274  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[274]), .rdlo_in(a3_wr[402]),  .coef_in(coef[144]), .rdup_out(a4_wr[274]), .rdlo_out(a4_wr[402]));
			radix2 #(.width(width)) rd_st3_275  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[275]), .rdlo_in(a3_wr[403]),  .coef_in(coef[152]), .rdup_out(a4_wr[275]), .rdlo_out(a4_wr[403]));
			radix2 #(.width(width)) rd_st3_276  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[276]), .rdlo_in(a3_wr[404]),  .coef_in(coef[160]), .rdup_out(a4_wr[276]), .rdlo_out(a4_wr[404]));
			radix2 #(.width(width)) rd_st3_277  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[277]), .rdlo_in(a3_wr[405]),  .coef_in(coef[168]), .rdup_out(a4_wr[277]), .rdlo_out(a4_wr[405]));
			radix2 #(.width(width)) rd_st3_278  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[278]), .rdlo_in(a3_wr[406]),  .coef_in(coef[176]), .rdup_out(a4_wr[278]), .rdlo_out(a4_wr[406]));
			radix2 #(.width(width)) rd_st3_279  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[279]), .rdlo_in(a3_wr[407]),  .coef_in(coef[184]), .rdup_out(a4_wr[279]), .rdlo_out(a4_wr[407]));
			radix2 #(.width(width)) rd_st3_280  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[280]), .rdlo_in(a3_wr[408]),  .coef_in(coef[192]), .rdup_out(a4_wr[280]), .rdlo_out(a4_wr[408]));
			radix2 #(.width(width)) rd_st3_281  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[281]), .rdlo_in(a3_wr[409]),  .coef_in(coef[200]), .rdup_out(a4_wr[281]), .rdlo_out(a4_wr[409]));
			radix2 #(.width(width)) rd_st3_282  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[282]), .rdlo_in(a3_wr[410]),  .coef_in(coef[208]), .rdup_out(a4_wr[282]), .rdlo_out(a4_wr[410]));
			radix2 #(.width(width)) rd_st3_283  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[283]), .rdlo_in(a3_wr[411]),  .coef_in(coef[216]), .rdup_out(a4_wr[283]), .rdlo_out(a4_wr[411]));
			radix2 #(.width(width)) rd_st3_284  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[284]), .rdlo_in(a3_wr[412]),  .coef_in(coef[224]), .rdup_out(a4_wr[284]), .rdlo_out(a4_wr[412]));
			radix2 #(.width(width)) rd_st3_285  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[285]), .rdlo_in(a3_wr[413]),  .coef_in(coef[232]), .rdup_out(a4_wr[285]), .rdlo_out(a4_wr[413]));
			radix2 #(.width(width)) rd_st3_286  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[286]), .rdlo_in(a3_wr[414]),  .coef_in(coef[240]), .rdup_out(a4_wr[286]), .rdlo_out(a4_wr[414]));
			radix2 #(.width(width)) rd_st3_287  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[287]), .rdlo_in(a3_wr[415]),  .coef_in(coef[248]), .rdup_out(a4_wr[287]), .rdlo_out(a4_wr[415]));
			radix2 #(.width(width)) rd_st3_288  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[288]), .rdlo_in(a3_wr[416]),  .coef_in(coef[256]), .rdup_out(a4_wr[288]), .rdlo_out(a4_wr[416]));
			radix2 #(.width(width)) rd_st3_289  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[289]), .rdlo_in(a3_wr[417]),  .coef_in(coef[264]), .rdup_out(a4_wr[289]), .rdlo_out(a4_wr[417]));
			radix2 #(.width(width)) rd_st3_290  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[290]), .rdlo_in(a3_wr[418]),  .coef_in(coef[272]), .rdup_out(a4_wr[290]), .rdlo_out(a4_wr[418]));
			radix2 #(.width(width)) rd_st3_291  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[291]), .rdlo_in(a3_wr[419]),  .coef_in(coef[280]), .rdup_out(a4_wr[291]), .rdlo_out(a4_wr[419]));
			radix2 #(.width(width)) rd_st3_292  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[292]), .rdlo_in(a3_wr[420]),  .coef_in(coef[288]), .rdup_out(a4_wr[292]), .rdlo_out(a4_wr[420]));
			radix2 #(.width(width)) rd_st3_293  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[293]), .rdlo_in(a3_wr[421]),  .coef_in(coef[296]), .rdup_out(a4_wr[293]), .rdlo_out(a4_wr[421]));
			radix2 #(.width(width)) rd_st3_294  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[294]), .rdlo_in(a3_wr[422]),  .coef_in(coef[304]), .rdup_out(a4_wr[294]), .rdlo_out(a4_wr[422]));
			radix2 #(.width(width)) rd_st3_295  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[295]), .rdlo_in(a3_wr[423]),  .coef_in(coef[312]), .rdup_out(a4_wr[295]), .rdlo_out(a4_wr[423]));
			radix2 #(.width(width)) rd_st3_296  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[296]), .rdlo_in(a3_wr[424]),  .coef_in(coef[320]), .rdup_out(a4_wr[296]), .rdlo_out(a4_wr[424]));
			radix2 #(.width(width)) rd_st3_297  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[297]), .rdlo_in(a3_wr[425]),  .coef_in(coef[328]), .rdup_out(a4_wr[297]), .rdlo_out(a4_wr[425]));
			radix2 #(.width(width)) rd_st3_298  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[298]), .rdlo_in(a3_wr[426]),  .coef_in(coef[336]), .rdup_out(a4_wr[298]), .rdlo_out(a4_wr[426]));
			radix2 #(.width(width)) rd_st3_299  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[299]), .rdlo_in(a3_wr[427]),  .coef_in(coef[344]), .rdup_out(a4_wr[299]), .rdlo_out(a4_wr[427]));
			radix2 #(.width(width)) rd_st3_300  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[300]), .rdlo_in(a3_wr[428]),  .coef_in(coef[352]), .rdup_out(a4_wr[300]), .rdlo_out(a4_wr[428]));
			radix2 #(.width(width)) rd_st3_301  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[301]), .rdlo_in(a3_wr[429]),  .coef_in(coef[360]), .rdup_out(a4_wr[301]), .rdlo_out(a4_wr[429]));
			radix2 #(.width(width)) rd_st3_302  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[302]), .rdlo_in(a3_wr[430]),  .coef_in(coef[368]), .rdup_out(a4_wr[302]), .rdlo_out(a4_wr[430]));
			radix2 #(.width(width)) rd_st3_303  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[303]), .rdlo_in(a3_wr[431]),  .coef_in(coef[376]), .rdup_out(a4_wr[303]), .rdlo_out(a4_wr[431]));
			radix2 #(.width(width)) rd_st3_304  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[304]), .rdlo_in(a3_wr[432]),  .coef_in(coef[384]), .rdup_out(a4_wr[304]), .rdlo_out(a4_wr[432]));
			radix2 #(.width(width)) rd_st3_305  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[305]), .rdlo_in(a3_wr[433]),  .coef_in(coef[392]), .rdup_out(a4_wr[305]), .rdlo_out(a4_wr[433]));
			radix2 #(.width(width)) rd_st3_306  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[306]), .rdlo_in(a3_wr[434]),  .coef_in(coef[400]), .rdup_out(a4_wr[306]), .rdlo_out(a4_wr[434]));
			radix2 #(.width(width)) rd_st3_307  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[307]), .rdlo_in(a3_wr[435]),  .coef_in(coef[408]), .rdup_out(a4_wr[307]), .rdlo_out(a4_wr[435]));
			radix2 #(.width(width)) rd_st3_308  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[308]), .rdlo_in(a3_wr[436]),  .coef_in(coef[416]), .rdup_out(a4_wr[308]), .rdlo_out(a4_wr[436]));
			radix2 #(.width(width)) rd_st3_309  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[309]), .rdlo_in(a3_wr[437]),  .coef_in(coef[424]), .rdup_out(a4_wr[309]), .rdlo_out(a4_wr[437]));
			radix2 #(.width(width)) rd_st3_310  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[310]), .rdlo_in(a3_wr[438]),  .coef_in(coef[432]), .rdup_out(a4_wr[310]), .rdlo_out(a4_wr[438]));
			radix2 #(.width(width)) rd_st3_311  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[311]), .rdlo_in(a3_wr[439]),  .coef_in(coef[440]), .rdup_out(a4_wr[311]), .rdlo_out(a4_wr[439]));
			radix2 #(.width(width)) rd_st3_312  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[312]), .rdlo_in(a3_wr[440]),  .coef_in(coef[448]), .rdup_out(a4_wr[312]), .rdlo_out(a4_wr[440]));
			radix2 #(.width(width)) rd_st3_313  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[313]), .rdlo_in(a3_wr[441]),  .coef_in(coef[456]), .rdup_out(a4_wr[313]), .rdlo_out(a4_wr[441]));
			radix2 #(.width(width)) rd_st3_314  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[314]), .rdlo_in(a3_wr[442]),  .coef_in(coef[464]), .rdup_out(a4_wr[314]), .rdlo_out(a4_wr[442]));
			radix2 #(.width(width)) rd_st3_315  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[315]), .rdlo_in(a3_wr[443]),  .coef_in(coef[472]), .rdup_out(a4_wr[315]), .rdlo_out(a4_wr[443]));
			radix2 #(.width(width)) rd_st3_316  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[316]), .rdlo_in(a3_wr[444]),  .coef_in(coef[480]), .rdup_out(a4_wr[316]), .rdlo_out(a4_wr[444]));
			radix2 #(.width(width)) rd_st3_317  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[317]), .rdlo_in(a3_wr[445]),  .coef_in(coef[488]), .rdup_out(a4_wr[317]), .rdlo_out(a4_wr[445]));
			radix2 #(.width(width)) rd_st3_318  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[318]), .rdlo_in(a3_wr[446]),  .coef_in(coef[496]), .rdup_out(a4_wr[318]), .rdlo_out(a4_wr[446]));
			radix2 #(.width(width)) rd_st3_319  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[319]), .rdlo_in(a3_wr[447]),  .coef_in(coef[504]), .rdup_out(a4_wr[319]), .rdlo_out(a4_wr[447]));
			radix2 #(.width(width)) rd_st3_320  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[320]), .rdlo_in(a3_wr[448]),  .coef_in(coef[512]), .rdup_out(a4_wr[320]), .rdlo_out(a4_wr[448]));
			radix2 #(.width(width)) rd_st3_321  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[321]), .rdlo_in(a3_wr[449]),  .coef_in(coef[520]), .rdup_out(a4_wr[321]), .rdlo_out(a4_wr[449]));
			radix2 #(.width(width)) rd_st3_322  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[322]), .rdlo_in(a3_wr[450]),  .coef_in(coef[528]), .rdup_out(a4_wr[322]), .rdlo_out(a4_wr[450]));
			radix2 #(.width(width)) rd_st3_323  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[323]), .rdlo_in(a3_wr[451]),  .coef_in(coef[536]), .rdup_out(a4_wr[323]), .rdlo_out(a4_wr[451]));
			radix2 #(.width(width)) rd_st3_324  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[324]), .rdlo_in(a3_wr[452]),  .coef_in(coef[544]), .rdup_out(a4_wr[324]), .rdlo_out(a4_wr[452]));
			radix2 #(.width(width)) rd_st3_325  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[325]), .rdlo_in(a3_wr[453]),  .coef_in(coef[552]), .rdup_out(a4_wr[325]), .rdlo_out(a4_wr[453]));
			radix2 #(.width(width)) rd_st3_326  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[326]), .rdlo_in(a3_wr[454]),  .coef_in(coef[560]), .rdup_out(a4_wr[326]), .rdlo_out(a4_wr[454]));
			radix2 #(.width(width)) rd_st3_327  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[327]), .rdlo_in(a3_wr[455]),  .coef_in(coef[568]), .rdup_out(a4_wr[327]), .rdlo_out(a4_wr[455]));
			radix2 #(.width(width)) rd_st3_328  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[328]), .rdlo_in(a3_wr[456]),  .coef_in(coef[576]), .rdup_out(a4_wr[328]), .rdlo_out(a4_wr[456]));
			radix2 #(.width(width)) rd_st3_329  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[329]), .rdlo_in(a3_wr[457]),  .coef_in(coef[584]), .rdup_out(a4_wr[329]), .rdlo_out(a4_wr[457]));
			radix2 #(.width(width)) rd_st3_330  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[330]), .rdlo_in(a3_wr[458]),  .coef_in(coef[592]), .rdup_out(a4_wr[330]), .rdlo_out(a4_wr[458]));
			radix2 #(.width(width)) rd_st3_331  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[331]), .rdlo_in(a3_wr[459]),  .coef_in(coef[600]), .rdup_out(a4_wr[331]), .rdlo_out(a4_wr[459]));
			radix2 #(.width(width)) rd_st3_332  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[332]), .rdlo_in(a3_wr[460]),  .coef_in(coef[608]), .rdup_out(a4_wr[332]), .rdlo_out(a4_wr[460]));
			radix2 #(.width(width)) rd_st3_333  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[333]), .rdlo_in(a3_wr[461]),  .coef_in(coef[616]), .rdup_out(a4_wr[333]), .rdlo_out(a4_wr[461]));
			radix2 #(.width(width)) rd_st3_334  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[334]), .rdlo_in(a3_wr[462]),  .coef_in(coef[624]), .rdup_out(a4_wr[334]), .rdlo_out(a4_wr[462]));
			radix2 #(.width(width)) rd_st3_335  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[335]), .rdlo_in(a3_wr[463]),  .coef_in(coef[632]), .rdup_out(a4_wr[335]), .rdlo_out(a4_wr[463]));
			radix2 #(.width(width)) rd_st3_336  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[336]), .rdlo_in(a3_wr[464]),  .coef_in(coef[640]), .rdup_out(a4_wr[336]), .rdlo_out(a4_wr[464]));
			radix2 #(.width(width)) rd_st3_337  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[337]), .rdlo_in(a3_wr[465]),  .coef_in(coef[648]), .rdup_out(a4_wr[337]), .rdlo_out(a4_wr[465]));
			radix2 #(.width(width)) rd_st3_338  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[338]), .rdlo_in(a3_wr[466]),  .coef_in(coef[656]), .rdup_out(a4_wr[338]), .rdlo_out(a4_wr[466]));
			radix2 #(.width(width)) rd_st3_339  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[339]), .rdlo_in(a3_wr[467]),  .coef_in(coef[664]), .rdup_out(a4_wr[339]), .rdlo_out(a4_wr[467]));
			radix2 #(.width(width)) rd_st3_340  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[340]), .rdlo_in(a3_wr[468]),  .coef_in(coef[672]), .rdup_out(a4_wr[340]), .rdlo_out(a4_wr[468]));
			radix2 #(.width(width)) rd_st3_341  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[341]), .rdlo_in(a3_wr[469]),  .coef_in(coef[680]), .rdup_out(a4_wr[341]), .rdlo_out(a4_wr[469]));
			radix2 #(.width(width)) rd_st3_342  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[342]), .rdlo_in(a3_wr[470]),  .coef_in(coef[688]), .rdup_out(a4_wr[342]), .rdlo_out(a4_wr[470]));
			radix2 #(.width(width)) rd_st3_343  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[343]), .rdlo_in(a3_wr[471]),  .coef_in(coef[696]), .rdup_out(a4_wr[343]), .rdlo_out(a4_wr[471]));
			radix2 #(.width(width)) rd_st3_344  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[344]), .rdlo_in(a3_wr[472]),  .coef_in(coef[704]), .rdup_out(a4_wr[344]), .rdlo_out(a4_wr[472]));
			radix2 #(.width(width)) rd_st3_345  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[345]), .rdlo_in(a3_wr[473]),  .coef_in(coef[712]), .rdup_out(a4_wr[345]), .rdlo_out(a4_wr[473]));
			radix2 #(.width(width)) rd_st3_346  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[346]), .rdlo_in(a3_wr[474]),  .coef_in(coef[720]), .rdup_out(a4_wr[346]), .rdlo_out(a4_wr[474]));
			radix2 #(.width(width)) rd_st3_347  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[347]), .rdlo_in(a3_wr[475]),  .coef_in(coef[728]), .rdup_out(a4_wr[347]), .rdlo_out(a4_wr[475]));
			radix2 #(.width(width)) rd_st3_348  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[348]), .rdlo_in(a3_wr[476]),  .coef_in(coef[736]), .rdup_out(a4_wr[348]), .rdlo_out(a4_wr[476]));
			radix2 #(.width(width)) rd_st3_349  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[349]), .rdlo_in(a3_wr[477]),  .coef_in(coef[744]), .rdup_out(a4_wr[349]), .rdlo_out(a4_wr[477]));
			radix2 #(.width(width)) rd_st3_350  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[350]), .rdlo_in(a3_wr[478]),  .coef_in(coef[752]), .rdup_out(a4_wr[350]), .rdlo_out(a4_wr[478]));
			radix2 #(.width(width)) rd_st3_351  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[351]), .rdlo_in(a3_wr[479]),  .coef_in(coef[760]), .rdup_out(a4_wr[351]), .rdlo_out(a4_wr[479]));
			radix2 #(.width(width)) rd_st3_352  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[352]), .rdlo_in(a3_wr[480]),  .coef_in(coef[768]), .rdup_out(a4_wr[352]), .rdlo_out(a4_wr[480]));
			radix2 #(.width(width)) rd_st3_353  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[353]), .rdlo_in(a3_wr[481]),  .coef_in(coef[776]), .rdup_out(a4_wr[353]), .rdlo_out(a4_wr[481]));
			radix2 #(.width(width)) rd_st3_354  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[354]), .rdlo_in(a3_wr[482]),  .coef_in(coef[784]), .rdup_out(a4_wr[354]), .rdlo_out(a4_wr[482]));
			radix2 #(.width(width)) rd_st3_355  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[355]), .rdlo_in(a3_wr[483]),  .coef_in(coef[792]), .rdup_out(a4_wr[355]), .rdlo_out(a4_wr[483]));
			radix2 #(.width(width)) rd_st3_356  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[356]), .rdlo_in(a3_wr[484]),  .coef_in(coef[800]), .rdup_out(a4_wr[356]), .rdlo_out(a4_wr[484]));
			radix2 #(.width(width)) rd_st3_357  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[357]), .rdlo_in(a3_wr[485]),  .coef_in(coef[808]), .rdup_out(a4_wr[357]), .rdlo_out(a4_wr[485]));
			radix2 #(.width(width)) rd_st3_358  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[358]), .rdlo_in(a3_wr[486]),  .coef_in(coef[816]), .rdup_out(a4_wr[358]), .rdlo_out(a4_wr[486]));
			radix2 #(.width(width)) rd_st3_359  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[359]), .rdlo_in(a3_wr[487]),  .coef_in(coef[824]), .rdup_out(a4_wr[359]), .rdlo_out(a4_wr[487]));
			radix2 #(.width(width)) rd_st3_360  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[360]), .rdlo_in(a3_wr[488]),  .coef_in(coef[832]), .rdup_out(a4_wr[360]), .rdlo_out(a4_wr[488]));
			radix2 #(.width(width)) rd_st3_361  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[361]), .rdlo_in(a3_wr[489]),  .coef_in(coef[840]), .rdup_out(a4_wr[361]), .rdlo_out(a4_wr[489]));
			radix2 #(.width(width)) rd_st3_362  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[362]), .rdlo_in(a3_wr[490]),  .coef_in(coef[848]), .rdup_out(a4_wr[362]), .rdlo_out(a4_wr[490]));
			radix2 #(.width(width)) rd_st3_363  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[363]), .rdlo_in(a3_wr[491]),  .coef_in(coef[856]), .rdup_out(a4_wr[363]), .rdlo_out(a4_wr[491]));
			radix2 #(.width(width)) rd_st3_364  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[364]), .rdlo_in(a3_wr[492]),  .coef_in(coef[864]), .rdup_out(a4_wr[364]), .rdlo_out(a4_wr[492]));
			radix2 #(.width(width)) rd_st3_365  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[365]), .rdlo_in(a3_wr[493]),  .coef_in(coef[872]), .rdup_out(a4_wr[365]), .rdlo_out(a4_wr[493]));
			radix2 #(.width(width)) rd_st3_366  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[366]), .rdlo_in(a3_wr[494]),  .coef_in(coef[880]), .rdup_out(a4_wr[366]), .rdlo_out(a4_wr[494]));
			radix2 #(.width(width)) rd_st3_367  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[367]), .rdlo_in(a3_wr[495]),  .coef_in(coef[888]), .rdup_out(a4_wr[367]), .rdlo_out(a4_wr[495]));
			radix2 #(.width(width)) rd_st3_368  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[368]), .rdlo_in(a3_wr[496]),  .coef_in(coef[896]), .rdup_out(a4_wr[368]), .rdlo_out(a4_wr[496]));
			radix2 #(.width(width)) rd_st3_369  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[369]), .rdlo_in(a3_wr[497]),  .coef_in(coef[904]), .rdup_out(a4_wr[369]), .rdlo_out(a4_wr[497]));
			radix2 #(.width(width)) rd_st3_370  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[370]), .rdlo_in(a3_wr[498]),  .coef_in(coef[912]), .rdup_out(a4_wr[370]), .rdlo_out(a4_wr[498]));
			radix2 #(.width(width)) rd_st3_371  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[371]), .rdlo_in(a3_wr[499]),  .coef_in(coef[920]), .rdup_out(a4_wr[371]), .rdlo_out(a4_wr[499]));
			radix2 #(.width(width)) rd_st3_372  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[372]), .rdlo_in(a3_wr[500]),  .coef_in(coef[928]), .rdup_out(a4_wr[372]), .rdlo_out(a4_wr[500]));
			radix2 #(.width(width)) rd_st3_373  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[373]), .rdlo_in(a3_wr[501]),  .coef_in(coef[936]), .rdup_out(a4_wr[373]), .rdlo_out(a4_wr[501]));
			radix2 #(.width(width)) rd_st3_374  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[374]), .rdlo_in(a3_wr[502]),  .coef_in(coef[944]), .rdup_out(a4_wr[374]), .rdlo_out(a4_wr[502]));
			radix2 #(.width(width)) rd_st3_375  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[375]), .rdlo_in(a3_wr[503]),  .coef_in(coef[952]), .rdup_out(a4_wr[375]), .rdlo_out(a4_wr[503]));
			radix2 #(.width(width)) rd_st3_376  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[376]), .rdlo_in(a3_wr[504]),  .coef_in(coef[960]), .rdup_out(a4_wr[376]), .rdlo_out(a4_wr[504]));
			radix2 #(.width(width)) rd_st3_377  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[377]), .rdlo_in(a3_wr[505]),  .coef_in(coef[968]), .rdup_out(a4_wr[377]), .rdlo_out(a4_wr[505]));
			radix2 #(.width(width)) rd_st3_378  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[378]), .rdlo_in(a3_wr[506]),  .coef_in(coef[976]), .rdup_out(a4_wr[378]), .rdlo_out(a4_wr[506]));
			radix2 #(.width(width)) rd_st3_379  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[379]), .rdlo_in(a3_wr[507]),  .coef_in(coef[984]), .rdup_out(a4_wr[379]), .rdlo_out(a4_wr[507]));
			radix2 #(.width(width)) rd_st3_380  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[380]), .rdlo_in(a3_wr[508]),  .coef_in(coef[992]), .rdup_out(a4_wr[380]), .rdlo_out(a4_wr[508]));
			radix2 #(.width(width)) rd_st3_381  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[381]), .rdlo_in(a3_wr[509]),  .coef_in(coef[1000]), .rdup_out(a4_wr[381]), .rdlo_out(a4_wr[509]));
			radix2 #(.width(width)) rd_st3_382  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[382]), .rdlo_in(a3_wr[510]),  .coef_in(coef[1008]), .rdup_out(a4_wr[382]), .rdlo_out(a4_wr[510]));
			radix2 #(.width(width)) rd_st3_383  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[383]), .rdlo_in(a3_wr[511]),  .coef_in(coef[1016]), .rdup_out(a4_wr[383]), .rdlo_out(a4_wr[511]));
			radix2 #(.width(width)) rd_st3_512  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[512]), .rdlo_in(a3_wr[640]),  .coef_in(coef[0]), .rdup_out(a4_wr[512]), .rdlo_out(a4_wr[640]));
			radix2 #(.width(width)) rd_st3_513  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[513]), .rdlo_in(a3_wr[641]),  .coef_in(coef[8]), .rdup_out(a4_wr[513]), .rdlo_out(a4_wr[641]));
			radix2 #(.width(width)) rd_st3_514  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[514]), .rdlo_in(a3_wr[642]),  .coef_in(coef[16]), .rdup_out(a4_wr[514]), .rdlo_out(a4_wr[642]));
			radix2 #(.width(width)) rd_st3_515  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[515]), .rdlo_in(a3_wr[643]),  .coef_in(coef[24]), .rdup_out(a4_wr[515]), .rdlo_out(a4_wr[643]));
			radix2 #(.width(width)) rd_st3_516  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[516]), .rdlo_in(a3_wr[644]),  .coef_in(coef[32]), .rdup_out(a4_wr[516]), .rdlo_out(a4_wr[644]));
			radix2 #(.width(width)) rd_st3_517  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[517]), .rdlo_in(a3_wr[645]),  .coef_in(coef[40]), .rdup_out(a4_wr[517]), .rdlo_out(a4_wr[645]));
			radix2 #(.width(width)) rd_st3_518  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[518]), .rdlo_in(a3_wr[646]),  .coef_in(coef[48]), .rdup_out(a4_wr[518]), .rdlo_out(a4_wr[646]));
			radix2 #(.width(width)) rd_st3_519  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[519]), .rdlo_in(a3_wr[647]),  .coef_in(coef[56]), .rdup_out(a4_wr[519]), .rdlo_out(a4_wr[647]));
			radix2 #(.width(width)) rd_st3_520  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[520]), .rdlo_in(a3_wr[648]),  .coef_in(coef[64]), .rdup_out(a4_wr[520]), .rdlo_out(a4_wr[648]));
			radix2 #(.width(width)) rd_st3_521  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[521]), .rdlo_in(a3_wr[649]),  .coef_in(coef[72]), .rdup_out(a4_wr[521]), .rdlo_out(a4_wr[649]));
			radix2 #(.width(width)) rd_st3_522  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[522]), .rdlo_in(a3_wr[650]),  .coef_in(coef[80]), .rdup_out(a4_wr[522]), .rdlo_out(a4_wr[650]));
			radix2 #(.width(width)) rd_st3_523  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[523]), .rdlo_in(a3_wr[651]),  .coef_in(coef[88]), .rdup_out(a4_wr[523]), .rdlo_out(a4_wr[651]));
			radix2 #(.width(width)) rd_st3_524  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[524]), .rdlo_in(a3_wr[652]),  .coef_in(coef[96]), .rdup_out(a4_wr[524]), .rdlo_out(a4_wr[652]));
			radix2 #(.width(width)) rd_st3_525  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[525]), .rdlo_in(a3_wr[653]),  .coef_in(coef[104]), .rdup_out(a4_wr[525]), .rdlo_out(a4_wr[653]));
			radix2 #(.width(width)) rd_st3_526  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[526]), .rdlo_in(a3_wr[654]),  .coef_in(coef[112]), .rdup_out(a4_wr[526]), .rdlo_out(a4_wr[654]));
			radix2 #(.width(width)) rd_st3_527  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[527]), .rdlo_in(a3_wr[655]),  .coef_in(coef[120]), .rdup_out(a4_wr[527]), .rdlo_out(a4_wr[655]));
			radix2 #(.width(width)) rd_st3_528  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[528]), .rdlo_in(a3_wr[656]),  .coef_in(coef[128]), .rdup_out(a4_wr[528]), .rdlo_out(a4_wr[656]));
			radix2 #(.width(width)) rd_st3_529  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[529]), .rdlo_in(a3_wr[657]),  .coef_in(coef[136]), .rdup_out(a4_wr[529]), .rdlo_out(a4_wr[657]));
			radix2 #(.width(width)) rd_st3_530  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[530]), .rdlo_in(a3_wr[658]),  .coef_in(coef[144]), .rdup_out(a4_wr[530]), .rdlo_out(a4_wr[658]));
			radix2 #(.width(width)) rd_st3_531  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[531]), .rdlo_in(a3_wr[659]),  .coef_in(coef[152]), .rdup_out(a4_wr[531]), .rdlo_out(a4_wr[659]));
			radix2 #(.width(width)) rd_st3_532  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[532]), .rdlo_in(a3_wr[660]),  .coef_in(coef[160]), .rdup_out(a4_wr[532]), .rdlo_out(a4_wr[660]));
			radix2 #(.width(width)) rd_st3_533  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[533]), .rdlo_in(a3_wr[661]),  .coef_in(coef[168]), .rdup_out(a4_wr[533]), .rdlo_out(a4_wr[661]));
			radix2 #(.width(width)) rd_st3_534  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[534]), .rdlo_in(a3_wr[662]),  .coef_in(coef[176]), .rdup_out(a4_wr[534]), .rdlo_out(a4_wr[662]));
			radix2 #(.width(width)) rd_st3_535  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[535]), .rdlo_in(a3_wr[663]),  .coef_in(coef[184]), .rdup_out(a4_wr[535]), .rdlo_out(a4_wr[663]));
			radix2 #(.width(width)) rd_st3_536  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[536]), .rdlo_in(a3_wr[664]),  .coef_in(coef[192]), .rdup_out(a4_wr[536]), .rdlo_out(a4_wr[664]));
			radix2 #(.width(width)) rd_st3_537  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[537]), .rdlo_in(a3_wr[665]),  .coef_in(coef[200]), .rdup_out(a4_wr[537]), .rdlo_out(a4_wr[665]));
			radix2 #(.width(width)) rd_st3_538  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[538]), .rdlo_in(a3_wr[666]),  .coef_in(coef[208]), .rdup_out(a4_wr[538]), .rdlo_out(a4_wr[666]));
			radix2 #(.width(width)) rd_st3_539  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[539]), .rdlo_in(a3_wr[667]),  .coef_in(coef[216]), .rdup_out(a4_wr[539]), .rdlo_out(a4_wr[667]));
			radix2 #(.width(width)) rd_st3_540  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[540]), .rdlo_in(a3_wr[668]),  .coef_in(coef[224]), .rdup_out(a4_wr[540]), .rdlo_out(a4_wr[668]));
			radix2 #(.width(width)) rd_st3_541  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[541]), .rdlo_in(a3_wr[669]),  .coef_in(coef[232]), .rdup_out(a4_wr[541]), .rdlo_out(a4_wr[669]));
			radix2 #(.width(width)) rd_st3_542  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[542]), .rdlo_in(a3_wr[670]),  .coef_in(coef[240]), .rdup_out(a4_wr[542]), .rdlo_out(a4_wr[670]));
			radix2 #(.width(width)) rd_st3_543  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[543]), .rdlo_in(a3_wr[671]),  .coef_in(coef[248]), .rdup_out(a4_wr[543]), .rdlo_out(a4_wr[671]));
			radix2 #(.width(width)) rd_st3_544  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[544]), .rdlo_in(a3_wr[672]),  .coef_in(coef[256]), .rdup_out(a4_wr[544]), .rdlo_out(a4_wr[672]));
			radix2 #(.width(width)) rd_st3_545  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[545]), .rdlo_in(a3_wr[673]),  .coef_in(coef[264]), .rdup_out(a4_wr[545]), .rdlo_out(a4_wr[673]));
			radix2 #(.width(width)) rd_st3_546  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[546]), .rdlo_in(a3_wr[674]),  .coef_in(coef[272]), .rdup_out(a4_wr[546]), .rdlo_out(a4_wr[674]));
			radix2 #(.width(width)) rd_st3_547  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[547]), .rdlo_in(a3_wr[675]),  .coef_in(coef[280]), .rdup_out(a4_wr[547]), .rdlo_out(a4_wr[675]));
			radix2 #(.width(width)) rd_st3_548  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[548]), .rdlo_in(a3_wr[676]),  .coef_in(coef[288]), .rdup_out(a4_wr[548]), .rdlo_out(a4_wr[676]));
			radix2 #(.width(width)) rd_st3_549  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[549]), .rdlo_in(a3_wr[677]),  .coef_in(coef[296]), .rdup_out(a4_wr[549]), .rdlo_out(a4_wr[677]));
			radix2 #(.width(width)) rd_st3_550  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[550]), .rdlo_in(a3_wr[678]),  .coef_in(coef[304]), .rdup_out(a4_wr[550]), .rdlo_out(a4_wr[678]));
			radix2 #(.width(width)) rd_st3_551  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[551]), .rdlo_in(a3_wr[679]),  .coef_in(coef[312]), .rdup_out(a4_wr[551]), .rdlo_out(a4_wr[679]));
			radix2 #(.width(width)) rd_st3_552  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[552]), .rdlo_in(a3_wr[680]),  .coef_in(coef[320]), .rdup_out(a4_wr[552]), .rdlo_out(a4_wr[680]));
			radix2 #(.width(width)) rd_st3_553  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[553]), .rdlo_in(a3_wr[681]),  .coef_in(coef[328]), .rdup_out(a4_wr[553]), .rdlo_out(a4_wr[681]));
			radix2 #(.width(width)) rd_st3_554  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[554]), .rdlo_in(a3_wr[682]),  .coef_in(coef[336]), .rdup_out(a4_wr[554]), .rdlo_out(a4_wr[682]));
			radix2 #(.width(width)) rd_st3_555  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[555]), .rdlo_in(a3_wr[683]),  .coef_in(coef[344]), .rdup_out(a4_wr[555]), .rdlo_out(a4_wr[683]));
			radix2 #(.width(width)) rd_st3_556  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[556]), .rdlo_in(a3_wr[684]),  .coef_in(coef[352]), .rdup_out(a4_wr[556]), .rdlo_out(a4_wr[684]));
			radix2 #(.width(width)) rd_st3_557  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[557]), .rdlo_in(a3_wr[685]),  .coef_in(coef[360]), .rdup_out(a4_wr[557]), .rdlo_out(a4_wr[685]));
			radix2 #(.width(width)) rd_st3_558  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[558]), .rdlo_in(a3_wr[686]),  .coef_in(coef[368]), .rdup_out(a4_wr[558]), .rdlo_out(a4_wr[686]));
			radix2 #(.width(width)) rd_st3_559  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[559]), .rdlo_in(a3_wr[687]),  .coef_in(coef[376]), .rdup_out(a4_wr[559]), .rdlo_out(a4_wr[687]));
			radix2 #(.width(width)) rd_st3_560  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[560]), .rdlo_in(a3_wr[688]),  .coef_in(coef[384]), .rdup_out(a4_wr[560]), .rdlo_out(a4_wr[688]));
			radix2 #(.width(width)) rd_st3_561  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[561]), .rdlo_in(a3_wr[689]),  .coef_in(coef[392]), .rdup_out(a4_wr[561]), .rdlo_out(a4_wr[689]));
			radix2 #(.width(width)) rd_st3_562  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[562]), .rdlo_in(a3_wr[690]),  .coef_in(coef[400]), .rdup_out(a4_wr[562]), .rdlo_out(a4_wr[690]));
			radix2 #(.width(width)) rd_st3_563  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[563]), .rdlo_in(a3_wr[691]),  .coef_in(coef[408]), .rdup_out(a4_wr[563]), .rdlo_out(a4_wr[691]));
			radix2 #(.width(width)) rd_st3_564  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[564]), .rdlo_in(a3_wr[692]),  .coef_in(coef[416]), .rdup_out(a4_wr[564]), .rdlo_out(a4_wr[692]));
			radix2 #(.width(width)) rd_st3_565  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[565]), .rdlo_in(a3_wr[693]),  .coef_in(coef[424]), .rdup_out(a4_wr[565]), .rdlo_out(a4_wr[693]));
			radix2 #(.width(width)) rd_st3_566  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[566]), .rdlo_in(a3_wr[694]),  .coef_in(coef[432]), .rdup_out(a4_wr[566]), .rdlo_out(a4_wr[694]));
			radix2 #(.width(width)) rd_st3_567  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[567]), .rdlo_in(a3_wr[695]),  .coef_in(coef[440]), .rdup_out(a4_wr[567]), .rdlo_out(a4_wr[695]));
			radix2 #(.width(width)) rd_st3_568  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[568]), .rdlo_in(a3_wr[696]),  .coef_in(coef[448]), .rdup_out(a4_wr[568]), .rdlo_out(a4_wr[696]));
			radix2 #(.width(width)) rd_st3_569  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[569]), .rdlo_in(a3_wr[697]),  .coef_in(coef[456]), .rdup_out(a4_wr[569]), .rdlo_out(a4_wr[697]));
			radix2 #(.width(width)) rd_st3_570  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[570]), .rdlo_in(a3_wr[698]),  .coef_in(coef[464]), .rdup_out(a4_wr[570]), .rdlo_out(a4_wr[698]));
			radix2 #(.width(width)) rd_st3_571  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[571]), .rdlo_in(a3_wr[699]),  .coef_in(coef[472]), .rdup_out(a4_wr[571]), .rdlo_out(a4_wr[699]));
			radix2 #(.width(width)) rd_st3_572  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[572]), .rdlo_in(a3_wr[700]),  .coef_in(coef[480]), .rdup_out(a4_wr[572]), .rdlo_out(a4_wr[700]));
			radix2 #(.width(width)) rd_st3_573  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[573]), .rdlo_in(a3_wr[701]),  .coef_in(coef[488]), .rdup_out(a4_wr[573]), .rdlo_out(a4_wr[701]));
			radix2 #(.width(width)) rd_st3_574  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[574]), .rdlo_in(a3_wr[702]),  .coef_in(coef[496]), .rdup_out(a4_wr[574]), .rdlo_out(a4_wr[702]));
			radix2 #(.width(width)) rd_st3_575  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[575]), .rdlo_in(a3_wr[703]),  .coef_in(coef[504]), .rdup_out(a4_wr[575]), .rdlo_out(a4_wr[703]));
			radix2 #(.width(width)) rd_st3_576  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[576]), .rdlo_in(a3_wr[704]),  .coef_in(coef[512]), .rdup_out(a4_wr[576]), .rdlo_out(a4_wr[704]));
			radix2 #(.width(width)) rd_st3_577  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[577]), .rdlo_in(a3_wr[705]),  .coef_in(coef[520]), .rdup_out(a4_wr[577]), .rdlo_out(a4_wr[705]));
			radix2 #(.width(width)) rd_st3_578  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[578]), .rdlo_in(a3_wr[706]),  .coef_in(coef[528]), .rdup_out(a4_wr[578]), .rdlo_out(a4_wr[706]));
			radix2 #(.width(width)) rd_st3_579  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[579]), .rdlo_in(a3_wr[707]),  .coef_in(coef[536]), .rdup_out(a4_wr[579]), .rdlo_out(a4_wr[707]));
			radix2 #(.width(width)) rd_st3_580  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[580]), .rdlo_in(a3_wr[708]),  .coef_in(coef[544]), .rdup_out(a4_wr[580]), .rdlo_out(a4_wr[708]));
			radix2 #(.width(width)) rd_st3_581  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[581]), .rdlo_in(a3_wr[709]),  .coef_in(coef[552]), .rdup_out(a4_wr[581]), .rdlo_out(a4_wr[709]));
			radix2 #(.width(width)) rd_st3_582  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[582]), .rdlo_in(a3_wr[710]),  .coef_in(coef[560]), .rdup_out(a4_wr[582]), .rdlo_out(a4_wr[710]));
			radix2 #(.width(width)) rd_st3_583  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[583]), .rdlo_in(a3_wr[711]),  .coef_in(coef[568]), .rdup_out(a4_wr[583]), .rdlo_out(a4_wr[711]));
			radix2 #(.width(width)) rd_st3_584  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[584]), .rdlo_in(a3_wr[712]),  .coef_in(coef[576]), .rdup_out(a4_wr[584]), .rdlo_out(a4_wr[712]));
			radix2 #(.width(width)) rd_st3_585  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[585]), .rdlo_in(a3_wr[713]),  .coef_in(coef[584]), .rdup_out(a4_wr[585]), .rdlo_out(a4_wr[713]));
			radix2 #(.width(width)) rd_st3_586  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[586]), .rdlo_in(a3_wr[714]),  .coef_in(coef[592]), .rdup_out(a4_wr[586]), .rdlo_out(a4_wr[714]));
			radix2 #(.width(width)) rd_st3_587  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[587]), .rdlo_in(a3_wr[715]),  .coef_in(coef[600]), .rdup_out(a4_wr[587]), .rdlo_out(a4_wr[715]));
			radix2 #(.width(width)) rd_st3_588  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[588]), .rdlo_in(a3_wr[716]),  .coef_in(coef[608]), .rdup_out(a4_wr[588]), .rdlo_out(a4_wr[716]));
			radix2 #(.width(width)) rd_st3_589  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[589]), .rdlo_in(a3_wr[717]),  .coef_in(coef[616]), .rdup_out(a4_wr[589]), .rdlo_out(a4_wr[717]));
			radix2 #(.width(width)) rd_st3_590  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[590]), .rdlo_in(a3_wr[718]),  .coef_in(coef[624]), .rdup_out(a4_wr[590]), .rdlo_out(a4_wr[718]));
			radix2 #(.width(width)) rd_st3_591  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[591]), .rdlo_in(a3_wr[719]),  .coef_in(coef[632]), .rdup_out(a4_wr[591]), .rdlo_out(a4_wr[719]));
			radix2 #(.width(width)) rd_st3_592  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[592]), .rdlo_in(a3_wr[720]),  .coef_in(coef[640]), .rdup_out(a4_wr[592]), .rdlo_out(a4_wr[720]));
			radix2 #(.width(width)) rd_st3_593  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[593]), .rdlo_in(a3_wr[721]),  .coef_in(coef[648]), .rdup_out(a4_wr[593]), .rdlo_out(a4_wr[721]));
			radix2 #(.width(width)) rd_st3_594  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[594]), .rdlo_in(a3_wr[722]),  .coef_in(coef[656]), .rdup_out(a4_wr[594]), .rdlo_out(a4_wr[722]));
			radix2 #(.width(width)) rd_st3_595  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[595]), .rdlo_in(a3_wr[723]),  .coef_in(coef[664]), .rdup_out(a4_wr[595]), .rdlo_out(a4_wr[723]));
			radix2 #(.width(width)) rd_st3_596  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[596]), .rdlo_in(a3_wr[724]),  .coef_in(coef[672]), .rdup_out(a4_wr[596]), .rdlo_out(a4_wr[724]));
			radix2 #(.width(width)) rd_st3_597  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[597]), .rdlo_in(a3_wr[725]),  .coef_in(coef[680]), .rdup_out(a4_wr[597]), .rdlo_out(a4_wr[725]));
			radix2 #(.width(width)) rd_st3_598  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[598]), .rdlo_in(a3_wr[726]),  .coef_in(coef[688]), .rdup_out(a4_wr[598]), .rdlo_out(a4_wr[726]));
			radix2 #(.width(width)) rd_st3_599  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[599]), .rdlo_in(a3_wr[727]),  .coef_in(coef[696]), .rdup_out(a4_wr[599]), .rdlo_out(a4_wr[727]));
			radix2 #(.width(width)) rd_st3_600  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[600]), .rdlo_in(a3_wr[728]),  .coef_in(coef[704]), .rdup_out(a4_wr[600]), .rdlo_out(a4_wr[728]));
			radix2 #(.width(width)) rd_st3_601  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[601]), .rdlo_in(a3_wr[729]),  .coef_in(coef[712]), .rdup_out(a4_wr[601]), .rdlo_out(a4_wr[729]));
			radix2 #(.width(width)) rd_st3_602  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[602]), .rdlo_in(a3_wr[730]),  .coef_in(coef[720]), .rdup_out(a4_wr[602]), .rdlo_out(a4_wr[730]));
			radix2 #(.width(width)) rd_st3_603  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[603]), .rdlo_in(a3_wr[731]),  .coef_in(coef[728]), .rdup_out(a4_wr[603]), .rdlo_out(a4_wr[731]));
			radix2 #(.width(width)) rd_st3_604  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[604]), .rdlo_in(a3_wr[732]),  .coef_in(coef[736]), .rdup_out(a4_wr[604]), .rdlo_out(a4_wr[732]));
			radix2 #(.width(width)) rd_st3_605  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[605]), .rdlo_in(a3_wr[733]),  .coef_in(coef[744]), .rdup_out(a4_wr[605]), .rdlo_out(a4_wr[733]));
			radix2 #(.width(width)) rd_st3_606  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[606]), .rdlo_in(a3_wr[734]),  .coef_in(coef[752]), .rdup_out(a4_wr[606]), .rdlo_out(a4_wr[734]));
			radix2 #(.width(width)) rd_st3_607  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[607]), .rdlo_in(a3_wr[735]),  .coef_in(coef[760]), .rdup_out(a4_wr[607]), .rdlo_out(a4_wr[735]));
			radix2 #(.width(width)) rd_st3_608  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[608]), .rdlo_in(a3_wr[736]),  .coef_in(coef[768]), .rdup_out(a4_wr[608]), .rdlo_out(a4_wr[736]));
			radix2 #(.width(width)) rd_st3_609  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[609]), .rdlo_in(a3_wr[737]),  .coef_in(coef[776]), .rdup_out(a4_wr[609]), .rdlo_out(a4_wr[737]));
			radix2 #(.width(width)) rd_st3_610  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[610]), .rdlo_in(a3_wr[738]),  .coef_in(coef[784]), .rdup_out(a4_wr[610]), .rdlo_out(a4_wr[738]));
			radix2 #(.width(width)) rd_st3_611  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[611]), .rdlo_in(a3_wr[739]),  .coef_in(coef[792]), .rdup_out(a4_wr[611]), .rdlo_out(a4_wr[739]));
			radix2 #(.width(width)) rd_st3_612  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[612]), .rdlo_in(a3_wr[740]),  .coef_in(coef[800]), .rdup_out(a4_wr[612]), .rdlo_out(a4_wr[740]));
			radix2 #(.width(width)) rd_st3_613  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[613]), .rdlo_in(a3_wr[741]),  .coef_in(coef[808]), .rdup_out(a4_wr[613]), .rdlo_out(a4_wr[741]));
			radix2 #(.width(width)) rd_st3_614  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[614]), .rdlo_in(a3_wr[742]),  .coef_in(coef[816]), .rdup_out(a4_wr[614]), .rdlo_out(a4_wr[742]));
			radix2 #(.width(width)) rd_st3_615  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[615]), .rdlo_in(a3_wr[743]),  .coef_in(coef[824]), .rdup_out(a4_wr[615]), .rdlo_out(a4_wr[743]));
			radix2 #(.width(width)) rd_st3_616  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[616]), .rdlo_in(a3_wr[744]),  .coef_in(coef[832]), .rdup_out(a4_wr[616]), .rdlo_out(a4_wr[744]));
			radix2 #(.width(width)) rd_st3_617  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[617]), .rdlo_in(a3_wr[745]),  .coef_in(coef[840]), .rdup_out(a4_wr[617]), .rdlo_out(a4_wr[745]));
			radix2 #(.width(width)) rd_st3_618  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[618]), .rdlo_in(a3_wr[746]),  .coef_in(coef[848]), .rdup_out(a4_wr[618]), .rdlo_out(a4_wr[746]));
			radix2 #(.width(width)) rd_st3_619  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[619]), .rdlo_in(a3_wr[747]),  .coef_in(coef[856]), .rdup_out(a4_wr[619]), .rdlo_out(a4_wr[747]));
			radix2 #(.width(width)) rd_st3_620  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[620]), .rdlo_in(a3_wr[748]),  .coef_in(coef[864]), .rdup_out(a4_wr[620]), .rdlo_out(a4_wr[748]));
			radix2 #(.width(width)) rd_st3_621  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[621]), .rdlo_in(a3_wr[749]),  .coef_in(coef[872]), .rdup_out(a4_wr[621]), .rdlo_out(a4_wr[749]));
			radix2 #(.width(width)) rd_st3_622  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[622]), .rdlo_in(a3_wr[750]),  .coef_in(coef[880]), .rdup_out(a4_wr[622]), .rdlo_out(a4_wr[750]));
			radix2 #(.width(width)) rd_st3_623  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[623]), .rdlo_in(a3_wr[751]),  .coef_in(coef[888]), .rdup_out(a4_wr[623]), .rdlo_out(a4_wr[751]));
			radix2 #(.width(width)) rd_st3_624  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[624]), .rdlo_in(a3_wr[752]),  .coef_in(coef[896]), .rdup_out(a4_wr[624]), .rdlo_out(a4_wr[752]));
			radix2 #(.width(width)) rd_st3_625  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[625]), .rdlo_in(a3_wr[753]),  .coef_in(coef[904]), .rdup_out(a4_wr[625]), .rdlo_out(a4_wr[753]));
			radix2 #(.width(width)) rd_st3_626  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[626]), .rdlo_in(a3_wr[754]),  .coef_in(coef[912]), .rdup_out(a4_wr[626]), .rdlo_out(a4_wr[754]));
			radix2 #(.width(width)) rd_st3_627  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[627]), .rdlo_in(a3_wr[755]),  .coef_in(coef[920]), .rdup_out(a4_wr[627]), .rdlo_out(a4_wr[755]));
			radix2 #(.width(width)) rd_st3_628  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[628]), .rdlo_in(a3_wr[756]),  .coef_in(coef[928]), .rdup_out(a4_wr[628]), .rdlo_out(a4_wr[756]));
			radix2 #(.width(width)) rd_st3_629  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[629]), .rdlo_in(a3_wr[757]),  .coef_in(coef[936]), .rdup_out(a4_wr[629]), .rdlo_out(a4_wr[757]));
			radix2 #(.width(width)) rd_st3_630  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[630]), .rdlo_in(a3_wr[758]),  .coef_in(coef[944]), .rdup_out(a4_wr[630]), .rdlo_out(a4_wr[758]));
			radix2 #(.width(width)) rd_st3_631  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[631]), .rdlo_in(a3_wr[759]),  .coef_in(coef[952]), .rdup_out(a4_wr[631]), .rdlo_out(a4_wr[759]));
			radix2 #(.width(width)) rd_st3_632  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[632]), .rdlo_in(a3_wr[760]),  .coef_in(coef[960]), .rdup_out(a4_wr[632]), .rdlo_out(a4_wr[760]));
			radix2 #(.width(width)) rd_st3_633  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[633]), .rdlo_in(a3_wr[761]),  .coef_in(coef[968]), .rdup_out(a4_wr[633]), .rdlo_out(a4_wr[761]));
			radix2 #(.width(width)) rd_st3_634  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[634]), .rdlo_in(a3_wr[762]),  .coef_in(coef[976]), .rdup_out(a4_wr[634]), .rdlo_out(a4_wr[762]));
			radix2 #(.width(width)) rd_st3_635  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[635]), .rdlo_in(a3_wr[763]),  .coef_in(coef[984]), .rdup_out(a4_wr[635]), .rdlo_out(a4_wr[763]));
			radix2 #(.width(width)) rd_st3_636  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[636]), .rdlo_in(a3_wr[764]),  .coef_in(coef[992]), .rdup_out(a4_wr[636]), .rdlo_out(a4_wr[764]));
			radix2 #(.width(width)) rd_st3_637  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[637]), .rdlo_in(a3_wr[765]),  .coef_in(coef[1000]), .rdup_out(a4_wr[637]), .rdlo_out(a4_wr[765]));
			radix2 #(.width(width)) rd_st3_638  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[638]), .rdlo_in(a3_wr[766]),  .coef_in(coef[1008]), .rdup_out(a4_wr[638]), .rdlo_out(a4_wr[766]));
			radix2 #(.width(width)) rd_st3_639  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[639]), .rdlo_in(a3_wr[767]),  .coef_in(coef[1016]), .rdup_out(a4_wr[639]), .rdlo_out(a4_wr[767]));
			radix2 #(.width(width)) rd_st3_768  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[768]), .rdlo_in(a3_wr[896]),  .coef_in(coef[0]), .rdup_out(a4_wr[768]), .rdlo_out(a4_wr[896]));
			radix2 #(.width(width)) rd_st3_769  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[769]), .rdlo_in(a3_wr[897]),  .coef_in(coef[8]), .rdup_out(a4_wr[769]), .rdlo_out(a4_wr[897]));
			radix2 #(.width(width)) rd_st3_770  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[770]), .rdlo_in(a3_wr[898]),  .coef_in(coef[16]), .rdup_out(a4_wr[770]), .rdlo_out(a4_wr[898]));
			radix2 #(.width(width)) rd_st3_771  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[771]), .rdlo_in(a3_wr[899]),  .coef_in(coef[24]), .rdup_out(a4_wr[771]), .rdlo_out(a4_wr[899]));
			radix2 #(.width(width)) rd_st3_772  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[772]), .rdlo_in(a3_wr[900]),  .coef_in(coef[32]), .rdup_out(a4_wr[772]), .rdlo_out(a4_wr[900]));
			radix2 #(.width(width)) rd_st3_773  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[773]), .rdlo_in(a3_wr[901]),  .coef_in(coef[40]), .rdup_out(a4_wr[773]), .rdlo_out(a4_wr[901]));
			radix2 #(.width(width)) rd_st3_774  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[774]), .rdlo_in(a3_wr[902]),  .coef_in(coef[48]), .rdup_out(a4_wr[774]), .rdlo_out(a4_wr[902]));
			radix2 #(.width(width)) rd_st3_775  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[775]), .rdlo_in(a3_wr[903]),  .coef_in(coef[56]), .rdup_out(a4_wr[775]), .rdlo_out(a4_wr[903]));
			radix2 #(.width(width)) rd_st3_776  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[776]), .rdlo_in(a3_wr[904]),  .coef_in(coef[64]), .rdup_out(a4_wr[776]), .rdlo_out(a4_wr[904]));
			radix2 #(.width(width)) rd_st3_777  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[777]), .rdlo_in(a3_wr[905]),  .coef_in(coef[72]), .rdup_out(a4_wr[777]), .rdlo_out(a4_wr[905]));
			radix2 #(.width(width)) rd_st3_778  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[778]), .rdlo_in(a3_wr[906]),  .coef_in(coef[80]), .rdup_out(a4_wr[778]), .rdlo_out(a4_wr[906]));
			radix2 #(.width(width)) rd_st3_779  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[779]), .rdlo_in(a3_wr[907]),  .coef_in(coef[88]), .rdup_out(a4_wr[779]), .rdlo_out(a4_wr[907]));
			radix2 #(.width(width)) rd_st3_780  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[780]), .rdlo_in(a3_wr[908]),  .coef_in(coef[96]), .rdup_out(a4_wr[780]), .rdlo_out(a4_wr[908]));
			radix2 #(.width(width)) rd_st3_781  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[781]), .rdlo_in(a3_wr[909]),  .coef_in(coef[104]), .rdup_out(a4_wr[781]), .rdlo_out(a4_wr[909]));
			radix2 #(.width(width)) rd_st3_782  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[782]), .rdlo_in(a3_wr[910]),  .coef_in(coef[112]), .rdup_out(a4_wr[782]), .rdlo_out(a4_wr[910]));
			radix2 #(.width(width)) rd_st3_783  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[783]), .rdlo_in(a3_wr[911]),  .coef_in(coef[120]), .rdup_out(a4_wr[783]), .rdlo_out(a4_wr[911]));
			radix2 #(.width(width)) rd_st3_784  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[784]), .rdlo_in(a3_wr[912]),  .coef_in(coef[128]), .rdup_out(a4_wr[784]), .rdlo_out(a4_wr[912]));
			radix2 #(.width(width)) rd_st3_785  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[785]), .rdlo_in(a3_wr[913]),  .coef_in(coef[136]), .rdup_out(a4_wr[785]), .rdlo_out(a4_wr[913]));
			radix2 #(.width(width)) rd_st3_786  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[786]), .rdlo_in(a3_wr[914]),  .coef_in(coef[144]), .rdup_out(a4_wr[786]), .rdlo_out(a4_wr[914]));
			radix2 #(.width(width)) rd_st3_787  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[787]), .rdlo_in(a3_wr[915]),  .coef_in(coef[152]), .rdup_out(a4_wr[787]), .rdlo_out(a4_wr[915]));
			radix2 #(.width(width)) rd_st3_788  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[788]), .rdlo_in(a3_wr[916]),  .coef_in(coef[160]), .rdup_out(a4_wr[788]), .rdlo_out(a4_wr[916]));
			radix2 #(.width(width)) rd_st3_789  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[789]), .rdlo_in(a3_wr[917]),  .coef_in(coef[168]), .rdup_out(a4_wr[789]), .rdlo_out(a4_wr[917]));
			radix2 #(.width(width)) rd_st3_790  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[790]), .rdlo_in(a3_wr[918]),  .coef_in(coef[176]), .rdup_out(a4_wr[790]), .rdlo_out(a4_wr[918]));
			radix2 #(.width(width)) rd_st3_791  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[791]), .rdlo_in(a3_wr[919]),  .coef_in(coef[184]), .rdup_out(a4_wr[791]), .rdlo_out(a4_wr[919]));
			radix2 #(.width(width)) rd_st3_792  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[792]), .rdlo_in(a3_wr[920]),  .coef_in(coef[192]), .rdup_out(a4_wr[792]), .rdlo_out(a4_wr[920]));
			radix2 #(.width(width)) rd_st3_793  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[793]), .rdlo_in(a3_wr[921]),  .coef_in(coef[200]), .rdup_out(a4_wr[793]), .rdlo_out(a4_wr[921]));
			radix2 #(.width(width)) rd_st3_794  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[794]), .rdlo_in(a3_wr[922]),  .coef_in(coef[208]), .rdup_out(a4_wr[794]), .rdlo_out(a4_wr[922]));
			radix2 #(.width(width)) rd_st3_795  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[795]), .rdlo_in(a3_wr[923]),  .coef_in(coef[216]), .rdup_out(a4_wr[795]), .rdlo_out(a4_wr[923]));
			radix2 #(.width(width)) rd_st3_796  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[796]), .rdlo_in(a3_wr[924]),  .coef_in(coef[224]), .rdup_out(a4_wr[796]), .rdlo_out(a4_wr[924]));
			radix2 #(.width(width)) rd_st3_797  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[797]), .rdlo_in(a3_wr[925]),  .coef_in(coef[232]), .rdup_out(a4_wr[797]), .rdlo_out(a4_wr[925]));
			radix2 #(.width(width)) rd_st3_798  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[798]), .rdlo_in(a3_wr[926]),  .coef_in(coef[240]), .rdup_out(a4_wr[798]), .rdlo_out(a4_wr[926]));
			radix2 #(.width(width)) rd_st3_799  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[799]), .rdlo_in(a3_wr[927]),  .coef_in(coef[248]), .rdup_out(a4_wr[799]), .rdlo_out(a4_wr[927]));
			radix2 #(.width(width)) rd_st3_800  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[800]), .rdlo_in(a3_wr[928]),  .coef_in(coef[256]), .rdup_out(a4_wr[800]), .rdlo_out(a4_wr[928]));
			radix2 #(.width(width)) rd_st3_801  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[801]), .rdlo_in(a3_wr[929]),  .coef_in(coef[264]), .rdup_out(a4_wr[801]), .rdlo_out(a4_wr[929]));
			radix2 #(.width(width)) rd_st3_802  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[802]), .rdlo_in(a3_wr[930]),  .coef_in(coef[272]), .rdup_out(a4_wr[802]), .rdlo_out(a4_wr[930]));
			radix2 #(.width(width)) rd_st3_803  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[803]), .rdlo_in(a3_wr[931]),  .coef_in(coef[280]), .rdup_out(a4_wr[803]), .rdlo_out(a4_wr[931]));
			radix2 #(.width(width)) rd_st3_804  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[804]), .rdlo_in(a3_wr[932]),  .coef_in(coef[288]), .rdup_out(a4_wr[804]), .rdlo_out(a4_wr[932]));
			radix2 #(.width(width)) rd_st3_805  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[805]), .rdlo_in(a3_wr[933]),  .coef_in(coef[296]), .rdup_out(a4_wr[805]), .rdlo_out(a4_wr[933]));
			radix2 #(.width(width)) rd_st3_806  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[806]), .rdlo_in(a3_wr[934]),  .coef_in(coef[304]), .rdup_out(a4_wr[806]), .rdlo_out(a4_wr[934]));
			radix2 #(.width(width)) rd_st3_807  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[807]), .rdlo_in(a3_wr[935]),  .coef_in(coef[312]), .rdup_out(a4_wr[807]), .rdlo_out(a4_wr[935]));
			radix2 #(.width(width)) rd_st3_808  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[808]), .rdlo_in(a3_wr[936]),  .coef_in(coef[320]), .rdup_out(a4_wr[808]), .rdlo_out(a4_wr[936]));
			radix2 #(.width(width)) rd_st3_809  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[809]), .rdlo_in(a3_wr[937]),  .coef_in(coef[328]), .rdup_out(a4_wr[809]), .rdlo_out(a4_wr[937]));
			radix2 #(.width(width)) rd_st3_810  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[810]), .rdlo_in(a3_wr[938]),  .coef_in(coef[336]), .rdup_out(a4_wr[810]), .rdlo_out(a4_wr[938]));
			radix2 #(.width(width)) rd_st3_811  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[811]), .rdlo_in(a3_wr[939]),  .coef_in(coef[344]), .rdup_out(a4_wr[811]), .rdlo_out(a4_wr[939]));
			radix2 #(.width(width)) rd_st3_812  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[812]), .rdlo_in(a3_wr[940]),  .coef_in(coef[352]), .rdup_out(a4_wr[812]), .rdlo_out(a4_wr[940]));
			radix2 #(.width(width)) rd_st3_813  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[813]), .rdlo_in(a3_wr[941]),  .coef_in(coef[360]), .rdup_out(a4_wr[813]), .rdlo_out(a4_wr[941]));
			radix2 #(.width(width)) rd_st3_814  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[814]), .rdlo_in(a3_wr[942]),  .coef_in(coef[368]), .rdup_out(a4_wr[814]), .rdlo_out(a4_wr[942]));
			radix2 #(.width(width)) rd_st3_815  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[815]), .rdlo_in(a3_wr[943]),  .coef_in(coef[376]), .rdup_out(a4_wr[815]), .rdlo_out(a4_wr[943]));
			radix2 #(.width(width)) rd_st3_816  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[816]), .rdlo_in(a3_wr[944]),  .coef_in(coef[384]), .rdup_out(a4_wr[816]), .rdlo_out(a4_wr[944]));
			radix2 #(.width(width)) rd_st3_817  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[817]), .rdlo_in(a3_wr[945]),  .coef_in(coef[392]), .rdup_out(a4_wr[817]), .rdlo_out(a4_wr[945]));
			radix2 #(.width(width)) rd_st3_818  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[818]), .rdlo_in(a3_wr[946]),  .coef_in(coef[400]), .rdup_out(a4_wr[818]), .rdlo_out(a4_wr[946]));
			radix2 #(.width(width)) rd_st3_819  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[819]), .rdlo_in(a3_wr[947]),  .coef_in(coef[408]), .rdup_out(a4_wr[819]), .rdlo_out(a4_wr[947]));
			radix2 #(.width(width)) rd_st3_820  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[820]), .rdlo_in(a3_wr[948]),  .coef_in(coef[416]), .rdup_out(a4_wr[820]), .rdlo_out(a4_wr[948]));
			radix2 #(.width(width)) rd_st3_821  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[821]), .rdlo_in(a3_wr[949]),  .coef_in(coef[424]), .rdup_out(a4_wr[821]), .rdlo_out(a4_wr[949]));
			radix2 #(.width(width)) rd_st3_822  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[822]), .rdlo_in(a3_wr[950]),  .coef_in(coef[432]), .rdup_out(a4_wr[822]), .rdlo_out(a4_wr[950]));
			radix2 #(.width(width)) rd_st3_823  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[823]), .rdlo_in(a3_wr[951]),  .coef_in(coef[440]), .rdup_out(a4_wr[823]), .rdlo_out(a4_wr[951]));
			radix2 #(.width(width)) rd_st3_824  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[824]), .rdlo_in(a3_wr[952]),  .coef_in(coef[448]), .rdup_out(a4_wr[824]), .rdlo_out(a4_wr[952]));
			radix2 #(.width(width)) rd_st3_825  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[825]), .rdlo_in(a3_wr[953]),  .coef_in(coef[456]), .rdup_out(a4_wr[825]), .rdlo_out(a4_wr[953]));
			radix2 #(.width(width)) rd_st3_826  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[826]), .rdlo_in(a3_wr[954]),  .coef_in(coef[464]), .rdup_out(a4_wr[826]), .rdlo_out(a4_wr[954]));
			radix2 #(.width(width)) rd_st3_827  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[827]), .rdlo_in(a3_wr[955]),  .coef_in(coef[472]), .rdup_out(a4_wr[827]), .rdlo_out(a4_wr[955]));
			radix2 #(.width(width)) rd_st3_828  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[828]), .rdlo_in(a3_wr[956]),  .coef_in(coef[480]), .rdup_out(a4_wr[828]), .rdlo_out(a4_wr[956]));
			radix2 #(.width(width)) rd_st3_829  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[829]), .rdlo_in(a3_wr[957]),  .coef_in(coef[488]), .rdup_out(a4_wr[829]), .rdlo_out(a4_wr[957]));
			radix2 #(.width(width)) rd_st3_830  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[830]), .rdlo_in(a3_wr[958]),  .coef_in(coef[496]), .rdup_out(a4_wr[830]), .rdlo_out(a4_wr[958]));
			radix2 #(.width(width)) rd_st3_831  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[831]), .rdlo_in(a3_wr[959]),  .coef_in(coef[504]), .rdup_out(a4_wr[831]), .rdlo_out(a4_wr[959]));
			radix2 #(.width(width)) rd_st3_832  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[832]), .rdlo_in(a3_wr[960]),  .coef_in(coef[512]), .rdup_out(a4_wr[832]), .rdlo_out(a4_wr[960]));
			radix2 #(.width(width)) rd_st3_833  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[833]), .rdlo_in(a3_wr[961]),  .coef_in(coef[520]), .rdup_out(a4_wr[833]), .rdlo_out(a4_wr[961]));
			radix2 #(.width(width)) rd_st3_834  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[834]), .rdlo_in(a3_wr[962]),  .coef_in(coef[528]), .rdup_out(a4_wr[834]), .rdlo_out(a4_wr[962]));
			radix2 #(.width(width)) rd_st3_835  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[835]), .rdlo_in(a3_wr[963]),  .coef_in(coef[536]), .rdup_out(a4_wr[835]), .rdlo_out(a4_wr[963]));
			radix2 #(.width(width)) rd_st3_836  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[836]), .rdlo_in(a3_wr[964]),  .coef_in(coef[544]), .rdup_out(a4_wr[836]), .rdlo_out(a4_wr[964]));
			radix2 #(.width(width)) rd_st3_837  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[837]), .rdlo_in(a3_wr[965]),  .coef_in(coef[552]), .rdup_out(a4_wr[837]), .rdlo_out(a4_wr[965]));
			radix2 #(.width(width)) rd_st3_838  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[838]), .rdlo_in(a3_wr[966]),  .coef_in(coef[560]), .rdup_out(a4_wr[838]), .rdlo_out(a4_wr[966]));
			radix2 #(.width(width)) rd_st3_839  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[839]), .rdlo_in(a3_wr[967]),  .coef_in(coef[568]), .rdup_out(a4_wr[839]), .rdlo_out(a4_wr[967]));
			radix2 #(.width(width)) rd_st3_840  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[840]), .rdlo_in(a3_wr[968]),  .coef_in(coef[576]), .rdup_out(a4_wr[840]), .rdlo_out(a4_wr[968]));
			radix2 #(.width(width)) rd_st3_841  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[841]), .rdlo_in(a3_wr[969]),  .coef_in(coef[584]), .rdup_out(a4_wr[841]), .rdlo_out(a4_wr[969]));
			radix2 #(.width(width)) rd_st3_842  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[842]), .rdlo_in(a3_wr[970]),  .coef_in(coef[592]), .rdup_out(a4_wr[842]), .rdlo_out(a4_wr[970]));
			radix2 #(.width(width)) rd_st3_843  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[843]), .rdlo_in(a3_wr[971]),  .coef_in(coef[600]), .rdup_out(a4_wr[843]), .rdlo_out(a4_wr[971]));
			radix2 #(.width(width)) rd_st3_844  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[844]), .rdlo_in(a3_wr[972]),  .coef_in(coef[608]), .rdup_out(a4_wr[844]), .rdlo_out(a4_wr[972]));
			radix2 #(.width(width)) rd_st3_845  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[845]), .rdlo_in(a3_wr[973]),  .coef_in(coef[616]), .rdup_out(a4_wr[845]), .rdlo_out(a4_wr[973]));
			radix2 #(.width(width)) rd_st3_846  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[846]), .rdlo_in(a3_wr[974]),  .coef_in(coef[624]), .rdup_out(a4_wr[846]), .rdlo_out(a4_wr[974]));
			radix2 #(.width(width)) rd_st3_847  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[847]), .rdlo_in(a3_wr[975]),  .coef_in(coef[632]), .rdup_out(a4_wr[847]), .rdlo_out(a4_wr[975]));
			radix2 #(.width(width)) rd_st3_848  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[848]), .rdlo_in(a3_wr[976]),  .coef_in(coef[640]), .rdup_out(a4_wr[848]), .rdlo_out(a4_wr[976]));
			radix2 #(.width(width)) rd_st3_849  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[849]), .rdlo_in(a3_wr[977]),  .coef_in(coef[648]), .rdup_out(a4_wr[849]), .rdlo_out(a4_wr[977]));
			radix2 #(.width(width)) rd_st3_850  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[850]), .rdlo_in(a3_wr[978]),  .coef_in(coef[656]), .rdup_out(a4_wr[850]), .rdlo_out(a4_wr[978]));
			radix2 #(.width(width)) rd_st3_851  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[851]), .rdlo_in(a3_wr[979]),  .coef_in(coef[664]), .rdup_out(a4_wr[851]), .rdlo_out(a4_wr[979]));
			radix2 #(.width(width)) rd_st3_852  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[852]), .rdlo_in(a3_wr[980]),  .coef_in(coef[672]), .rdup_out(a4_wr[852]), .rdlo_out(a4_wr[980]));
			radix2 #(.width(width)) rd_st3_853  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[853]), .rdlo_in(a3_wr[981]),  .coef_in(coef[680]), .rdup_out(a4_wr[853]), .rdlo_out(a4_wr[981]));
			radix2 #(.width(width)) rd_st3_854  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[854]), .rdlo_in(a3_wr[982]),  .coef_in(coef[688]), .rdup_out(a4_wr[854]), .rdlo_out(a4_wr[982]));
			radix2 #(.width(width)) rd_st3_855  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[855]), .rdlo_in(a3_wr[983]),  .coef_in(coef[696]), .rdup_out(a4_wr[855]), .rdlo_out(a4_wr[983]));
			radix2 #(.width(width)) rd_st3_856  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[856]), .rdlo_in(a3_wr[984]),  .coef_in(coef[704]), .rdup_out(a4_wr[856]), .rdlo_out(a4_wr[984]));
			radix2 #(.width(width)) rd_st3_857  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[857]), .rdlo_in(a3_wr[985]),  .coef_in(coef[712]), .rdup_out(a4_wr[857]), .rdlo_out(a4_wr[985]));
			radix2 #(.width(width)) rd_st3_858  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[858]), .rdlo_in(a3_wr[986]),  .coef_in(coef[720]), .rdup_out(a4_wr[858]), .rdlo_out(a4_wr[986]));
			radix2 #(.width(width)) rd_st3_859  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[859]), .rdlo_in(a3_wr[987]),  .coef_in(coef[728]), .rdup_out(a4_wr[859]), .rdlo_out(a4_wr[987]));
			radix2 #(.width(width)) rd_st3_860  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[860]), .rdlo_in(a3_wr[988]),  .coef_in(coef[736]), .rdup_out(a4_wr[860]), .rdlo_out(a4_wr[988]));
			radix2 #(.width(width)) rd_st3_861  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[861]), .rdlo_in(a3_wr[989]),  .coef_in(coef[744]), .rdup_out(a4_wr[861]), .rdlo_out(a4_wr[989]));
			radix2 #(.width(width)) rd_st3_862  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[862]), .rdlo_in(a3_wr[990]),  .coef_in(coef[752]), .rdup_out(a4_wr[862]), .rdlo_out(a4_wr[990]));
			radix2 #(.width(width)) rd_st3_863  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[863]), .rdlo_in(a3_wr[991]),  .coef_in(coef[760]), .rdup_out(a4_wr[863]), .rdlo_out(a4_wr[991]));
			radix2 #(.width(width)) rd_st3_864  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[864]), .rdlo_in(a3_wr[992]),  .coef_in(coef[768]), .rdup_out(a4_wr[864]), .rdlo_out(a4_wr[992]));
			radix2 #(.width(width)) rd_st3_865  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[865]), .rdlo_in(a3_wr[993]),  .coef_in(coef[776]), .rdup_out(a4_wr[865]), .rdlo_out(a4_wr[993]));
			radix2 #(.width(width)) rd_st3_866  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[866]), .rdlo_in(a3_wr[994]),  .coef_in(coef[784]), .rdup_out(a4_wr[866]), .rdlo_out(a4_wr[994]));
			radix2 #(.width(width)) rd_st3_867  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[867]), .rdlo_in(a3_wr[995]),  .coef_in(coef[792]), .rdup_out(a4_wr[867]), .rdlo_out(a4_wr[995]));
			radix2 #(.width(width)) rd_st3_868  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[868]), .rdlo_in(a3_wr[996]),  .coef_in(coef[800]), .rdup_out(a4_wr[868]), .rdlo_out(a4_wr[996]));
			radix2 #(.width(width)) rd_st3_869  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[869]), .rdlo_in(a3_wr[997]),  .coef_in(coef[808]), .rdup_out(a4_wr[869]), .rdlo_out(a4_wr[997]));
			radix2 #(.width(width)) rd_st3_870  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[870]), .rdlo_in(a3_wr[998]),  .coef_in(coef[816]), .rdup_out(a4_wr[870]), .rdlo_out(a4_wr[998]));
			radix2 #(.width(width)) rd_st3_871  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[871]), .rdlo_in(a3_wr[999]),  .coef_in(coef[824]), .rdup_out(a4_wr[871]), .rdlo_out(a4_wr[999]));
			radix2 #(.width(width)) rd_st3_872  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[872]), .rdlo_in(a3_wr[1000]),  .coef_in(coef[832]), .rdup_out(a4_wr[872]), .rdlo_out(a4_wr[1000]));
			radix2 #(.width(width)) rd_st3_873  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[873]), .rdlo_in(a3_wr[1001]),  .coef_in(coef[840]), .rdup_out(a4_wr[873]), .rdlo_out(a4_wr[1001]));
			radix2 #(.width(width)) rd_st3_874  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[874]), .rdlo_in(a3_wr[1002]),  .coef_in(coef[848]), .rdup_out(a4_wr[874]), .rdlo_out(a4_wr[1002]));
			radix2 #(.width(width)) rd_st3_875  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[875]), .rdlo_in(a3_wr[1003]),  .coef_in(coef[856]), .rdup_out(a4_wr[875]), .rdlo_out(a4_wr[1003]));
			radix2 #(.width(width)) rd_st3_876  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[876]), .rdlo_in(a3_wr[1004]),  .coef_in(coef[864]), .rdup_out(a4_wr[876]), .rdlo_out(a4_wr[1004]));
			radix2 #(.width(width)) rd_st3_877  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[877]), .rdlo_in(a3_wr[1005]),  .coef_in(coef[872]), .rdup_out(a4_wr[877]), .rdlo_out(a4_wr[1005]));
			radix2 #(.width(width)) rd_st3_878  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[878]), .rdlo_in(a3_wr[1006]),  .coef_in(coef[880]), .rdup_out(a4_wr[878]), .rdlo_out(a4_wr[1006]));
			radix2 #(.width(width)) rd_st3_879  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[879]), .rdlo_in(a3_wr[1007]),  .coef_in(coef[888]), .rdup_out(a4_wr[879]), .rdlo_out(a4_wr[1007]));
			radix2 #(.width(width)) rd_st3_880  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[880]), .rdlo_in(a3_wr[1008]),  .coef_in(coef[896]), .rdup_out(a4_wr[880]), .rdlo_out(a4_wr[1008]));
			radix2 #(.width(width)) rd_st3_881  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[881]), .rdlo_in(a3_wr[1009]),  .coef_in(coef[904]), .rdup_out(a4_wr[881]), .rdlo_out(a4_wr[1009]));
			radix2 #(.width(width)) rd_st3_882  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[882]), .rdlo_in(a3_wr[1010]),  .coef_in(coef[912]), .rdup_out(a4_wr[882]), .rdlo_out(a4_wr[1010]));
			radix2 #(.width(width)) rd_st3_883  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[883]), .rdlo_in(a3_wr[1011]),  .coef_in(coef[920]), .rdup_out(a4_wr[883]), .rdlo_out(a4_wr[1011]));
			radix2 #(.width(width)) rd_st3_884  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[884]), .rdlo_in(a3_wr[1012]),  .coef_in(coef[928]), .rdup_out(a4_wr[884]), .rdlo_out(a4_wr[1012]));
			radix2 #(.width(width)) rd_st3_885  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[885]), .rdlo_in(a3_wr[1013]),  .coef_in(coef[936]), .rdup_out(a4_wr[885]), .rdlo_out(a4_wr[1013]));
			radix2 #(.width(width)) rd_st3_886  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[886]), .rdlo_in(a3_wr[1014]),  .coef_in(coef[944]), .rdup_out(a4_wr[886]), .rdlo_out(a4_wr[1014]));
			radix2 #(.width(width)) rd_st3_887  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[887]), .rdlo_in(a3_wr[1015]),  .coef_in(coef[952]), .rdup_out(a4_wr[887]), .rdlo_out(a4_wr[1015]));
			radix2 #(.width(width)) rd_st3_888  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[888]), .rdlo_in(a3_wr[1016]),  .coef_in(coef[960]), .rdup_out(a4_wr[888]), .rdlo_out(a4_wr[1016]));
			radix2 #(.width(width)) rd_st3_889  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[889]), .rdlo_in(a3_wr[1017]),  .coef_in(coef[968]), .rdup_out(a4_wr[889]), .rdlo_out(a4_wr[1017]));
			radix2 #(.width(width)) rd_st3_890  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[890]), .rdlo_in(a3_wr[1018]),  .coef_in(coef[976]), .rdup_out(a4_wr[890]), .rdlo_out(a4_wr[1018]));
			radix2 #(.width(width)) rd_st3_891  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[891]), .rdlo_in(a3_wr[1019]),  .coef_in(coef[984]), .rdup_out(a4_wr[891]), .rdlo_out(a4_wr[1019]));
			radix2 #(.width(width)) rd_st3_892  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[892]), .rdlo_in(a3_wr[1020]),  .coef_in(coef[992]), .rdup_out(a4_wr[892]), .rdlo_out(a4_wr[1020]));
			radix2 #(.width(width)) rd_st3_893  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[893]), .rdlo_in(a3_wr[1021]),  .coef_in(coef[1000]), .rdup_out(a4_wr[893]), .rdlo_out(a4_wr[1021]));
			radix2 #(.width(width)) rd_st3_894  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[894]), .rdlo_in(a3_wr[1022]),  .coef_in(coef[1008]), .rdup_out(a4_wr[894]), .rdlo_out(a4_wr[1022]));
			radix2 #(.width(width)) rd_st3_895  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[895]), .rdlo_in(a3_wr[1023]),  .coef_in(coef[1016]), .rdup_out(a4_wr[895]), .rdlo_out(a4_wr[1023]));
			radix2 #(.width(width)) rd_st3_1024  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1024]), .rdlo_in(a3_wr[1152]),  .coef_in(coef[0]), .rdup_out(a4_wr[1024]), .rdlo_out(a4_wr[1152]));
			radix2 #(.width(width)) rd_st3_1025  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1025]), .rdlo_in(a3_wr[1153]),  .coef_in(coef[8]), .rdup_out(a4_wr[1025]), .rdlo_out(a4_wr[1153]));
			radix2 #(.width(width)) rd_st3_1026  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1026]), .rdlo_in(a3_wr[1154]),  .coef_in(coef[16]), .rdup_out(a4_wr[1026]), .rdlo_out(a4_wr[1154]));
			radix2 #(.width(width)) rd_st3_1027  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1027]), .rdlo_in(a3_wr[1155]),  .coef_in(coef[24]), .rdup_out(a4_wr[1027]), .rdlo_out(a4_wr[1155]));
			radix2 #(.width(width)) rd_st3_1028  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1028]), .rdlo_in(a3_wr[1156]),  .coef_in(coef[32]), .rdup_out(a4_wr[1028]), .rdlo_out(a4_wr[1156]));
			radix2 #(.width(width)) rd_st3_1029  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1029]), .rdlo_in(a3_wr[1157]),  .coef_in(coef[40]), .rdup_out(a4_wr[1029]), .rdlo_out(a4_wr[1157]));
			radix2 #(.width(width)) rd_st3_1030  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1030]), .rdlo_in(a3_wr[1158]),  .coef_in(coef[48]), .rdup_out(a4_wr[1030]), .rdlo_out(a4_wr[1158]));
			radix2 #(.width(width)) rd_st3_1031  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1031]), .rdlo_in(a3_wr[1159]),  .coef_in(coef[56]), .rdup_out(a4_wr[1031]), .rdlo_out(a4_wr[1159]));
			radix2 #(.width(width)) rd_st3_1032  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1032]), .rdlo_in(a3_wr[1160]),  .coef_in(coef[64]), .rdup_out(a4_wr[1032]), .rdlo_out(a4_wr[1160]));
			radix2 #(.width(width)) rd_st3_1033  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1033]), .rdlo_in(a3_wr[1161]),  .coef_in(coef[72]), .rdup_out(a4_wr[1033]), .rdlo_out(a4_wr[1161]));
			radix2 #(.width(width)) rd_st3_1034  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1034]), .rdlo_in(a3_wr[1162]),  .coef_in(coef[80]), .rdup_out(a4_wr[1034]), .rdlo_out(a4_wr[1162]));
			radix2 #(.width(width)) rd_st3_1035  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1035]), .rdlo_in(a3_wr[1163]),  .coef_in(coef[88]), .rdup_out(a4_wr[1035]), .rdlo_out(a4_wr[1163]));
			radix2 #(.width(width)) rd_st3_1036  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1036]), .rdlo_in(a3_wr[1164]),  .coef_in(coef[96]), .rdup_out(a4_wr[1036]), .rdlo_out(a4_wr[1164]));
			radix2 #(.width(width)) rd_st3_1037  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1037]), .rdlo_in(a3_wr[1165]),  .coef_in(coef[104]), .rdup_out(a4_wr[1037]), .rdlo_out(a4_wr[1165]));
			radix2 #(.width(width)) rd_st3_1038  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1038]), .rdlo_in(a3_wr[1166]),  .coef_in(coef[112]), .rdup_out(a4_wr[1038]), .rdlo_out(a4_wr[1166]));
			radix2 #(.width(width)) rd_st3_1039  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1039]), .rdlo_in(a3_wr[1167]),  .coef_in(coef[120]), .rdup_out(a4_wr[1039]), .rdlo_out(a4_wr[1167]));
			radix2 #(.width(width)) rd_st3_1040  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1040]), .rdlo_in(a3_wr[1168]),  .coef_in(coef[128]), .rdup_out(a4_wr[1040]), .rdlo_out(a4_wr[1168]));
			radix2 #(.width(width)) rd_st3_1041  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1041]), .rdlo_in(a3_wr[1169]),  .coef_in(coef[136]), .rdup_out(a4_wr[1041]), .rdlo_out(a4_wr[1169]));
			radix2 #(.width(width)) rd_st3_1042  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1042]), .rdlo_in(a3_wr[1170]),  .coef_in(coef[144]), .rdup_out(a4_wr[1042]), .rdlo_out(a4_wr[1170]));
			radix2 #(.width(width)) rd_st3_1043  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1043]), .rdlo_in(a3_wr[1171]),  .coef_in(coef[152]), .rdup_out(a4_wr[1043]), .rdlo_out(a4_wr[1171]));
			radix2 #(.width(width)) rd_st3_1044  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1044]), .rdlo_in(a3_wr[1172]),  .coef_in(coef[160]), .rdup_out(a4_wr[1044]), .rdlo_out(a4_wr[1172]));
			radix2 #(.width(width)) rd_st3_1045  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1045]), .rdlo_in(a3_wr[1173]),  .coef_in(coef[168]), .rdup_out(a4_wr[1045]), .rdlo_out(a4_wr[1173]));
			radix2 #(.width(width)) rd_st3_1046  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1046]), .rdlo_in(a3_wr[1174]),  .coef_in(coef[176]), .rdup_out(a4_wr[1046]), .rdlo_out(a4_wr[1174]));
			radix2 #(.width(width)) rd_st3_1047  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1047]), .rdlo_in(a3_wr[1175]),  .coef_in(coef[184]), .rdup_out(a4_wr[1047]), .rdlo_out(a4_wr[1175]));
			radix2 #(.width(width)) rd_st3_1048  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1048]), .rdlo_in(a3_wr[1176]),  .coef_in(coef[192]), .rdup_out(a4_wr[1048]), .rdlo_out(a4_wr[1176]));
			radix2 #(.width(width)) rd_st3_1049  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1049]), .rdlo_in(a3_wr[1177]),  .coef_in(coef[200]), .rdup_out(a4_wr[1049]), .rdlo_out(a4_wr[1177]));
			radix2 #(.width(width)) rd_st3_1050  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1050]), .rdlo_in(a3_wr[1178]),  .coef_in(coef[208]), .rdup_out(a4_wr[1050]), .rdlo_out(a4_wr[1178]));
			radix2 #(.width(width)) rd_st3_1051  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1051]), .rdlo_in(a3_wr[1179]),  .coef_in(coef[216]), .rdup_out(a4_wr[1051]), .rdlo_out(a4_wr[1179]));
			radix2 #(.width(width)) rd_st3_1052  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1052]), .rdlo_in(a3_wr[1180]),  .coef_in(coef[224]), .rdup_out(a4_wr[1052]), .rdlo_out(a4_wr[1180]));
			radix2 #(.width(width)) rd_st3_1053  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1053]), .rdlo_in(a3_wr[1181]),  .coef_in(coef[232]), .rdup_out(a4_wr[1053]), .rdlo_out(a4_wr[1181]));
			radix2 #(.width(width)) rd_st3_1054  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1054]), .rdlo_in(a3_wr[1182]),  .coef_in(coef[240]), .rdup_out(a4_wr[1054]), .rdlo_out(a4_wr[1182]));
			radix2 #(.width(width)) rd_st3_1055  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1055]), .rdlo_in(a3_wr[1183]),  .coef_in(coef[248]), .rdup_out(a4_wr[1055]), .rdlo_out(a4_wr[1183]));
			radix2 #(.width(width)) rd_st3_1056  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1056]), .rdlo_in(a3_wr[1184]),  .coef_in(coef[256]), .rdup_out(a4_wr[1056]), .rdlo_out(a4_wr[1184]));
			radix2 #(.width(width)) rd_st3_1057  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1057]), .rdlo_in(a3_wr[1185]),  .coef_in(coef[264]), .rdup_out(a4_wr[1057]), .rdlo_out(a4_wr[1185]));
			radix2 #(.width(width)) rd_st3_1058  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1058]), .rdlo_in(a3_wr[1186]),  .coef_in(coef[272]), .rdup_out(a4_wr[1058]), .rdlo_out(a4_wr[1186]));
			radix2 #(.width(width)) rd_st3_1059  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1059]), .rdlo_in(a3_wr[1187]),  .coef_in(coef[280]), .rdup_out(a4_wr[1059]), .rdlo_out(a4_wr[1187]));
			radix2 #(.width(width)) rd_st3_1060  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1060]), .rdlo_in(a3_wr[1188]),  .coef_in(coef[288]), .rdup_out(a4_wr[1060]), .rdlo_out(a4_wr[1188]));
			radix2 #(.width(width)) rd_st3_1061  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1061]), .rdlo_in(a3_wr[1189]),  .coef_in(coef[296]), .rdup_out(a4_wr[1061]), .rdlo_out(a4_wr[1189]));
			radix2 #(.width(width)) rd_st3_1062  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1062]), .rdlo_in(a3_wr[1190]),  .coef_in(coef[304]), .rdup_out(a4_wr[1062]), .rdlo_out(a4_wr[1190]));
			radix2 #(.width(width)) rd_st3_1063  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1063]), .rdlo_in(a3_wr[1191]),  .coef_in(coef[312]), .rdup_out(a4_wr[1063]), .rdlo_out(a4_wr[1191]));
			radix2 #(.width(width)) rd_st3_1064  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1064]), .rdlo_in(a3_wr[1192]),  .coef_in(coef[320]), .rdup_out(a4_wr[1064]), .rdlo_out(a4_wr[1192]));
			radix2 #(.width(width)) rd_st3_1065  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1065]), .rdlo_in(a3_wr[1193]),  .coef_in(coef[328]), .rdup_out(a4_wr[1065]), .rdlo_out(a4_wr[1193]));
			radix2 #(.width(width)) rd_st3_1066  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1066]), .rdlo_in(a3_wr[1194]),  .coef_in(coef[336]), .rdup_out(a4_wr[1066]), .rdlo_out(a4_wr[1194]));
			radix2 #(.width(width)) rd_st3_1067  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1067]), .rdlo_in(a3_wr[1195]),  .coef_in(coef[344]), .rdup_out(a4_wr[1067]), .rdlo_out(a4_wr[1195]));
			radix2 #(.width(width)) rd_st3_1068  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1068]), .rdlo_in(a3_wr[1196]),  .coef_in(coef[352]), .rdup_out(a4_wr[1068]), .rdlo_out(a4_wr[1196]));
			radix2 #(.width(width)) rd_st3_1069  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1069]), .rdlo_in(a3_wr[1197]),  .coef_in(coef[360]), .rdup_out(a4_wr[1069]), .rdlo_out(a4_wr[1197]));
			radix2 #(.width(width)) rd_st3_1070  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1070]), .rdlo_in(a3_wr[1198]),  .coef_in(coef[368]), .rdup_out(a4_wr[1070]), .rdlo_out(a4_wr[1198]));
			radix2 #(.width(width)) rd_st3_1071  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1071]), .rdlo_in(a3_wr[1199]),  .coef_in(coef[376]), .rdup_out(a4_wr[1071]), .rdlo_out(a4_wr[1199]));
			radix2 #(.width(width)) rd_st3_1072  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1072]), .rdlo_in(a3_wr[1200]),  .coef_in(coef[384]), .rdup_out(a4_wr[1072]), .rdlo_out(a4_wr[1200]));
			radix2 #(.width(width)) rd_st3_1073  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1073]), .rdlo_in(a3_wr[1201]),  .coef_in(coef[392]), .rdup_out(a4_wr[1073]), .rdlo_out(a4_wr[1201]));
			radix2 #(.width(width)) rd_st3_1074  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1074]), .rdlo_in(a3_wr[1202]),  .coef_in(coef[400]), .rdup_out(a4_wr[1074]), .rdlo_out(a4_wr[1202]));
			radix2 #(.width(width)) rd_st3_1075  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1075]), .rdlo_in(a3_wr[1203]),  .coef_in(coef[408]), .rdup_out(a4_wr[1075]), .rdlo_out(a4_wr[1203]));
			radix2 #(.width(width)) rd_st3_1076  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1076]), .rdlo_in(a3_wr[1204]),  .coef_in(coef[416]), .rdup_out(a4_wr[1076]), .rdlo_out(a4_wr[1204]));
			radix2 #(.width(width)) rd_st3_1077  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1077]), .rdlo_in(a3_wr[1205]),  .coef_in(coef[424]), .rdup_out(a4_wr[1077]), .rdlo_out(a4_wr[1205]));
			radix2 #(.width(width)) rd_st3_1078  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1078]), .rdlo_in(a3_wr[1206]),  .coef_in(coef[432]), .rdup_out(a4_wr[1078]), .rdlo_out(a4_wr[1206]));
			radix2 #(.width(width)) rd_st3_1079  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1079]), .rdlo_in(a3_wr[1207]),  .coef_in(coef[440]), .rdup_out(a4_wr[1079]), .rdlo_out(a4_wr[1207]));
			radix2 #(.width(width)) rd_st3_1080  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1080]), .rdlo_in(a3_wr[1208]),  .coef_in(coef[448]), .rdup_out(a4_wr[1080]), .rdlo_out(a4_wr[1208]));
			radix2 #(.width(width)) rd_st3_1081  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1081]), .rdlo_in(a3_wr[1209]),  .coef_in(coef[456]), .rdup_out(a4_wr[1081]), .rdlo_out(a4_wr[1209]));
			radix2 #(.width(width)) rd_st3_1082  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1082]), .rdlo_in(a3_wr[1210]),  .coef_in(coef[464]), .rdup_out(a4_wr[1082]), .rdlo_out(a4_wr[1210]));
			radix2 #(.width(width)) rd_st3_1083  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1083]), .rdlo_in(a3_wr[1211]),  .coef_in(coef[472]), .rdup_out(a4_wr[1083]), .rdlo_out(a4_wr[1211]));
			radix2 #(.width(width)) rd_st3_1084  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1084]), .rdlo_in(a3_wr[1212]),  .coef_in(coef[480]), .rdup_out(a4_wr[1084]), .rdlo_out(a4_wr[1212]));
			radix2 #(.width(width)) rd_st3_1085  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1085]), .rdlo_in(a3_wr[1213]),  .coef_in(coef[488]), .rdup_out(a4_wr[1085]), .rdlo_out(a4_wr[1213]));
			radix2 #(.width(width)) rd_st3_1086  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1086]), .rdlo_in(a3_wr[1214]),  .coef_in(coef[496]), .rdup_out(a4_wr[1086]), .rdlo_out(a4_wr[1214]));
			radix2 #(.width(width)) rd_st3_1087  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1087]), .rdlo_in(a3_wr[1215]),  .coef_in(coef[504]), .rdup_out(a4_wr[1087]), .rdlo_out(a4_wr[1215]));
			radix2 #(.width(width)) rd_st3_1088  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1088]), .rdlo_in(a3_wr[1216]),  .coef_in(coef[512]), .rdup_out(a4_wr[1088]), .rdlo_out(a4_wr[1216]));
			radix2 #(.width(width)) rd_st3_1089  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1089]), .rdlo_in(a3_wr[1217]),  .coef_in(coef[520]), .rdup_out(a4_wr[1089]), .rdlo_out(a4_wr[1217]));
			radix2 #(.width(width)) rd_st3_1090  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1090]), .rdlo_in(a3_wr[1218]),  .coef_in(coef[528]), .rdup_out(a4_wr[1090]), .rdlo_out(a4_wr[1218]));
			radix2 #(.width(width)) rd_st3_1091  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1091]), .rdlo_in(a3_wr[1219]),  .coef_in(coef[536]), .rdup_out(a4_wr[1091]), .rdlo_out(a4_wr[1219]));
			radix2 #(.width(width)) rd_st3_1092  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1092]), .rdlo_in(a3_wr[1220]),  .coef_in(coef[544]), .rdup_out(a4_wr[1092]), .rdlo_out(a4_wr[1220]));
			radix2 #(.width(width)) rd_st3_1093  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1093]), .rdlo_in(a3_wr[1221]),  .coef_in(coef[552]), .rdup_out(a4_wr[1093]), .rdlo_out(a4_wr[1221]));
			radix2 #(.width(width)) rd_st3_1094  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1094]), .rdlo_in(a3_wr[1222]),  .coef_in(coef[560]), .rdup_out(a4_wr[1094]), .rdlo_out(a4_wr[1222]));
			radix2 #(.width(width)) rd_st3_1095  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1095]), .rdlo_in(a3_wr[1223]),  .coef_in(coef[568]), .rdup_out(a4_wr[1095]), .rdlo_out(a4_wr[1223]));
			radix2 #(.width(width)) rd_st3_1096  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1096]), .rdlo_in(a3_wr[1224]),  .coef_in(coef[576]), .rdup_out(a4_wr[1096]), .rdlo_out(a4_wr[1224]));
			radix2 #(.width(width)) rd_st3_1097  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1097]), .rdlo_in(a3_wr[1225]),  .coef_in(coef[584]), .rdup_out(a4_wr[1097]), .rdlo_out(a4_wr[1225]));
			radix2 #(.width(width)) rd_st3_1098  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1098]), .rdlo_in(a3_wr[1226]),  .coef_in(coef[592]), .rdup_out(a4_wr[1098]), .rdlo_out(a4_wr[1226]));
			radix2 #(.width(width)) rd_st3_1099  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1099]), .rdlo_in(a3_wr[1227]),  .coef_in(coef[600]), .rdup_out(a4_wr[1099]), .rdlo_out(a4_wr[1227]));
			radix2 #(.width(width)) rd_st3_1100  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1100]), .rdlo_in(a3_wr[1228]),  .coef_in(coef[608]), .rdup_out(a4_wr[1100]), .rdlo_out(a4_wr[1228]));
			radix2 #(.width(width)) rd_st3_1101  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1101]), .rdlo_in(a3_wr[1229]),  .coef_in(coef[616]), .rdup_out(a4_wr[1101]), .rdlo_out(a4_wr[1229]));
			radix2 #(.width(width)) rd_st3_1102  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1102]), .rdlo_in(a3_wr[1230]),  .coef_in(coef[624]), .rdup_out(a4_wr[1102]), .rdlo_out(a4_wr[1230]));
			radix2 #(.width(width)) rd_st3_1103  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1103]), .rdlo_in(a3_wr[1231]),  .coef_in(coef[632]), .rdup_out(a4_wr[1103]), .rdlo_out(a4_wr[1231]));
			radix2 #(.width(width)) rd_st3_1104  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1104]), .rdlo_in(a3_wr[1232]),  .coef_in(coef[640]), .rdup_out(a4_wr[1104]), .rdlo_out(a4_wr[1232]));
			radix2 #(.width(width)) rd_st3_1105  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1105]), .rdlo_in(a3_wr[1233]),  .coef_in(coef[648]), .rdup_out(a4_wr[1105]), .rdlo_out(a4_wr[1233]));
			radix2 #(.width(width)) rd_st3_1106  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1106]), .rdlo_in(a3_wr[1234]),  .coef_in(coef[656]), .rdup_out(a4_wr[1106]), .rdlo_out(a4_wr[1234]));
			radix2 #(.width(width)) rd_st3_1107  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1107]), .rdlo_in(a3_wr[1235]),  .coef_in(coef[664]), .rdup_out(a4_wr[1107]), .rdlo_out(a4_wr[1235]));
			radix2 #(.width(width)) rd_st3_1108  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1108]), .rdlo_in(a3_wr[1236]),  .coef_in(coef[672]), .rdup_out(a4_wr[1108]), .rdlo_out(a4_wr[1236]));
			radix2 #(.width(width)) rd_st3_1109  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1109]), .rdlo_in(a3_wr[1237]),  .coef_in(coef[680]), .rdup_out(a4_wr[1109]), .rdlo_out(a4_wr[1237]));
			radix2 #(.width(width)) rd_st3_1110  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1110]), .rdlo_in(a3_wr[1238]),  .coef_in(coef[688]), .rdup_out(a4_wr[1110]), .rdlo_out(a4_wr[1238]));
			radix2 #(.width(width)) rd_st3_1111  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1111]), .rdlo_in(a3_wr[1239]),  .coef_in(coef[696]), .rdup_out(a4_wr[1111]), .rdlo_out(a4_wr[1239]));
			radix2 #(.width(width)) rd_st3_1112  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1112]), .rdlo_in(a3_wr[1240]),  .coef_in(coef[704]), .rdup_out(a4_wr[1112]), .rdlo_out(a4_wr[1240]));
			radix2 #(.width(width)) rd_st3_1113  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1113]), .rdlo_in(a3_wr[1241]),  .coef_in(coef[712]), .rdup_out(a4_wr[1113]), .rdlo_out(a4_wr[1241]));
			radix2 #(.width(width)) rd_st3_1114  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1114]), .rdlo_in(a3_wr[1242]),  .coef_in(coef[720]), .rdup_out(a4_wr[1114]), .rdlo_out(a4_wr[1242]));
			radix2 #(.width(width)) rd_st3_1115  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1115]), .rdlo_in(a3_wr[1243]),  .coef_in(coef[728]), .rdup_out(a4_wr[1115]), .rdlo_out(a4_wr[1243]));
			radix2 #(.width(width)) rd_st3_1116  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1116]), .rdlo_in(a3_wr[1244]),  .coef_in(coef[736]), .rdup_out(a4_wr[1116]), .rdlo_out(a4_wr[1244]));
			radix2 #(.width(width)) rd_st3_1117  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1117]), .rdlo_in(a3_wr[1245]),  .coef_in(coef[744]), .rdup_out(a4_wr[1117]), .rdlo_out(a4_wr[1245]));
			radix2 #(.width(width)) rd_st3_1118  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1118]), .rdlo_in(a3_wr[1246]),  .coef_in(coef[752]), .rdup_out(a4_wr[1118]), .rdlo_out(a4_wr[1246]));
			radix2 #(.width(width)) rd_st3_1119  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1119]), .rdlo_in(a3_wr[1247]),  .coef_in(coef[760]), .rdup_out(a4_wr[1119]), .rdlo_out(a4_wr[1247]));
			radix2 #(.width(width)) rd_st3_1120  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1120]), .rdlo_in(a3_wr[1248]),  .coef_in(coef[768]), .rdup_out(a4_wr[1120]), .rdlo_out(a4_wr[1248]));
			radix2 #(.width(width)) rd_st3_1121  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1121]), .rdlo_in(a3_wr[1249]),  .coef_in(coef[776]), .rdup_out(a4_wr[1121]), .rdlo_out(a4_wr[1249]));
			radix2 #(.width(width)) rd_st3_1122  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1122]), .rdlo_in(a3_wr[1250]),  .coef_in(coef[784]), .rdup_out(a4_wr[1122]), .rdlo_out(a4_wr[1250]));
			radix2 #(.width(width)) rd_st3_1123  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1123]), .rdlo_in(a3_wr[1251]),  .coef_in(coef[792]), .rdup_out(a4_wr[1123]), .rdlo_out(a4_wr[1251]));
			radix2 #(.width(width)) rd_st3_1124  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1124]), .rdlo_in(a3_wr[1252]),  .coef_in(coef[800]), .rdup_out(a4_wr[1124]), .rdlo_out(a4_wr[1252]));
			radix2 #(.width(width)) rd_st3_1125  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1125]), .rdlo_in(a3_wr[1253]),  .coef_in(coef[808]), .rdup_out(a4_wr[1125]), .rdlo_out(a4_wr[1253]));
			radix2 #(.width(width)) rd_st3_1126  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1126]), .rdlo_in(a3_wr[1254]),  .coef_in(coef[816]), .rdup_out(a4_wr[1126]), .rdlo_out(a4_wr[1254]));
			radix2 #(.width(width)) rd_st3_1127  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1127]), .rdlo_in(a3_wr[1255]),  .coef_in(coef[824]), .rdup_out(a4_wr[1127]), .rdlo_out(a4_wr[1255]));
			radix2 #(.width(width)) rd_st3_1128  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1128]), .rdlo_in(a3_wr[1256]),  .coef_in(coef[832]), .rdup_out(a4_wr[1128]), .rdlo_out(a4_wr[1256]));
			radix2 #(.width(width)) rd_st3_1129  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1129]), .rdlo_in(a3_wr[1257]),  .coef_in(coef[840]), .rdup_out(a4_wr[1129]), .rdlo_out(a4_wr[1257]));
			radix2 #(.width(width)) rd_st3_1130  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1130]), .rdlo_in(a3_wr[1258]),  .coef_in(coef[848]), .rdup_out(a4_wr[1130]), .rdlo_out(a4_wr[1258]));
			radix2 #(.width(width)) rd_st3_1131  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1131]), .rdlo_in(a3_wr[1259]),  .coef_in(coef[856]), .rdup_out(a4_wr[1131]), .rdlo_out(a4_wr[1259]));
			radix2 #(.width(width)) rd_st3_1132  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1132]), .rdlo_in(a3_wr[1260]),  .coef_in(coef[864]), .rdup_out(a4_wr[1132]), .rdlo_out(a4_wr[1260]));
			radix2 #(.width(width)) rd_st3_1133  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1133]), .rdlo_in(a3_wr[1261]),  .coef_in(coef[872]), .rdup_out(a4_wr[1133]), .rdlo_out(a4_wr[1261]));
			radix2 #(.width(width)) rd_st3_1134  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1134]), .rdlo_in(a3_wr[1262]),  .coef_in(coef[880]), .rdup_out(a4_wr[1134]), .rdlo_out(a4_wr[1262]));
			radix2 #(.width(width)) rd_st3_1135  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1135]), .rdlo_in(a3_wr[1263]),  .coef_in(coef[888]), .rdup_out(a4_wr[1135]), .rdlo_out(a4_wr[1263]));
			radix2 #(.width(width)) rd_st3_1136  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1136]), .rdlo_in(a3_wr[1264]),  .coef_in(coef[896]), .rdup_out(a4_wr[1136]), .rdlo_out(a4_wr[1264]));
			radix2 #(.width(width)) rd_st3_1137  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1137]), .rdlo_in(a3_wr[1265]),  .coef_in(coef[904]), .rdup_out(a4_wr[1137]), .rdlo_out(a4_wr[1265]));
			radix2 #(.width(width)) rd_st3_1138  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1138]), .rdlo_in(a3_wr[1266]),  .coef_in(coef[912]), .rdup_out(a4_wr[1138]), .rdlo_out(a4_wr[1266]));
			radix2 #(.width(width)) rd_st3_1139  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1139]), .rdlo_in(a3_wr[1267]),  .coef_in(coef[920]), .rdup_out(a4_wr[1139]), .rdlo_out(a4_wr[1267]));
			radix2 #(.width(width)) rd_st3_1140  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1140]), .rdlo_in(a3_wr[1268]),  .coef_in(coef[928]), .rdup_out(a4_wr[1140]), .rdlo_out(a4_wr[1268]));
			radix2 #(.width(width)) rd_st3_1141  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1141]), .rdlo_in(a3_wr[1269]),  .coef_in(coef[936]), .rdup_out(a4_wr[1141]), .rdlo_out(a4_wr[1269]));
			radix2 #(.width(width)) rd_st3_1142  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1142]), .rdlo_in(a3_wr[1270]),  .coef_in(coef[944]), .rdup_out(a4_wr[1142]), .rdlo_out(a4_wr[1270]));
			radix2 #(.width(width)) rd_st3_1143  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1143]), .rdlo_in(a3_wr[1271]),  .coef_in(coef[952]), .rdup_out(a4_wr[1143]), .rdlo_out(a4_wr[1271]));
			radix2 #(.width(width)) rd_st3_1144  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1144]), .rdlo_in(a3_wr[1272]),  .coef_in(coef[960]), .rdup_out(a4_wr[1144]), .rdlo_out(a4_wr[1272]));
			radix2 #(.width(width)) rd_st3_1145  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1145]), .rdlo_in(a3_wr[1273]),  .coef_in(coef[968]), .rdup_out(a4_wr[1145]), .rdlo_out(a4_wr[1273]));
			radix2 #(.width(width)) rd_st3_1146  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1146]), .rdlo_in(a3_wr[1274]),  .coef_in(coef[976]), .rdup_out(a4_wr[1146]), .rdlo_out(a4_wr[1274]));
			radix2 #(.width(width)) rd_st3_1147  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1147]), .rdlo_in(a3_wr[1275]),  .coef_in(coef[984]), .rdup_out(a4_wr[1147]), .rdlo_out(a4_wr[1275]));
			radix2 #(.width(width)) rd_st3_1148  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1148]), .rdlo_in(a3_wr[1276]),  .coef_in(coef[992]), .rdup_out(a4_wr[1148]), .rdlo_out(a4_wr[1276]));
			radix2 #(.width(width)) rd_st3_1149  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1149]), .rdlo_in(a3_wr[1277]),  .coef_in(coef[1000]), .rdup_out(a4_wr[1149]), .rdlo_out(a4_wr[1277]));
			radix2 #(.width(width)) rd_st3_1150  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1150]), .rdlo_in(a3_wr[1278]),  .coef_in(coef[1008]), .rdup_out(a4_wr[1150]), .rdlo_out(a4_wr[1278]));
			radix2 #(.width(width)) rd_st3_1151  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1151]), .rdlo_in(a3_wr[1279]),  .coef_in(coef[1016]), .rdup_out(a4_wr[1151]), .rdlo_out(a4_wr[1279]));
			radix2 #(.width(width)) rd_st3_1280  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1280]), .rdlo_in(a3_wr[1408]),  .coef_in(coef[0]), .rdup_out(a4_wr[1280]), .rdlo_out(a4_wr[1408]));
			radix2 #(.width(width)) rd_st3_1281  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1281]), .rdlo_in(a3_wr[1409]),  .coef_in(coef[8]), .rdup_out(a4_wr[1281]), .rdlo_out(a4_wr[1409]));
			radix2 #(.width(width)) rd_st3_1282  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1282]), .rdlo_in(a3_wr[1410]),  .coef_in(coef[16]), .rdup_out(a4_wr[1282]), .rdlo_out(a4_wr[1410]));
			radix2 #(.width(width)) rd_st3_1283  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1283]), .rdlo_in(a3_wr[1411]),  .coef_in(coef[24]), .rdup_out(a4_wr[1283]), .rdlo_out(a4_wr[1411]));
			radix2 #(.width(width)) rd_st3_1284  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1284]), .rdlo_in(a3_wr[1412]),  .coef_in(coef[32]), .rdup_out(a4_wr[1284]), .rdlo_out(a4_wr[1412]));
			radix2 #(.width(width)) rd_st3_1285  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1285]), .rdlo_in(a3_wr[1413]),  .coef_in(coef[40]), .rdup_out(a4_wr[1285]), .rdlo_out(a4_wr[1413]));
			radix2 #(.width(width)) rd_st3_1286  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1286]), .rdlo_in(a3_wr[1414]),  .coef_in(coef[48]), .rdup_out(a4_wr[1286]), .rdlo_out(a4_wr[1414]));
			radix2 #(.width(width)) rd_st3_1287  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1287]), .rdlo_in(a3_wr[1415]),  .coef_in(coef[56]), .rdup_out(a4_wr[1287]), .rdlo_out(a4_wr[1415]));
			radix2 #(.width(width)) rd_st3_1288  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1288]), .rdlo_in(a3_wr[1416]),  .coef_in(coef[64]), .rdup_out(a4_wr[1288]), .rdlo_out(a4_wr[1416]));
			radix2 #(.width(width)) rd_st3_1289  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1289]), .rdlo_in(a3_wr[1417]),  .coef_in(coef[72]), .rdup_out(a4_wr[1289]), .rdlo_out(a4_wr[1417]));
			radix2 #(.width(width)) rd_st3_1290  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1290]), .rdlo_in(a3_wr[1418]),  .coef_in(coef[80]), .rdup_out(a4_wr[1290]), .rdlo_out(a4_wr[1418]));
			radix2 #(.width(width)) rd_st3_1291  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1291]), .rdlo_in(a3_wr[1419]),  .coef_in(coef[88]), .rdup_out(a4_wr[1291]), .rdlo_out(a4_wr[1419]));
			radix2 #(.width(width)) rd_st3_1292  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1292]), .rdlo_in(a3_wr[1420]),  .coef_in(coef[96]), .rdup_out(a4_wr[1292]), .rdlo_out(a4_wr[1420]));
			radix2 #(.width(width)) rd_st3_1293  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1293]), .rdlo_in(a3_wr[1421]),  .coef_in(coef[104]), .rdup_out(a4_wr[1293]), .rdlo_out(a4_wr[1421]));
			radix2 #(.width(width)) rd_st3_1294  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1294]), .rdlo_in(a3_wr[1422]),  .coef_in(coef[112]), .rdup_out(a4_wr[1294]), .rdlo_out(a4_wr[1422]));
			radix2 #(.width(width)) rd_st3_1295  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1295]), .rdlo_in(a3_wr[1423]),  .coef_in(coef[120]), .rdup_out(a4_wr[1295]), .rdlo_out(a4_wr[1423]));
			radix2 #(.width(width)) rd_st3_1296  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1296]), .rdlo_in(a3_wr[1424]),  .coef_in(coef[128]), .rdup_out(a4_wr[1296]), .rdlo_out(a4_wr[1424]));
			radix2 #(.width(width)) rd_st3_1297  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1297]), .rdlo_in(a3_wr[1425]),  .coef_in(coef[136]), .rdup_out(a4_wr[1297]), .rdlo_out(a4_wr[1425]));
			radix2 #(.width(width)) rd_st3_1298  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1298]), .rdlo_in(a3_wr[1426]),  .coef_in(coef[144]), .rdup_out(a4_wr[1298]), .rdlo_out(a4_wr[1426]));
			radix2 #(.width(width)) rd_st3_1299  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1299]), .rdlo_in(a3_wr[1427]),  .coef_in(coef[152]), .rdup_out(a4_wr[1299]), .rdlo_out(a4_wr[1427]));
			radix2 #(.width(width)) rd_st3_1300  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1300]), .rdlo_in(a3_wr[1428]),  .coef_in(coef[160]), .rdup_out(a4_wr[1300]), .rdlo_out(a4_wr[1428]));
			radix2 #(.width(width)) rd_st3_1301  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1301]), .rdlo_in(a3_wr[1429]),  .coef_in(coef[168]), .rdup_out(a4_wr[1301]), .rdlo_out(a4_wr[1429]));
			radix2 #(.width(width)) rd_st3_1302  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1302]), .rdlo_in(a3_wr[1430]),  .coef_in(coef[176]), .rdup_out(a4_wr[1302]), .rdlo_out(a4_wr[1430]));
			radix2 #(.width(width)) rd_st3_1303  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1303]), .rdlo_in(a3_wr[1431]),  .coef_in(coef[184]), .rdup_out(a4_wr[1303]), .rdlo_out(a4_wr[1431]));
			radix2 #(.width(width)) rd_st3_1304  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1304]), .rdlo_in(a3_wr[1432]),  .coef_in(coef[192]), .rdup_out(a4_wr[1304]), .rdlo_out(a4_wr[1432]));
			radix2 #(.width(width)) rd_st3_1305  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1305]), .rdlo_in(a3_wr[1433]),  .coef_in(coef[200]), .rdup_out(a4_wr[1305]), .rdlo_out(a4_wr[1433]));
			radix2 #(.width(width)) rd_st3_1306  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1306]), .rdlo_in(a3_wr[1434]),  .coef_in(coef[208]), .rdup_out(a4_wr[1306]), .rdlo_out(a4_wr[1434]));
			radix2 #(.width(width)) rd_st3_1307  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1307]), .rdlo_in(a3_wr[1435]),  .coef_in(coef[216]), .rdup_out(a4_wr[1307]), .rdlo_out(a4_wr[1435]));
			radix2 #(.width(width)) rd_st3_1308  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1308]), .rdlo_in(a3_wr[1436]),  .coef_in(coef[224]), .rdup_out(a4_wr[1308]), .rdlo_out(a4_wr[1436]));
			radix2 #(.width(width)) rd_st3_1309  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1309]), .rdlo_in(a3_wr[1437]),  .coef_in(coef[232]), .rdup_out(a4_wr[1309]), .rdlo_out(a4_wr[1437]));
			radix2 #(.width(width)) rd_st3_1310  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1310]), .rdlo_in(a3_wr[1438]),  .coef_in(coef[240]), .rdup_out(a4_wr[1310]), .rdlo_out(a4_wr[1438]));
			radix2 #(.width(width)) rd_st3_1311  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1311]), .rdlo_in(a3_wr[1439]),  .coef_in(coef[248]), .rdup_out(a4_wr[1311]), .rdlo_out(a4_wr[1439]));
			radix2 #(.width(width)) rd_st3_1312  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1312]), .rdlo_in(a3_wr[1440]),  .coef_in(coef[256]), .rdup_out(a4_wr[1312]), .rdlo_out(a4_wr[1440]));
			radix2 #(.width(width)) rd_st3_1313  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1313]), .rdlo_in(a3_wr[1441]),  .coef_in(coef[264]), .rdup_out(a4_wr[1313]), .rdlo_out(a4_wr[1441]));
			radix2 #(.width(width)) rd_st3_1314  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1314]), .rdlo_in(a3_wr[1442]),  .coef_in(coef[272]), .rdup_out(a4_wr[1314]), .rdlo_out(a4_wr[1442]));
			radix2 #(.width(width)) rd_st3_1315  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1315]), .rdlo_in(a3_wr[1443]),  .coef_in(coef[280]), .rdup_out(a4_wr[1315]), .rdlo_out(a4_wr[1443]));
			radix2 #(.width(width)) rd_st3_1316  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1316]), .rdlo_in(a3_wr[1444]),  .coef_in(coef[288]), .rdup_out(a4_wr[1316]), .rdlo_out(a4_wr[1444]));
			radix2 #(.width(width)) rd_st3_1317  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1317]), .rdlo_in(a3_wr[1445]),  .coef_in(coef[296]), .rdup_out(a4_wr[1317]), .rdlo_out(a4_wr[1445]));
			radix2 #(.width(width)) rd_st3_1318  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1318]), .rdlo_in(a3_wr[1446]),  .coef_in(coef[304]), .rdup_out(a4_wr[1318]), .rdlo_out(a4_wr[1446]));
			radix2 #(.width(width)) rd_st3_1319  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1319]), .rdlo_in(a3_wr[1447]),  .coef_in(coef[312]), .rdup_out(a4_wr[1319]), .rdlo_out(a4_wr[1447]));
			radix2 #(.width(width)) rd_st3_1320  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1320]), .rdlo_in(a3_wr[1448]),  .coef_in(coef[320]), .rdup_out(a4_wr[1320]), .rdlo_out(a4_wr[1448]));
			radix2 #(.width(width)) rd_st3_1321  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1321]), .rdlo_in(a3_wr[1449]),  .coef_in(coef[328]), .rdup_out(a4_wr[1321]), .rdlo_out(a4_wr[1449]));
			radix2 #(.width(width)) rd_st3_1322  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1322]), .rdlo_in(a3_wr[1450]),  .coef_in(coef[336]), .rdup_out(a4_wr[1322]), .rdlo_out(a4_wr[1450]));
			radix2 #(.width(width)) rd_st3_1323  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1323]), .rdlo_in(a3_wr[1451]),  .coef_in(coef[344]), .rdup_out(a4_wr[1323]), .rdlo_out(a4_wr[1451]));
			radix2 #(.width(width)) rd_st3_1324  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1324]), .rdlo_in(a3_wr[1452]),  .coef_in(coef[352]), .rdup_out(a4_wr[1324]), .rdlo_out(a4_wr[1452]));
			radix2 #(.width(width)) rd_st3_1325  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1325]), .rdlo_in(a3_wr[1453]),  .coef_in(coef[360]), .rdup_out(a4_wr[1325]), .rdlo_out(a4_wr[1453]));
			radix2 #(.width(width)) rd_st3_1326  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1326]), .rdlo_in(a3_wr[1454]),  .coef_in(coef[368]), .rdup_out(a4_wr[1326]), .rdlo_out(a4_wr[1454]));
			radix2 #(.width(width)) rd_st3_1327  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1327]), .rdlo_in(a3_wr[1455]),  .coef_in(coef[376]), .rdup_out(a4_wr[1327]), .rdlo_out(a4_wr[1455]));
			radix2 #(.width(width)) rd_st3_1328  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1328]), .rdlo_in(a3_wr[1456]),  .coef_in(coef[384]), .rdup_out(a4_wr[1328]), .rdlo_out(a4_wr[1456]));
			radix2 #(.width(width)) rd_st3_1329  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1329]), .rdlo_in(a3_wr[1457]),  .coef_in(coef[392]), .rdup_out(a4_wr[1329]), .rdlo_out(a4_wr[1457]));
			radix2 #(.width(width)) rd_st3_1330  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1330]), .rdlo_in(a3_wr[1458]),  .coef_in(coef[400]), .rdup_out(a4_wr[1330]), .rdlo_out(a4_wr[1458]));
			radix2 #(.width(width)) rd_st3_1331  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1331]), .rdlo_in(a3_wr[1459]),  .coef_in(coef[408]), .rdup_out(a4_wr[1331]), .rdlo_out(a4_wr[1459]));
			radix2 #(.width(width)) rd_st3_1332  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1332]), .rdlo_in(a3_wr[1460]),  .coef_in(coef[416]), .rdup_out(a4_wr[1332]), .rdlo_out(a4_wr[1460]));
			radix2 #(.width(width)) rd_st3_1333  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1333]), .rdlo_in(a3_wr[1461]),  .coef_in(coef[424]), .rdup_out(a4_wr[1333]), .rdlo_out(a4_wr[1461]));
			radix2 #(.width(width)) rd_st3_1334  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1334]), .rdlo_in(a3_wr[1462]),  .coef_in(coef[432]), .rdup_out(a4_wr[1334]), .rdlo_out(a4_wr[1462]));
			radix2 #(.width(width)) rd_st3_1335  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1335]), .rdlo_in(a3_wr[1463]),  .coef_in(coef[440]), .rdup_out(a4_wr[1335]), .rdlo_out(a4_wr[1463]));
			radix2 #(.width(width)) rd_st3_1336  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1336]), .rdlo_in(a3_wr[1464]),  .coef_in(coef[448]), .rdup_out(a4_wr[1336]), .rdlo_out(a4_wr[1464]));
			radix2 #(.width(width)) rd_st3_1337  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1337]), .rdlo_in(a3_wr[1465]),  .coef_in(coef[456]), .rdup_out(a4_wr[1337]), .rdlo_out(a4_wr[1465]));
			radix2 #(.width(width)) rd_st3_1338  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1338]), .rdlo_in(a3_wr[1466]),  .coef_in(coef[464]), .rdup_out(a4_wr[1338]), .rdlo_out(a4_wr[1466]));
			radix2 #(.width(width)) rd_st3_1339  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1339]), .rdlo_in(a3_wr[1467]),  .coef_in(coef[472]), .rdup_out(a4_wr[1339]), .rdlo_out(a4_wr[1467]));
			radix2 #(.width(width)) rd_st3_1340  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1340]), .rdlo_in(a3_wr[1468]),  .coef_in(coef[480]), .rdup_out(a4_wr[1340]), .rdlo_out(a4_wr[1468]));
			radix2 #(.width(width)) rd_st3_1341  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1341]), .rdlo_in(a3_wr[1469]),  .coef_in(coef[488]), .rdup_out(a4_wr[1341]), .rdlo_out(a4_wr[1469]));
			radix2 #(.width(width)) rd_st3_1342  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1342]), .rdlo_in(a3_wr[1470]),  .coef_in(coef[496]), .rdup_out(a4_wr[1342]), .rdlo_out(a4_wr[1470]));
			radix2 #(.width(width)) rd_st3_1343  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1343]), .rdlo_in(a3_wr[1471]),  .coef_in(coef[504]), .rdup_out(a4_wr[1343]), .rdlo_out(a4_wr[1471]));
			radix2 #(.width(width)) rd_st3_1344  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1344]), .rdlo_in(a3_wr[1472]),  .coef_in(coef[512]), .rdup_out(a4_wr[1344]), .rdlo_out(a4_wr[1472]));
			radix2 #(.width(width)) rd_st3_1345  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1345]), .rdlo_in(a3_wr[1473]),  .coef_in(coef[520]), .rdup_out(a4_wr[1345]), .rdlo_out(a4_wr[1473]));
			radix2 #(.width(width)) rd_st3_1346  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1346]), .rdlo_in(a3_wr[1474]),  .coef_in(coef[528]), .rdup_out(a4_wr[1346]), .rdlo_out(a4_wr[1474]));
			radix2 #(.width(width)) rd_st3_1347  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1347]), .rdlo_in(a3_wr[1475]),  .coef_in(coef[536]), .rdup_out(a4_wr[1347]), .rdlo_out(a4_wr[1475]));
			radix2 #(.width(width)) rd_st3_1348  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1348]), .rdlo_in(a3_wr[1476]),  .coef_in(coef[544]), .rdup_out(a4_wr[1348]), .rdlo_out(a4_wr[1476]));
			radix2 #(.width(width)) rd_st3_1349  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1349]), .rdlo_in(a3_wr[1477]),  .coef_in(coef[552]), .rdup_out(a4_wr[1349]), .rdlo_out(a4_wr[1477]));
			radix2 #(.width(width)) rd_st3_1350  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1350]), .rdlo_in(a3_wr[1478]),  .coef_in(coef[560]), .rdup_out(a4_wr[1350]), .rdlo_out(a4_wr[1478]));
			radix2 #(.width(width)) rd_st3_1351  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1351]), .rdlo_in(a3_wr[1479]),  .coef_in(coef[568]), .rdup_out(a4_wr[1351]), .rdlo_out(a4_wr[1479]));
			radix2 #(.width(width)) rd_st3_1352  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1352]), .rdlo_in(a3_wr[1480]),  .coef_in(coef[576]), .rdup_out(a4_wr[1352]), .rdlo_out(a4_wr[1480]));
			radix2 #(.width(width)) rd_st3_1353  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1353]), .rdlo_in(a3_wr[1481]),  .coef_in(coef[584]), .rdup_out(a4_wr[1353]), .rdlo_out(a4_wr[1481]));
			radix2 #(.width(width)) rd_st3_1354  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1354]), .rdlo_in(a3_wr[1482]),  .coef_in(coef[592]), .rdup_out(a4_wr[1354]), .rdlo_out(a4_wr[1482]));
			radix2 #(.width(width)) rd_st3_1355  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1355]), .rdlo_in(a3_wr[1483]),  .coef_in(coef[600]), .rdup_out(a4_wr[1355]), .rdlo_out(a4_wr[1483]));
			radix2 #(.width(width)) rd_st3_1356  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1356]), .rdlo_in(a3_wr[1484]),  .coef_in(coef[608]), .rdup_out(a4_wr[1356]), .rdlo_out(a4_wr[1484]));
			radix2 #(.width(width)) rd_st3_1357  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1357]), .rdlo_in(a3_wr[1485]),  .coef_in(coef[616]), .rdup_out(a4_wr[1357]), .rdlo_out(a4_wr[1485]));
			radix2 #(.width(width)) rd_st3_1358  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1358]), .rdlo_in(a3_wr[1486]),  .coef_in(coef[624]), .rdup_out(a4_wr[1358]), .rdlo_out(a4_wr[1486]));
			radix2 #(.width(width)) rd_st3_1359  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1359]), .rdlo_in(a3_wr[1487]),  .coef_in(coef[632]), .rdup_out(a4_wr[1359]), .rdlo_out(a4_wr[1487]));
			radix2 #(.width(width)) rd_st3_1360  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1360]), .rdlo_in(a3_wr[1488]),  .coef_in(coef[640]), .rdup_out(a4_wr[1360]), .rdlo_out(a4_wr[1488]));
			radix2 #(.width(width)) rd_st3_1361  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1361]), .rdlo_in(a3_wr[1489]),  .coef_in(coef[648]), .rdup_out(a4_wr[1361]), .rdlo_out(a4_wr[1489]));
			radix2 #(.width(width)) rd_st3_1362  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1362]), .rdlo_in(a3_wr[1490]),  .coef_in(coef[656]), .rdup_out(a4_wr[1362]), .rdlo_out(a4_wr[1490]));
			radix2 #(.width(width)) rd_st3_1363  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1363]), .rdlo_in(a3_wr[1491]),  .coef_in(coef[664]), .rdup_out(a4_wr[1363]), .rdlo_out(a4_wr[1491]));
			radix2 #(.width(width)) rd_st3_1364  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1364]), .rdlo_in(a3_wr[1492]),  .coef_in(coef[672]), .rdup_out(a4_wr[1364]), .rdlo_out(a4_wr[1492]));
			radix2 #(.width(width)) rd_st3_1365  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1365]), .rdlo_in(a3_wr[1493]),  .coef_in(coef[680]), .rdup_out(a4_wr[1365]), .rdlo_out(a4_wr[1493]));
			radix2 #(.width(width)) rd_st3_1366  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1366]), .rdlo_in(a3_wr[1494]),  .coef_in(coef[688]), .rdup_out(a4_wr[1366]), .rdlo_out(a4_wr[1494]));
			radix2 #(.width(width)) rd_st3_1367  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1367]), .rdlo_in(a3_wr[1495]),  .coef_in(coef[696]), .rdup_out(a4_wr[1367]), .rdlo_out(a4_wr[1495]));
			radix2 #(.width(width)) rd_st3_1368  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1368]), .rdlo_in(a3_wr[1496]),  .coef_in(coef[704]), .rdup_out(a4_wr[1368]), .rdlo_out(a4_wr[1496]));
			radix2 #(.width(width)) rd_st3_1369  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1369]), .rdlo_in(a3_wr[1497]),  .coef_in(coef[712]), .rdup_out(a4_wr[1369]), .rdlo_out(a4_wr[1497]));
			radix2 #(.width(width)) rd_st3_1370  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1370]), .rdlo_in(a3_wr[1498]),  .coef_in(coef[720]), .rdup_out(a4_wr[1370]), .rdlo_out(a4_wr[1498]));
			radix2 #(.width(width)) rd_st3_1371  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1371]), .rdlo_in(a3_wr[1499]),  .coef_in(coef[728]), .rdup_out(a4_wr[1371]), .rdlo_out(a4_wr[1499]));
			radix2 #(.width(width)) rd_st3_1372  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1372]), .rdlo_in(a3_wr[1500]),  .coef_in(coef[736]), .rdup_out(a4_wr[1372]), .rdlo_out(a4_wr[1500]));
			radix2 #(.width(width)) rd_st3_1373  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1373]), .rdlo_in(a3_wr[1501]),  .coef_in(coef[744]), .rdup_out(a4_wr[1373]), .rdlo_out(a4_wr[1501]));
			radix2 #(.width(width)) rd_st3_1374  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1374]), .rdlo_in(a3_wr[1502]),  .coef_in(coef[752]), .rdup_out(a4_wr[1374]), .rdlo_out(a4_wr[1502]));
			radix2 #(.width(width)) rd_st3_1375  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1375]), .rdlo_in(a3_wr[1503]),  .coef_in(coef[760]), .rdup_out(a4_wr[1375]), .rdlo_out(a4_wr[1503]));
			radix2 #(.width(width)) rd_st3_1376  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1376]), .rdlo_in(a3_wr[1504]),  .coef_in(coef[768]), .rdup_out(a4_wr[1376]), .rdlo_out(a4_wr[1504]));
			radix2 #(.width(width)) rd_st3_1377  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1377]), .rdlo_in(a3_wr[1505]),  .coef_in(coef[776]), .rdup_out(a4_wr[1377]), .rdlo_out(a4_wr[1505]));
			radix2 #(.width(width)) rd_st3_1378  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1378]), .rdlo_in(a3_wr[1506]),  .coef_in(coef[784]), .rdup_out(a4_wr[1378]), .rdlo_out(a4_wr[1506]));
			radix2 #(.width(width)) rd_st3_1379  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1379]), .rdlo_in(a3_wr[1507]),  .coef_in(coef[792]), .rdup_out(a4_wr[1379]), .rdlo_out(a4_wr[1507]));
			radix2 #(.width(width)) rd_st3_1380  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1380]), .rdlo_in(a3_wr[1508]),  .coef_in(coef[800]), .rdup_out(a4_wr[1380]), .rdlo_out(a4_wr[1508]));
			radix2 #(.width(width)) rd_st3_1381  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1381]), .rdlo_in(a3_wr[1509]),  .coef_in(coef[808]), .rdup_out(a4_wr[1381]), .rdlo_out(a4_wr[1509]));
			radix2 #(.width(width)) rd_st3_1382  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1382]), .rdlo_in(a3_wr[1510]),  .coef_in(coef[816]), .rdup_out(a4_wr[1382]), .rdlo_out(a4_wr[1510]));
			radix2 #(.width(width)) rd_st3_1383  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1383]), .rdlo_in(a3_wr[1511]),  .coef_in(coef[824]), .rdup_out(a4_wr[1383]), .rdlo_out(a4_wr[1511]));
			radix2 #(.width(width)) rd_st3_1384  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1384]), .rdlo_in(a3_wr[1512]),  .coef_in(coef[832]), .rdup_out(a4_wr[1384]), .rdlo_out(a4_wr[1512]));
			radix2 #(.width(width)) rd_st3_1385  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1385]), .rdlo_in(a3_wr[1513]),  .coef_in(coef[840]), .rdup_out(a4_wr[1385]), .rdlo_out(a4_wr[1513]));
			radix2 #(.width(width)) rd_st3_1386  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1386]), .rdlo_in(a3_wr[1514]),  .coef_in(coef[848]), .rdup_out(a4_wr[1386]), .rdlo_out(a4_wr[1514]));
			radix2 #(.width(width)) rd_st3_1387  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1387]), .rdlo_in(a3_wr[1515]),  .coef_in(coef[856]), .rdup_out(a4_wr[1387]), .rdlo_out(a4_wr[1515]));
			radix2 #(.width(width)) rd_st3_1388  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1388]), .rdlo_in(a3_wr[1516]),  .coef_in(coef[864]), .rdup_out(a4_wr[1388]), .rdlo_out(a4_wr[1516]));
			radix2 #(.width(width)) rd_st3_1389  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1389]), .rdlo_in(a3_wr[1517]),  .coef_in(coef[872]), .rdup_out(a4_wr[1389]), .rdlo_out(a4_wr[1517]));
			radix2 #(.width(width)) rd_st3_1390  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1390]), .rdlo_in(a3_wr[1518]),  .coef_in(coef[880]), .rdup_out(a4_wr[1390]), .rdlo_out(a4_wr[1518]));
			radix2 #(.width(width)) rd_st3_1391  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1391]), .rdlo_in(a3_wr[1519]),  .coef_in(coef[888]), .rdup_out(a4_wr[1391]), .rdlo_out(a4_wr[1519]));
			radix2 #(.width(width)) rd_st3_1392  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1392]), .rdlo_in(a3_wr[1520]),  .coef_in(coef[896]), .rdup_out(a4_wr[1392]), .rdlo_out(a4_wr[1520]));
			radix2 #(.width(width)) rd_st3_1393  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1393]), .rdlo_in(a3_wr[1521]),  .coef_in(coef[904]), .rdup_out(a4_wr[1393]), .rdlo_out(a4_wr[1521]));
			radix2 #(.width(width)) rd_st3_1394  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1394]), .rdlo_in(a3_wr[1522]),  .coef_in(coef[912]), .rdup_out(a4_wr[1394]), .rdlo_out(a4_wr[1522]));
			radix2 #(.width(width)) rd_st3_1395  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1395]), .rdlo_in(a3_wr[1523]),  .coef_in(coef[920]), .rdup_out(a4_wr[1395]), .rdlo_out(a4_wr[1523]));
			radix2 #(.width(width)) rd_st3_1396  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1396]), .rdlo_in(a3_wr[1524]),  .coef_in(coef[928]), .rdup_out(a4_wr[1396]), .rdlo_out(a4_wr[1524]));
			radix2 #(.width(width)) rd_st3_1397  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1397]), .rdlo_in(a3_wr[1525]),  .coef_in(coef[936]), .rdup_out(a4_wr[1397]), .rdlo_out(a4_wr[1525]));
			radix2 #(.width(width)) rd_st3_1398  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1398]), .rdlo_in(a3_wr[1526]),  .coef_in(coef[944]), .rdup_out(a4_wr[1398]), .rdlo_out(a4_wr[1526]));
			radix2 #(.width(width)) rd_st3_1399  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1399]), .rdlo_in(a3_wr[1527]),  .coef_in(coef[952]), .rdup_out(a4_wr[1399]), .rdlo_out(a4_wr[1527]));
			radix2 #(.width(width)) rd_st3_1400  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1400]), .rdlo_in(a3_wr[1528]),  .coef_in(coef[960]), .rdup_out(a4_wr[1400]), .rdlo_out(a4_wr[1528]));
			radix2 #(.width(width)) rd_st3_1401  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1401]), .rdlo_in(a3_wr[1529]),  .coef_in(coef[968]), .rdup_out(a4_wr[1401]), .rdlo_out(a4_wr[1529]));
			radix2 #(.width(width)) rd_st3_1402  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1402]), .rdlo_in(a3_wr[1530]),  .coef_in(coef[976]), .rdup_out(a4_wr[1402]), .rdlo_out(a4_wr[1530]));
			radix2 #(.width(width)) rd_st3_1403  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1403]), .rdlo_in(a3_wr[1531]),  .coef_in(coef[984]), .rdup_out(a4_wr[1403]), .rdlo_out(a4_wr[1531]));
			radix2 #(.width(width)) rd_st3_1404  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1404]), .rdlo_in(a3_wr[1532]),  .coef_in(coef[992]), .rdup_out(a4_wr[1404]), .rdlo_out(a4_wr[1532]));
			radix2 #(.width(width)) rd_st3_1405  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1405]), .rdlo_in(a3_wr[1533]),  .coef_in(coef[1000]), .rdup_out(a4_wr[1405]), .rdlo_out(a4_wr[1533]));
			radix2 #(.width(width)) rd_st3_1406  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1406]), .rdlo_in(a3_wr[1534]),  .coef_in(coef[1008]), .rdup_out(a4_wr[1406]), .rdlo_out(a4_wr[1534]));
			radix2 #(.width(width)) rd_st3_1407  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1407]), .rdlo_in(a3_wr[1535]),  .coef_in(coef[1016]), .rdup_out(a4_wr[1407]), .rdlo_out(a4_wr[1535]));
			radix2 #(.width(width)) rd_st3_1536  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1536]), .rdlo_in(a3_wr[1664]),  .coef_in(coef[0]), .rdup_out(a4_wr[1536]), .rdlo_out(a4_wr[1664]));
			radix2 #(.width(width)) rd_st3_1537  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1537]), .rdlo_in(a3_wr[1665]),  .coef_in(coef[8]), .rdup_out(a4_wr[1537]), .rdlo_out(a4_wr[1665]));
			radix2 #(.width(width)) rd_st3_1538  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1538]), .rdlo_in(a3_wr[1666]),  .coef_in(coef[16]), .rdup_out(a4_wr[1538]), .rdlo_out(a4_wr[1666]));
			radix2 #(.width(width)) rd_st3_1539  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1539]), .rdlo_in(a3_wr[1667]),  .coef_in(coef[24]), .rdup_out(a4_wr[1539]), .rdlo_out(a4_wr[1667]));
			radix2 #(.width(width)) rd_st3_1540  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1540]), .rdlo_in(a3_wr[1668]),  .coef_in(coef[32]), .rdup_out(a4_wr[1540]), .rdlo_out(a4_wr[1668]));
			radix2 #(.width(width)) rd_st3_1541  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1541]), .rdlo_in(a3_wr[1669]),  .coef_in(coef[40]), .rdup_out(a4_wr[1541]), .rdlo_out(a4_wr[1669]));
			radix2 #(.width(width)) rd_st3_1542  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1542]), .rdlo_in(a3_wr[1670]),  .coef_in(coef[48]), .rdup_out(a4_wr[1542]), .rdlo_out(a4_wr[1670]));
			radix2 #(.width(width)) rd_st3_1543  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1543]), .rdlo_in(a3_wr[1671]),  .coef_in(coef[56]), .rdup_out(a4_wr[1543]), .rdlo_out(a4_wr[1671]));
			radix2 #(.width(width)) rd_st3_1544  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1544]), .rdlo_in(a3_wr[1672]),  .coef_in(coef[64]), .rdup_out(a4_wr[1544]), .rdlo_out(a4_wr[1672]));
			radix2 #(.width(width)) rd_st3_1545  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1545]), .rdlo_in(a3_wr[1673]),  .coef_in(coef[72]), .rdup_out(a4_wr[1545]), .rdlo_out(a4_wr[1673]));
			radix2 #(.width(width)) rd_st3_1546  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1546]), .rdlo_in(a3_wr[1674]),  .coef_in(coef[80]), .rdup_out(a4_wr[1546]), .rdlo_out(a4_wr[1674]));
			radix2 #(.width(width)) rd_st3_1547  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1547]), .rdlo_in(a3_wr[1675]),  .coef_in(coef[88]), .rdup_out(a4_wr[1547]), .rdlo_out(a4_wr[1675]));
			radix2 #(.width(width)) rd_st3_1548  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1548]), .rdlo_in(a3_wr[1676]),  .coef_in(coef[96]), .rdup_out(a4_wr[1548]), .rdlo_out(a4_wr[1676]));
			radix2 #(.width(width)) rd_st3_1549  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1549]), .rdlo_in(a3_wr[1677]),  .coef_in(coef[104]), .rdup_out(a4_wr[1549]), .rdlo_out(a4_wr[1677]));
			radix2 #(.width(width)) rd_st3_1550  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1550]), .rdlo_in(a3_wr[1678]),  .coef_in(coef[112]), .rdup_out(a4_wr[1550]), .rdlo_out(a4_wr[1678]));
			radix2 #(.width(width)) rd_st3_1551  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1551]), .rdlo_in(a3_wr[1679]),  .coef_in(coef[120]), .rdup_out(a4_wr[1551]), .rdlo_out(a4_wr[1679]));
			radix2 #(.width(width)) rd_st3_1552  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1552]), .rdlo_in(a3_wr[1680]),  .coef_in(coef[128]), .rdup_out(a4_wr[1552]), .rdlo_out(a4_wr[1680]));
			radix2 #(.width(width)) rd_st3_1553  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1553]), .rdlo_in(a3_wr[1681]),  .coef_in(coef[136]), .rdup_out(a4_wr[1553]), .rdlo_out(a4_wr[1681]));
			radix2 #(.width(width)) rd_st3_1554  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1554]), .rdlo_in(a3_wr[1682]),  .coef_in(coef[144]), .rdup_out(a4_wr[1554]), .rdlo_out(a4_wr[1682]));
			radix2 #(.width(width)) rd_st3_1555  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1555]), .rdlo_in(a3_wr[1683]),  .coef_in(coef[152]), .rdup_out(a4_wr[1555]), .rdlo_out(a4_wr[1683]));
			radix2 #(.width(width)) rd_st3_1556  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1556]), .rdlo_in(a3_wr[1684]),  .coef_in(coef[160]), .rdup_out(a4_wr[1556]), .rdlo_out(a4_wr[1684]));
			radix2 #(.width(width)) rd_st3_1557  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1557]), .rdlo_in(a3_wr[1685]),  .coef_in(coef[168]), .rdup_out(a4_wr[1557]), .rdlo_out(a4_wr[1685]));
			radix2 #(.width(width)) rd_st3_1558  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1558]), .rdlo_in(a3_wr[1686]),  .coef_in(coef[176]), .rdup_out(a4_wr[1558]), .rdlo_out(a4_wr[1686]));
			radix2 #(.width(width)) rd_st3_1559  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1559]), .rdlo_in(a3_wr[1687]),  .coef_in(coef[184]), .rdup_out(a4_wr[1559]), .rdlo_out(a4_wr[1687]));
			radix2 #(.width(width)) rd_st3_1560  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1560]), .rdlo_in(a3_wr[1688]),  .coef_in(coef[192]), .rdup_out(a4_wr[1560]), .rdlo_out(a4_wr[1688]));
			radix2 #(.width(width)) rd_st3_1561  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1561]), .rdlo_in(a3_wr[1689]),  .coef_in(coef[200]), .rdup_out(a4_wr[1561]), .rdlo_out(a4_wr[1689]));
			radix2 #(.width(width)) rd_st3_1562  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1562]), .rdlo_in(a3_wr[1690]),  .coef_in(coef[208]), .rdup_out(a4_wr[1562]), .rdlo_out(a4_wr[1690]));
			radix2 #(.width(width)) rd_st3_1563  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1563]), .rdlo_in(a3_wr[1691]),  .coef_in(coef[216]), .rdup_out(a4_wr[1563]), .rdlo_out(a4_wr[1691]));
			radix2 #(.width(width)) rd_st3_1564  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1564]), .rdlo_in(a3_wr[1692]),  .coef_in(coef[224]), .rdup_out(a4_wr[1564]), .rdlo_out(a4_wr[1692]));
			radix2 #(.width(width)) rd_st3_1565  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1565]), .rdlo_in(a3_wr[1693]),  .coef_in(coef[232]), .rdup_out(a4_wr[1565]), .rdlo_out(a4_wr[1693]));
			radix2 #(.width(width)) rd_st3_1566  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1566]), .rdlo_in(a3_wr[1694]),  .coef_in(coef[240]), .rdup_out(a4_wr[1566]), .rdlo_out(a4_wr[1694]));
			radix2 #(.width(width)) rd_st3_1567  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1567]), .rdlo_in(a3_wr[1695]),  .coef_in(coef[248]), .rdup_out(a4_wr[1567]), .rdlo_out(a4_wr[1695]));
			radix2 #(.width(width)) rd_st3_1568  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1568]), .rdlo_in(a3_wr[1696]),  .coef_in(coef[256]), .rdup_out(a4_wr[1568]), .rdlo_out(a4_wr[1696]));
			radix2 #(.width(width)) rd_st3_1569  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1569]), .rdlo_in(a3_wr[1697]),  .coef_in(coef[264]), .rdup_out(a4_wr[1569]), .rdlo_out(a4_wr[1697]));
			radix2 #(.width(width)) rd_st3_1570  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1570]), .rdlo_in(a3_wr[1698]),  .coef_in(coef[272]), .rdup_out(a4_wr[1570]), .rdlo_out(a4_wr[1698]));
			radix2 #(.width(width)) rd_st3_1571  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1571]), .rdlo_in(a3_wr[1699]),  .coef_in(coef[280]), .rdup_out(a4_wr[1571]), .rdlo_out(a4_wr[1699]));
			radix2 #(.width(width)) rd_st3_1572  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1572]), .rdlo_in(a3_wr[1700]),  .coef_in(coef[288]), .rdup_out(a4_wr[1572]), .rdlo_out(a4_wr[1700]));
			radix2 #(.width(width)) rd_st3_1573  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1573]), .rdlo_in(a3_wr[1701]),  .coef_in(coef[296]), .rdup_out(a4_wr[1573]), .rdlo_out(a4_wr[1701]));
			radix2 #(.width(width)) rd_st3_1574  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1574]), .rdlo_in(a3_wr[1702]),  .coef_in(coef[304]), .rdup_out(a4_wr[1574]), .rdlo_out(a4_wr[1702]));
			radix2 #(.width(width)) rd_st3_1575  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1575]), .rdlo_in(a3_wr[1703]),  .coef_in(coef[312]), .rdup_out(a4_wr[1575]), .rdlo_out(a4_wr[1703]));
			radix2 #(.width(width)) rd_st3_1576  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1576]), .rdlo_in(a3_wr[1704]),  .coef_in(coef[320]), .rdup_out(a4_wr[1576]), .rdlo_out(a4_wr[1704]));
			radix2 #(.width(width)) rd_st3_1577  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1577]), .rdlo_in(a3_wr[1705]),  .coef_in(coef[328]), .rdup_out(a4_wr[1577]), .rdlo_out(a4_wr[1705]));
			radix2 #(.width(width)) rd_st3_1578  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1578]), .rdlo_in(a3_wr[1706]),  .coef_in(coef[336]), .rdup_out(a4_wr[1578]), .rdlo_out(a4_wr[1706]));
			radix2 #(.width(width)) rd_st3_1579  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1579]), .rdlo_in(a3_wr[1707]),  .coef_in(coef[344]), .rdup_out(a4_wr[1579]), .rdlo_out(a4_wr[1707]));
			radix2 #(.width(width)) rd_st3_1580  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1580]), .rdlo_in(a3_wr[1708]),  .coef_in(coef[352]), .rdup_out(a4_wr[1580]), .rdlo_out(a4_wr[1708]));
			radix2 #(.width(width)) rd_st3_1581  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1581]), .rdlo_in(a3_wr[1709]),  .coef_in(coef[360]), .rdup_out(a4_wr[1581]), .rdlo_out(a4_wr[1709]));
			radix2 #(.width(width)) rd_st3_1582  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1582]), .rdlo_in(a3_wr[1710]),  .coef_in(coef[368]), .rdup_out(a4_wr[1582]), .rdlo_out(a4_wr[1710]));
			radix2 #(.width(width)) rd_st3_1583  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1583]), .rdlo_in(a3_wr[1711]),  .coef_in(coef[376]), .rdup_out(a4_wr[1583]), .rdlo_out(a4_wr[1711]));
			radix2 #(.width(width)) rd_st3_1584  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1584]), .rdlo_in(a3_wr[1712]),  .coef_in(coef[384]), .rdup_out(a4_wr[1584]), .rdlo_out(a4_wr[1712]));
			radix2 #(.width(width)) rd_st3_1585  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1585]), .rdlo_in(a3_wr[1713]),  .coef_in(coef[392]), .rdup_out(a4_wr[1585]), .rdlo_out(a4_wr[1713]));
			radix2 #(.width(width)) rd_st3_1586  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1586]), .rdlo_in(a3_wr[1714]),  .coef_in(coef[400]), .rdup_out(a4_wr[1586]), .rdlo_out(a4_wr[1714]));
			radix2 #(.width(width)) rd_st3_1587  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1587]), .rdlo_in(a3_wr[1715]),  .coef_in(coef[408]), .rdup_out(a4_wr[1587]), .rdlo_out(a4_wr[1715]));
			radix2 #(.width(width)) rd_st3_1588  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1588]), .rdlo_in(a3_wr[1716]),  .coef_in(coef[416]), .rdup_out(a4_wr[1588]), .rdlo_out(a4_wr[1716]));
			radix2 #(.width(width)) rd_st3_1589  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1589]), .rdlo_in(a3_wr[1717]),  .coef_in(coef[424]), .rdup_out(a4_wr[1589]), .rdlo_out(a4_wr[1717]));
			radix2 #(.width(width)) rd_st3_1590  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1590]), .rdlo_in(a3_wr[1718]),  .coef_in(coef[432]), .rdup_out(a4_wr[1590]), .rdlo_out(a4_wr[1718]));
			radix2 #(.width(width)) rd_st3_1591  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1591]), .rdlo_in(a3_wr[1719]),  .coef_in(coef[440]), .rdup_out(a4_wr[1591]), .rdlo_out(a4_wr[1719]));
			radix2 #(.width(width)) rd_st3_1592  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1592]), .rdlo_in(a3_wr[1720]),  .coef_in(coef[448]), .rdup_out(a4_wr[1592]), .rdlo_out(a4_wr[1720]));
			radix2 #(.width(width)) rd_st3_1593  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1593]), .rdlo_in(a3_wr[1721]),  .coef_in(coef[456]), .rdup_out(a4_wr[1593]), .rdlo_out(a4_wr[1721]));
			radix2 #(.width(width)) rd_st3_1594  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1594]), .rdlo_in(a3_wr[1722]),  .coef_in(coef[464]), .rdup_out(a4_wr[1594]), .rdlo_out(a4_wr[1722]));
			radix2 #(.width(width)) rd_st3_1595  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1595]), .rdlo_in(a3_wr[1723]),  .coef_in(coef[472]), .rdup_out(a4_wr[1595]), .rdlo_out(a4_wr[1723]));
			radix2 #(.width(width)) rd_st3_1596  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1596]), .rdlo_in(a3_wr[1724]),  .coef_in(coef[480]), .rdup_out(a4_wr[1596]), .rdlo_out(a4_wr[1724]));
			radix2 #(.width(width)) rd_st3_1597  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1597]), .rdlo_in(a3_wr[1725]),  .coef_in(coef[488]), .rdup_out(a4_wr[1597]), .rdlo_out(a4_wr[1725]));
			radix2 #(.width(width)) rd_st3_1598  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1598]), .rdlo_in(a3_wr[1726]),  .coef_in(coef[496]), .rdup_out(a4_wr[1598]), .rdlo_out(a4_wr[1726]));
			radix2 #(.width(width)) rd_st3_1599  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1599]), .rdlo_in(a3_wr[1727]),  .coef_in(coef[504]), .rdup_out(a4_wr[1599]), .rdlo_out(a4_wr[1727]));
			radix2 #(.width(width)) rd_st3_1600  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1600]), .rdlo_in(a3_wr[1728]),  .coef_in(coef[512]), .rdup_out(a4_wr[1600]), .rdlo_out(a4_wr[1728]));
			radix2 #(.width(width)) rd_st3_1601  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1601]), .rdlo_in(a3_wr[1729]),  .coef_in(coef[520]), .rdup_out(a4_wr[1601]), .rdlo_out(a4_wr[1729]));
			radix2 #(.width(width)) rd_st3_1602  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1602]), .rdlo_in(a3_wr[1730]),  .coef_in(coef[528]), .rdup_out(a4_wr[1602]), .rdlo_out(a4_wr[1730]));
			radix2 #(.width(width)) rd_st3_1603  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1603]), .rdlo_in(a3_wr[1731]),  .coef_in(coef[536]), .rdup_out(a4_wr[1603]), .rdlo_out(a4_wr[1731]));
			radix2 #(.width(width)) rd_st3_1604  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1604]), .rdlo_in(a3_wr[1732]),  .coef_in(coef[544]), .rdup_out(a4_wr[1604]), .rdlo_out(a4_wr[1732]));
			radix2 #(.width(width)) rd_st3_1605  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1605]), .rdlo_in(a3_wr[1733]),  .coef_in(coef[552]), .rdup_out(a4_wr[1605]), .rdlo_out(a4_wr[1733]));
			radix2 #(.width(width)) rd_st3_1606  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1606]), .rdlo_in(a3_wr[1734]),  .coef_in(coef[560]), .rdup_out(a4_wr[1606]), .rdlo_out(a4_wr[1734]));
			radix2 #(.width(width)) rd_st3_1607  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1607]), .rdlo_in(a3_wr[1735]),  .coef_in(coef[568]), .rdup_out(a4_wr[1607]), .rdlo_out(a4_wr[1735]));
			radix2 #(.width(width)) rd_st3_1608  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1608]), .rdlo_in(a3_wr[1736]),  .coef_in(coef[576]), .rdup_out(a4_wr[1608]), .rdlo_out(a4_wr[1736]));
			radix2 #(.width(width)) rd_st3_1609  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1609]), .rdlo_in(a3_wr[1737]),  .coef_in(coef[584]), .rdup_out(a4_wr[1609]), .rdlo_out(a4_wr[1737]));
			radix2 #(.width(width)) rd_st3_1610  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1610]), .rdlo_in(a3_wr[1738]),  .coef_in(coef[592]), .rdup_out(a4_wr[1610]), .rdlo_out(a4_wr[1738]));
			radix2 #(.width(width)) rd_st3_1611  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1611]), .rdlo_in(a3_wr[1739]),  .coef_in(coef[600]), .rdup_out(a4_wr[1611]), .rdlo_out(a4_wr[1739]));
			radix2 #(.width(width)) rd_st3_1612  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1612]), .rdlo_in(a3_wr[1740]),  .coef_in(coef[608]), .rdup_out(a4_wr[1612]), .rdlo_out(a4_wr[1740]));
			radix2 #(.width(width)) rd_st3_1613  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1613]), .rdlo_in(a3_wr[1741]),  .coef_in(coef[616]), .rdup_out(a4_wr[1613]), .rdlo_out(a4_wr[1741]));
			radix2 #(.width(width)) rd_st3_1614  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1614]), .rdlo_in(a3_wr[1742]),  .coef_in(coef[624]), .rdup_out(a4_wr[1614]), .rdlo_out(a4_wr[1742]));
			radix2 #(.width(width)) rd_st3_1615  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1615]), .rdlo_in(a3_wr[1743]),  .coef_in(coef[632]), .rdup_out(a4_wr[1615]), .rdlo_out(a4_wr[1743]));
			radix2 #(.width(width)) rd_st3_1616  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1616]), .rdlo_in(a3_wr[1744]),  .coef_in(coef[640]), .rdup_out(a4_wr[1616]), .rdlo_out(a4_wr[1744]));
			radix2 #(.width(width)) rd_st3_1617  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1617]), .rdlo_in(a3_wr[1745]),  .coef_in(coef[648]), .rdup_out(a4_wr[1617]), .rdlo_out(a4_wr[1745]));
			radix2 #(.width(width)) rd_st3_1618  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1618]), .rdlo_in(a3_wr[1746]),  .coef_in(coef[656]), .rdup_out(a4_wr[1618]), .rdlo_out(a4_wr[1746]));
			radix2 #(.width(width)) rd_st3_1619  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1619]), .rdlo_in(a3_wr[1747]),  .coef_in(coef[664]), .rdup_out(a4_wr[1619]), .rdlo_out(a4_wr[1747]));
			radix2 #(.width(width)) rd_st3_1620  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1620]), .rdlo_in(a3_wr[1748]),  .coef_in(coef[672]), .rdup_out(a4_wr[1620]), .rdlo_out(a4_wr[1748]));
			radix2 #(.width(width)) rd_st3_1621  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1621]), .rdlo_in(a3_wr[1749]),  .coef_in(coef[680]), .rdup_out(a4_wr[1621]), .rdlo_out(a4_wr[1749]));
			radix2 #(.width(width)) rd_st3_1622  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1622]), .rdlo_in(a3_wr[1750]),  .coef_in(coef[688]), .rdup_out(a4_wr[1622]), .rdlo_out(a4_wr[1750]));
			radix2 #(.width(width)) rd_st3_1623  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1623]), .rdlo_in(a3_wr[1751]),  .coef_in(coef[696]), .rdup_out(a4_wr[1623]), .rdlo_out(a4_wr[1751]));
			radix2 #(.width(width)) rd_st3_1624  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1624]), .rdlo_in(a3_wr[1752]),  .coef_in(coef[704]), .rdup_out(a4_wr[1624]), .rdlo_out(a4_wr[1752]));
			radix2 #(.width(width)) rd_st3_1625  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1625]), .rdlo_in(a3_wr[1753]),  .coef_in(coef[712]), .rdup_out(a4_wr[1625]), .rdlo_out(a4_wr[1753]));
			radix2 #(.width(width)) rd_st3_1626  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1626]), .rdlo_in(a3_wr[1754]),  .coef_in(coef[720]), .rdup_out(a4_wr[1626]), .rdlo_out(a4_wr[1754]));
			radix2 #(.width(width)) rd_st3_1627  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1627]), .rdlo_in(a3_wr[1755]),  .coef_in(coef[728]), .rdup_out(a4_wr[1627]), .rdlo_out(a4_wr[1755]));
			radix2 #(.width(width)) rd_st3_1628  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1628]), .rdlo_in(a3_wr[1756]),  .coef_in(coef[736]), .rdup_out(a4_wr[1628]), .rdlo_out(a4_wr[1756]));
			radix2 #(.width(width)) rd_st3_1629  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1629]), .rdlo_in(a3_wr[1757]),  .coef_in(coef[744]), .rdup_out(a4_wr[1629]), .rdlo_out(a4_wr[1757]));
			radix2 #(.width(width)) rd_st3_1630  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1630]), .rdlo_in(a3_wr[1758]),  .coef_in(coef[752]), .rdup_out(a4_wr[1630]), .rdlo_out(a4_wr[1758]));
			radix2 #(.width(width)) rd_st3_1631  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1631]), .rdlo_in(a3_wr[1759]),  .coef_in(coef[760]), .rdup_out(a4_wr[1631]), .rdlo_out(a4_wr[1759]));
			radix2 #(.width(width)) rd_st3_1632  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1632]), .rdlo_in(a3_wr[1760]),  .coef_in(coef[768]), .rdup_out(a4_wr[1632]), .rdlo_out(a4_wr[1760]));
			radix2 #(.width(width)) rd_st3_1633  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1633]), .rdlo_in(a3_wr[1761]),  .coef_in(coef[776]), .rdup_out(a4_wr[1633]), .rdlo_out(a4_wr[1761]));
			radix2 #(.width(width)) rd_st3_1634  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1634]), .rdlo_in(a3_wr[1762]),  .coef_in(coef[784]), .rdup_out(a4_wr[1634]), .rdlo_out(a4_wr[1762]));
			radix2 #(.width(width)) rd_st3_1635  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1635]), .rdlo_in(a3_wr[1763]),  .coef_in(coef[792]), .rdup_out(a4_wr[1635]), .rdlo_out(a4_wr[1763]));
			radix2 #(.width(width)) rd_st3_1636  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1636]), .rdlo_in(a3_wr[1764]),  .coef_in(coef[800]), .rdup_out(a4_wr[1636]), .rdlo_out(a4_wr[1764]));
			radix2 #(.width(width)) rd_st3_1637  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1637]), .rdlo_in(a3_wr[1765]),  .coef_in(coef[808]), .rdup_out(a4_wr[1637]), .rdlo_out(a4_wr[1765]));
			radix2 #(.width(width)) rd_st3_1638  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1638]), .rdlo_in(a3_wr[1766]),  .coef_in(coef[816]), .rdup_out(a4_wr[1638]), .rdlo_out(a4_wr[1766]));
			radix2 #(.width(width)) rd_st3_1639  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1639]), .rdlo_in(a3_wr[1767]),  .coef_in(coef[824]), .rdup_out(a4_wr[1639]), .rdlo_out(a4_wr[1767]));
			radix2 #(.width(width)) rd_st3_1640  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1640]), .rdlo_in(a3_wr[1768]),  .coef_in(coef[832]), .rdup_out(a4_wr[1640]), .rdlo_out(a4_wr[1768]));
			radix2 #(.width(width)) rd_st3_1641  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1641]), .rdlo_in(a3_wr[1769]),  .coef_in(coef[840]), .rdup_out(a4_wr[1641]), .rdlo_out(a4_wr[1769]));
			radix2 #(.width(width)) rd_st3_1642  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1642]), .rdlo_in(a3_wr[1770]),  .coef_in(coef[848]), .rdup_out(a4_wr[1642]), .rdlo_out(a4_wr[1770]));
			radix2 #(.width(width)) rd_st3_1643  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1643]), .rdlo_in(a3_wr[1771]),  .coef_in(coef[856]), .rdup_out(a4_wr[1643]), .rdlo_out(a4_wr[1771]));
			radix2 #(.width(width)) rd_st3_1644  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1644]), .rdlo_in(a3_wr[1772]),  .coef_in(coef[864]), .rdup_out(a4_wr[1644]), .rdlo_out(a4_wr[1772]));
			radix2 #(.width(width)) rd_st3_1645  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1645]), .rdlo_in(a3_wr[1773]),  .coef_in(coef[872]), .rdup_out(a4_wr[1645]), .rdlo_out(a4_wr[1773]));
			radix2 #(.width(width)) rd_st3_1646  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1646]), .rdlo_in(a3_wr[1774]),  .coef_in(coef[880]), .rdup_out(a4_wr[1646]), .rdlo_out(a4_wr[1774]));
			radix2 #(.width(width)) rd_st3_1647  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1647]), .rdlo_in(a3_wr[1775]),  .coef_in(coef[888]), .rdup_out(a4_wr[1647]), .rdlo_out(a4_wr[1775]));
			radix2 #(.width(width)) rd_st3_1648  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1648]), .rdlo_in(a3_wr[1776]),  .coef_in(coef[896]), .rdup_out(a4_wr[1648]), .rdlo_out(a4_wr[1776]));
			radix2 #(.width(width)) rd_st3_1649  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1649]), .rdlo_in(a3_wr[1777]),  .coef_in(coef[904]), .rdup_out(a4_wr[1649]), .rdlo_out(a4_wr[1777]));
			radix2 #(.width(width)) rd_st3_1650  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1650]), .rdlo_in(a3_wr[1778]),  .coef_in(coef[912]), .rdup_out(a4_wr[1650]), .rdlo_out(a4_wr[1778]));
			radix2 #(.width(width)) rd_st3_1651  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1651]), .rdlo_in(a3_wr[1779]),  .coef_in(coef[920]), .rdup_out(a4_wr[1651]), .rdlo_out(a4_wr[1779]));
			radix2 #(.width(width)) rd_st3_1652  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1652]), .rdlo_in(a3_wr[1780]),  .coef_in(coef[928]), .rdup_out(a4_wr[1652]), .rdlo_out(a4_wr[1780]));
			radix2 #(.width(width)) rd_st3_1653  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1653]), .rdlo_in(a3_wr[1781]),  .coef_in(coef[936]), .rdup_out(a4_wr[1653]), .rdlo_out(a4_wr[1781]));
			radix2 #(.width(width)) rd_st3_1654  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1654]), .rdlo_in(a3_wr[1782]),  .coef_in(coef[944]), .rdup_out(a4_wr[1654]), .rdlo_out(a4_wr[1782]));
			radix2 #(.width(width)) rd_st3_1655  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1655]), .rdlo_in(a3_wr[1783]),  .coef_in(coef[952]), .rdup_out(a4_wr[1655]), .rdlo_out(a4_wr[1783]));
			radix2 #(.width(width)) rd_st3_1656  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1656]), .rdlo_in(a3_wr[1784]),  .coef_in(coef[960]), .rdup_out(a4_wr[1656]), .rdlo_out(a4_wr[1784]));
			radix2 #(.width(width)) rd_st3_1657  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1657]), .rdlo_in(a3_wr[1785]),  .coef_in(coef[968]), .rdup_out(a4_wr[1657]), .rdlo_out(a4_wr[1785]));
			radix2 #(.width(width)) rd_st3_1658  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1658]), .rdlo_in(a3_wr[1786]),  .coef_in(coef[976]), .rdup_out(a4_wr[1658]), .rdlo_out(a4_wr[1786]));
			radix2 #(.width(width)) rd_st3_1659  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1659]), .rdlo_in(a3_wr[1787]),  .coef_in(coef[984]), .rdup_out(a4_wr[1659]), .rdlo_out(a4_wr[1787]));
			radix2 #(.width(width)) rd_st3_1660  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1660]), .rdlo_in(a3_wr[1788]),  .coef_in(coef[992]), .rdup_out(a4_wr[1660]), .rdlo_out(a4_wr[1788]));
			radix2 #(.width(width)) rd_st3_1661  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1661]), .rdlo_in(a3_wr[1789]),  .coef_in(coef[1000]), .rdup_out(a4_wr[1661]), .rdlo_out(a4_wr[1789]));
			radix2 #(.width(width)) rd_st3_1662  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1662]), .rdlo_in(a3_wr[1790]),  .coef_in(coef[1008]), .rdup_out(a4_wr[1662]), .rdlo_out(a4_wr[1790]));
			radix2 #(.width(width)) rd_st3_1663  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1663]), .rdlo_in(a3_wr[1791]),  .coef_in(coef[1016]), .rdup_out(a4_wr[1663]), .rdlo_out(a4_wr[1791]));
			radix2 #(.width(width)) rd_st3_1792  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1792]), .rdlo_in(a3_wr[1920]),  .coef_in(coef[0]), .rdup_out(a4_wr[1792]), .rdlo_out(a4_wr[1920]));
			radix2 #(.width(width)) rd_st3_1793  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1793]), .rdlo_in(a3_wr[1921]),  .coef_in(coef[8]), .rdup_out(a4_wr[1793]), .rdlo_out(a4_wr[1921]));
			radix2 #(.width(width)) rd_st3_1794  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1794]), .rdlo_in(a3_wr[1922]),  .coef_in(coef[16]), .rdup_out(a4_wr[1794]), .rdlo_out(a4_wr[1922]));
			radix2 #(.width(width)) rd_st3_1795  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1795]), .rdlo_in(a3_wr[1923]),  .coef_in(coef[24]), .rdup_out(a4_wr[1795]), .rdlo_out(a4_wr[1923]));
			radix2 #(.width(width)) rd_st3_1796  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1796]), .rdlo_in(a3_wr[1924]),  .coef_in(coef[32]), .rdup_out(a4_wr[1796]), .rdlo_out(a4_wr[1924]));
			radix2 #(.width(width)) rd_st3_1797  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1797]), .rdlo_in(a3_wr[1925]),  .coef_in(coef[40]), .rdup_out(a4_wr[1797]), .rdlo_out(a4_wr[1925]));
			radix2 #(.width(width)) rd_st3_1798  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1798]), .rdlo_in(a3_wr[1926]),  .coef_in(coef[48]), .rdup_out(a4_wr[1798]), .rdlo_out(a4_wr[1926]));
			radix2 #(.width(width)) rd_st3_1799  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1799]), .rdlo_in(a3_wr[1927]),  .coef_in(coef[56]), .rdup_out(a4_wr[1799]), .rdlo_out(a4_wr[1927]));
			radix2 #(.width(width)) rd_st3_1800  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1800]), .rdlo_in(a3_wr[1928]),  .coef_in(coef[64]), .rdup_out(a4_wr[1800]), .rdlo_out(a4_wr[1928]));
			radix2 #(.width(width)) rd_st3_1801  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1801]), .rdlo_in(a3_wr[1929]),  .coef_in(coef[72]), .rdup_out(a4_wr[1801]), .rdlo_out(a4_wr[1929]));
			radix2 #(.width(width)) rd_st3_1802  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1802]), .rdlo_in(a3_wr[1930]),  .coef_in(coef[80]), .rdup_out(a4_wr[1802]), .rdlo_out(a4_wr[1930]));
			radix2 #(.width(width)) rd_st3_1803  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1803]), .rdlo_in(a3_wr[1931]),  .coef_in(coef[88]), .rdup_out(a4_wr[1803]), .rdlo_out(a4_wr[1931]));
			radix2 #(.width(width)) rd_st3_1804  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1804]), .rdlo_in(a3_wr[1932]),  .coef_in(coef[96]), .rdup_out(a4_wr[1804]), .rdlo_out(a4_wr[1932]));
			radix2 #(.width(width)) rd_st3_1805  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1805]), .rdlo_in(a3_wr[1933]),  .coef_in(coef[104]), .rdup_out(a4_wr[1805]), .rdlo_out(a4_wr[1933]));
			radix2 #(.width(width)) rd_st3_1806  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1806]), .rdlo_in(a3_wr[1934]),  .coef_in(coef[112]), .rdup_out(a4_wr[1806]), .rdlo_out(a4_wr[1934]));
			radix2 #(.width(width)) rd_st3_1807  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1807]), .rdlo_in(a3_wr[1935]),  .coef_in(coef[120]), .rdup_out(a4_wr[1807]), .rdlo_out(a4_wr[1935]));
			radix2 #(.width(width)) rd_st3_1808  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1808]), .rdlo_in(a3_wr[1936]),  .coef_in(coef[128]), .rdup_out(a4_wr[1808]), .rdlo_out(a4_wr[1936]));
			radix2 #(.width(width)) rd_st3_1809  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1809]), .rdlo_in(a3_wr[1937]),  .coef_in(coef[136]), .rdup_out(a4_wr[1809]), .rdlo_out(a4_wr[1937]));
			radix2 #(.width(width)) rd_st3_1810  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1810]), .rdlo_in(a3_wr[1938]),  .coef_in(coef[144]), .rdup_out(a4_wr[1810]), .rdlo_out(a4_wr[1938]));
			radix2 #(.width(width)) rd_st3_1811  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1811]), .rdlo_in(a3_wr[1939]),  .coef_in(coef[152]), .rdup_out(a4_wr[1811]), .rdlo_out(a4_wr[1939]));
			radix2 #(.width(width)) rd_st3_1812  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1812]), .rdlo_in(a3_wr[1940]),  .coef_in(coef[160]), .rdup_out(a4_wr[1812]), .rdlo_out(a4_wr[1940]));
			radix2 #(.width(width)) rd_st3_1813  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1813]), .rdlo_in(a3_wr[1941]),  .coef_in(coef[168]), .rdup_out(a4_wr[1813]), .rdlo_out(a4_wr[1941]));
			radix2 #(.width(width)) rd_st3_1814  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1814]), .rdlo_in(a3_wr[1942]),  .coef_in(coef[176]), .rdup_out(a4_wr[1814]), .rdlo_out(a4_wr[1942]));
			radix2 #(.width(width)) rd_st3_1815  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1815]), .rdlo_in(a3_wr[1943]),  .coef_in(coef[184]), .rdup_out(a4_wr[1815]), .rdlo_out(a4_wr[1943]));
			radix2 #(.width(width)) rd_st3_1816  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1816]), .rdlo_in(a3_wr[1944]),  .coef_in(coef[192]), .rdup_out(a4_wr[1816]), .rdlo_out(a4_wr[1944]));
			radix2 #(.width(width)) rd_st3_1817  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1817]), .rdlo_in(a3_wr[1945]),  .coef_in(coef[200]), .rdup_out(a4_wr[1817]), .rdlo_out(a4_wr[1945]));
			radix2 #(.width(width)) rd_st3_1818  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1818]), .rdlo_in(a3_wr[1946]),  .coef_in(coef[208]), .rdup_out(a4_wr[1818]), .rdlo_out(a4_wr[1946]));
			radix2 #(.width(width)) rd_st3_1819  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1819]), .rdlo_in(a3_wr[1947]),  .coef_in(coef[216]), .rdup_out(a4_wr[1819]), .rdlo_out(a4_wr[1947]));
			radix2 #(.width(width)) rd_st3_1820  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1820]), .rdlo_in(a3_wr[1948]),  .coef_in(coef[224]), .rdup_out(a4_wr[1820]), .rdlo_out(a4_wr[1948]));
			radix2 #(.width(width)) rd_st3_1821  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1821]), .rdlo_in(a3_wr[1949]),  .coef_in(coef[232]), .rdup_out(a4_wr[1821]), .rdlo_out(a4_wr[1949]));
			radix2 #(.width(width)) rd_st3_1822  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1822]), .rdlo_in(a3_wr[1950]),  .coef_in(coef[240]), .rdup_out(a4_wr[1822]), .rdlo_out(a4_wr[1950]));
			radix2 #(.width(width)) rd_st3_1823  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1823]), .rdlo_in(a3_wr[1951]),  .coef_in(coef[248]), .rdup_out(a4_wr[1823]), .rdlo_out(a4_wr[1951]));
			radix2 #(.width(width)) rd_st3_1824  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1824]), .rdlo_in(a3_wr[1952]),  .coef_in(coef[256]), .rdup_out(a4_wr[1824]), .rdlo_out(a4_wr[1952]));
			radix2 #(.width(width)) rd_st3_1825  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1825]), .rdlo_in(a3_wr[1953]),  .coef_in(coef[264]), .rdup_out(a4_wr[1825]), .rdlo_out(a4_wr[1953]));
			radix2 #(.width(width)) rd_st3_1826  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1826]), .rdlo_in(a3_wr[1954]),  .coef_in(coef[272]), .rdup_out(a4_wr[1826]), .rdlo_out(a4_wr[1954]));
			radix2 #(.width(width)) rd_st3_1827  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1827]), .rdlo_in(a3_wr[1955]),  .coef_in(coef[280]), .rdup_out(a4_wr[1827]), .rdlo_out(a4_wr[1955]));
			radix2 #(.width(width)) rd_st3_1828  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1828]), .rdlo_in(a3_wr[1956]),  .coef_in(coef[288]), .rdup_out(a4_wr[1828]), .rdlo_out(a4_wr[1956]));
			radix2 #(.width(width)) rd_st3_1829  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1829]), .rdlo_in(a3_wr[1957]),  .coef_in(coef[296]), .rdup_out(a4_wr[1829]), .rdlo_out(a4_wr[1957]));
			radix2 #(.width(width)) rd_st3_1830  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1830]), .rdlo_in(a3_wr[1958]),  .coef_in(coef[304]), .rdup_out(a4_wr[1830]), .rdlo_out(a4_wr[1958]));
			radix2 #(.width(width)) rd_st3_1831  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1831]), .rdlo_in(a3_wr[1959]),  .coef_in(coef[312]), .rdup_out(a4_wr[1831]), .rdlo_out(a4_wr[1959]));
			radix2 #(.width(width)) rd_st3_1832  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1832]), .rdlo_in(a3_wr[1960]),  .coef_in(coef[320]), .rdup_out(a4_wr[1832]), .rdlo_out(a4_wr[1960]));
			radix2 #(.width(width)) rd_st3_1833  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1833]), .rdlo_in(a3_wr[1961]),  .coef_in(coef[328]), .rdup_out(a4_wr[1833]), .rdlo_out(a4_wr[1961]));
			radix2 #(.width(width)) rd_st3_1834  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1834]), .rdlo_in(a3_wr[1962]),  .coef_in(coef[336]), .rdup_out(a4_wr[1834]), .rdlo_out(a4_wr[1962]));
			radix2 #(.width(width)) rd_st3_1835  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1835]), .rdlo_in(a3_wr[1963]),  .coef_in(coef[344]), .rdup_out(a4_wr[1835]), .rdlo_out(a4_wr[1963]));
			radix2 #(.width(width)) rd_st3_1836  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1836]), .rdlo_in(a3_wr[1964]),  .coef_in(coef[352]), .rdup_out(a4_wr[1836]), .rdlo_out(a4_wr[1964]));
			radix2 #(.width(width)) rd_st3_1837  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1837]), .rdlo_in(a3_wr[1965]),  .coef_in(coef[360]), .rdup_out(a4_wr[1837]), .rdlo_out(a4_wr[1965]));
			radix2 #(.width(width)) rd_st3_1838  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1838]), .rdlo_in(a3_wr[1966]),  .coef_in(coef[368]), .rdup_out(a4_wr[1838]), .rdlo_out(a4_wr[1966]));
			radix2 #(.width(width)) rd_st3_1839  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1839]), .rdlo_in(a3_wr[1967]),  .coef_in(coef[376]), .rdup_out(a4_wr[1839]), .rdlo_out(a4_wr[1967]));
			radix2 #(.width(width)) rd_st3_1840  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1840]), .rdlo_in(a3_wr[1968]),  .coef_in(coef[384]), .rdup_out(a4_wr[1840]), .rdlo_out(a4_wr[1968]));
			radix2 #(.width(width)) rd_st3_1841  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1841]), .rdlo_in(a3_wr[1969]),  .coef_in(coef[392]), .rdup_out(a4_wr[1841]), .rdlo_out(a4_wr[1969]));
			radix2 #(.width(width)) rd_st3_1842  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1842]), .rdlo_in(a3_wr[1970]),  .coef_in(coef[400]), .rdup_out(a4_wr[1842]), .rdlo_out(a4_wr[1970]));
			radix2 #(.width(width)) rd_st3_1843  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1843]), .rdlo_in(a3_wr[1971]),  .coef_in(coef[408]), .rdup_out(a4_wr[1843]), .rdlo_out(a4_wr[1971]));
			radix2 #(.width(width)) rd_st3_1844  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1844]), .rdlo_in(a3_wr[1972]),  .coef_in(coef[416]), .rdup_out(a4_wr[1844]), .rdlo_out(a4_wr[1972]));
			radix2 #(.width(width)) rd_st3_1845  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1845]), .rdlo_in(a3_wr[1973]),  .coef_in(coef[424]), .rdup_out(a4_wr[1845]), .rdlo_out(a4_wr[1973]));
			radix2 #(.width(width)) rd_st3_1846  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1846]), .rdlo_in(a3_wr[1974]),  .coef_in(coef[432]), .rdup_out(a4_wr[1846]), .rdlo_out(a4_wr[1974]));
			radix2 #(.width(width)) rd_st3_1847  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1847]), .rdlo_in(a3_wr[1975]),  .coef_in(coef[440]), .rdup_out(a4_wr[1847]), .rdlo_out(a4_wr[1975]));
			radix2 #(.width(width)) rd_st3_1848  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1848]), .rdlo_in(a3_wr[1976]),  .coef_in(coef[448]), .rdup_out(a4_wr[1848]), .rdlo_out(a4_wr[1976]));
			radix2 #(.width(width)) rd_st3_1849  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1849]), .rdlo_in(a3_wr[1977]),  .coef_in(coef[456]), .rdup_out(a4_wr[1849]), .rdlo_out(a4_wr[1977]));
			radix2 #(.width(width)) rd_st3_1850  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1850]), .rdlo_in(a3_wr[1978]),  .coef_in(coef[464]), .rdup_out(a4_wr[1850]), .rdlo_out(a4_wr[1978]));
			radix2 #(.width(width)) rd_st3_1851  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1851]), .rdlo_in(a3_wr[1979]),  .coef_in(coef[472]), .rdup_out(a4_wr[1851]), .rdlo_out(a4_wr[1979]));
			radix2 #(.width(width)) rd_st3_1852  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1852]), .rdlo_in(a3_wr[1980]),  .coef_in(coef[480]), .rdup_out(a4_wr[1852]), .rdlo_out(a4_wr[1980]));
			radix2 #(.width(width)) rd_st3_1853  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1853]), .rdlo_in(a3_wr[1981]),  .coef_in(coef[488]), .rdup_out(a4_wr[1853]), .rdlo_out(a4_wr[1981]));
			radix2 #(.width(width)) rd_st3_1854  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1854]), .rdlo_in(a3_wr[1982]),  .coef_in(coef[496]), .rdup_out(a4_wr[1854]), .rdlo_out(a4_wr[1982]));
			radix2 #(.width(width)) rd_st3_1855  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1855]), .rdlo_in(a3_wr[1983]),  .coef_in(coef[504]), .rdup_out(a4_wr[1855]), .rdlo_out(a4_wr[1983]));
			radix2 #(.width(width)) rd_st3_1856  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1856]), .rdlo_in(a3_wr[1984]),  .coef_in(coef[512]), .rdup_out(a4_wr[1856]), .rdlo_out(a4_wr[1984]));
			radix2 #(.width(width)) rd_st3_1857  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1857]), .rdlo_in(a3_wr[1985]),  .coef_in(coef[520]), .rdup_out(a4_wr[1857]), .rdlo_out(a4_wr[1985]));
			radix2 #(.width(width)) rd_st3_1858  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1858]), .rdlo_in(a3_wr[1986]),  .coef_in(coef[528]), .rdup_out(a4_wr[1858]), .rdlo_out(a4_wr[1986]));
			radix2 #(.width(width)) rd_st3_1859  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1859]), .rdlo_in(a3_wr[1987]),  .coef_in(coef[536]), .rdup_out(a4_wr[1859]), .rdlo_out(a4_wr[1987]));
			radix2 #(.width(width)) rd_st3_1860  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1860]), .rdlo_in(a3_wr[1988]),  .coef_in(coef[544]), .rdup_out(a4_wr[1860]), .rdlo_out(a4_wr[1988]));
			radix2 #(.width(width)) rd_st3_1861  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1861]), .rdlo_in(a3_wr[1989]),  .coef_in(coef[552]), .rdup_out(a4_wr[1861]), .rdlo_out(a4_wr[1989]));
			radix2 #(.width(width)) rd_st3_1862  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1862]), .rdlo_in(a3_wr[1990]),  .coef_in(coef[560]), .rdup_out(a4_wr[1862]), .rdlo_out(a4_wr[1990]));
			radix2 #(.width(width)) rd_st3_1863  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1863]), .rdlo_in(a3_wr[1991]),  .coef_in(coef[568]), .rdup_out(a4_wr[1863]), .rdlo_out(a4_wr[1991]));
			radix2 #(.width(width)) rd_st3_1864  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1864]), .rdlo_in(a3_wr[1992]),  .coef_in(coef[576]), .rdup_out(a4_wr[1864]), .rdlo_out(a4_wr[1992]));
			radix2 #(.width(width)) rd_st3_1865  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1865]), .rdlo_in(a3_wr[1993]),  .coef_in(coef[584]), .rdup_out(a4_wr[1865]), .rdlo_out(a4_wr[1993]));
			radix2 #(.width(width)) rd_st3_1866  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1866]), .rdlo_in(a3_wr[1994]),  .coef_in(coef[592]), .rdup_out(a4_wr[1866]), .rdlo_out(a4_wr[1994]));
			radix2 #(.width(width)) rd_st3_1867  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1867]), .rdlo_in(a3_wr[1995]),  .coef_in(coef[600]), .rdup_out(a4_wr[1867]), .rdlo_out(a4_wr[1995]));
			radix2 #(.width(width)) rd_st3_1868  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1868]), .rdlo_in(a3_wr[1996]),  .coef_in(coef[608]), .rdup_out(a4_wr[1868]), .rdlo_out(a4_wr[1996]));
			radix2 #(.width(width)) rd_st3_1869  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1869]), .rdlo_in(a3_wr[1997]),  .coef_in(coef[616]), .rdup_out(a4_wr[1869]), .rdlo_out(a4_wr[1997]));
			radix2 #(.width(width)) rd_st3_1870  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1870]), .rdlo_in(a3_wr[1998]),  .coef_in(coef[624]), .rdup_out(a4_wr[1870]), .rdlo_out(a4_wr[1998]));
			radix2 #(.width(width)) rd_st3_1871  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1871]), .rdlo_in(a3_wr[1999]),  .coef_in(coef[632]), .rdup_out(a4_wr[1871]), .rdlo_out(a4_wr[1999]));
			radix2 #(.width(width)) rd_st3_1872  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1872]), .rdlo_in(a3_wr[2000]),  .coef_in(coef[640]), .rdup_out(a4_wr[1872]), .rdlo_out(a4_wr[2000]));
			radix2 #(.width(width)) rd_st3_1873  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1873]), .rdlo_in(a3_wr[2001]),  .coef_in(coef[648]), .rdup_out(a4_wr[1873]), .rdlo_out(a4_wr[2001]));
			radix2 #(.width(width)) rd_st3_1874  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1874]), .rdlo_in(a3_wr[2002]),  .coef_in(coef[656]), .rdup_out(a4_wr[1874]), .rdlo_out(a4_wr[2002]));
			radix2 #(.width(width)) rd_st3_1875  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1875]), .rdlo_in(a3_wr[2003]),  .coef_in(coef[664]), .rdup_out(a4_wr[1875]), .rdlo_out(a4_wr[2003]));
			radix2 #(.width(width)) rd_st3_1876  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1876]), .rdlo_in(a3_wr[2004]),  .coef_in(coef[672]), .rdup_out(a4_wr[1876]), .rdlo_out(a4_wr[2004]));
			radix2 #(.width(width)) rd_st3_1877  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1877]), .rdlo_in(a3_wr[2005]),  .coef_in(coef[680]), .rdup_out(a4_wr[1877]), .rdlo_out(a4_wr[2005]));
			radix2 #(.width(width)) rd_st3_1878  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1878]), .rdlo_in(a3_wr[2006]),  .coef_in(coef[688]), .rdup_out(a4_wr[1878]), .rdlo_out(a4_wr[2006]));
			radix2 #(.width(width)) rd_st3_1879  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1879]), .rdlo_in(a3_wr[2007]),  .coef_in(coef[696]), .rdup_out(a4_wr[1879]), .rdlo_out(a4_wr[2007]));
			radix2 #(.width(width)) rd_st3_1880  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1880]), .rdlo_in(a3_wr[2008]),  .coef_in(coef[704]), .rdup_out(a4_wr[1880]), .rdlo_out(a4_wr[2008]));
			radix2 #(.width(width)) rd_st3_1881  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1881]), .rdlo_in(a3_wr[2009]),  .coef_in(coef[712]), .rdup_out(a4_wr[1881]), .rdlo_out(a4_wr[2009]));
			radix2 #(.width(width)) rd_st3_1882  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1882]), .rdlo_in(a3_wr[2010]),  .coef_in(coef[720]), .rdup_out(a4_wr[1882]), .rdlo_out(a4_wr[2010]));
			radix2 #(.width(width)) rd_st3_1883  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1883]), .rdlo_in(a3_wr[2011]),  .coef_in(coef[728]), .rdup_out(a4_wr[1883]), .rdlo_out(a4_wr[2011]));
			radix2 #(.width(width)) rd_st3_1884  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1884]), .rdlo_in(a3_wr[2012]),  .coef_in(coef[736]), .rdup_out(a4_wr[1884]), .rdlo_out(a4_wr[2012]));
			radix2 #(.width(width)) rd_st3_1885  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1885]), .rdlo_in(a3_wr[2013]),  .coef_in(coef[744]), .rdup_out(a4_wr[1885]), .rdlo_out(a4_wr[2013]));
			radix2 #(.width(width)) rd_st3_1886  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1886]), .rdlo_in(a3_wr[2014]),  .coef_in(coef[752]), .rdup_out(a4_wr[1886]), .rdlo_out(a4_wr[2014]));
			radix2 #(.width(width)) rd_st3_1887  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1887]), .rdlo_in(a3_wr[2015]),  .coef_in(coef[760]), .rdup_out(a4_wr[1887]), .rdlo_out(a4_wr[2015]));
			radix2 #(.width(width)) rd_st3_1888  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1888]), .rdlo_in(a3_wr[2016]),  .coef_in(coef[768]), .rdup_out(a4_wr[1888]), .rdlo_out(a4_wr[2016]));
			radix2 #(.width(width)) rd_st3_1889  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1889]), .rdlo_in(a3_wr[2017]),  .coef_in(coef[776]), .rdup_out(a4_wr[1889]), .rdlo_out(a4_wr[2017]));
			radix2 #(.width(width)) rd_st3_1890  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1890]), .rdlo_in(a3_wr[2018]),  .coef_in(coef[784]), .rdup_out(a4_wr[1890]), .rdlo_out(a4_wr[2018]));
			radix2 #(.width(width)) rd_st3_1891  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1891]), .rdlo_in(a3_wr[2019]),  .coef_in(coef[792]), .rdup_out(a4_wr[1891]), .rdlo_out(a4_wr[2019]));
			radix2 #(.width(width)) rd_st3_1892  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1892]), .rdlo_in(a3_wr[2020]),  .coef_in(coef[800]), .rdup_out(a4_wr[1892]), .rdlo_out(a4_wr[2020]));
			radix2 #(.width(width)) rd_st3_1893  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1893]), .rdlo_in(a3_wr[2021]),  .coef_in(coef[808]), .rdup_out(a4_wr[1893]), .rdlo_out(a4_wr[2021]));
			radix2 #(.width(width)) rd_st3_1894  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1894]), .rdlo_in(a3_wr[2022]),  .coef_in(coef[816]), .rdup_out(a4_wr[1894]), .rdlo_out(a4_wr[2022]));
			radix2 #(.width(width)) rd_st3_1895  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1895]), .rdlo_in(a3_wr[2023]),  .coef_in(coef[824]), .rdup_out(a4_wr[1895]), .rdlo_out(a4_wr[2023]));
			radix2 #(.width(width)) rd_st3_1896  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1896]), .rdlo_in(a3_wr[2024]),  .coef_in(coef[832]), .rdup_out(a4_wr[1896]), .rdlo_out(a4_wr[2024]));
			radix2 #(.width(width)) rd_st3_1897  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1897]), .rdlo_in(a3_wr[2025]),  .coef_in(coef[840]), .rdup_out(a4_wr[1897]), .rdlo_out(a4_wr[2025]));
			radix2 #(.width(width)) rd_st3_1898  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1898]), .rdlo_in(a3_wr[2026]),  .coef_in(coef[848]), .rdup_out(a4_wr[1898]), .rdlo_out(a4_wr[2026]));
			radix2 #(.width(width)) rd_st3_1899  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1899]), .rdlo_in(a3_wr[2027]),  .coef_in(coef[856]), .rdup_out(a4_wr[1899]), .rdlo_out(a4_wr[2027]));
			radix2 #(.width(width)) rd_st3_1900  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1900]), .rdlo_in(a3_wr[2028]),  .coef_in(coef[864]), .rdup_out(a4_wr[1900]), .rdlo_out(a4_wr[2028]));
			radix2 #(.width(width)) rd_st3_1901  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1901]), .rdlo_in(a3_wr[2029]),  .coef_in(coef[872]), .rdup_out(a4_wr[1901]), .rdlo_out(a4_wr[2029]));
			radix2 #(.width(width)) rd_st3_1902  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1902]), .rdlo_in(a3_wr[2030]),  .coef_in(coef[880]), .rdup_out(a4_wr[1902]), .rdlo_out(a4_wr[2030]));
			radix2 #(.width(width)) rd_st3_1903  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1903]), .rdlo_in(a3_wr[2031]),  .coef_in(coef[888]), .rdup_out(a4_wr[1903]), .rdlo_out(a4_wr[2031]));
			radix2 #(.width(width)) rd_st3_1904  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1904]), .rdlo_in(a3_wr[2032]),  .coef_in(coef[896]), .rdup_out(a4_wr[1904]), .rdlo_out(a4_wr[2032]));
			radix2 #(.width(width)) rd_st3_1905  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1905]), .rdlo_in(a3_wr[2033]),  .coef_in(coef[904]), .rdup_out(a4_wr[1905]), .rdlo_out(a4_wr[2033]));
			radix2 #(.width(width)) rd_st3_1906  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1906]), .rdlo_in(a3_wr[2034]),  .coef_in(coef[912]), .rdup_out(a4_wr[1906]), .rdlo_out(a4_wr[2034]));
			radix2 #(.width(width)) rd_st3_1907  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1907]), .rdlo_in(a3_wr[2035]),  .coef_in(coef[920]), .rdup_out(a4_wr[1907]), .rdlo_out(a4_wr[2035]));
			radix2 #(.width(width)) rd_st3_1908  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1908]), .rdlo_in(a3_wr[2036]),  .coef_in(coef[928]), .rdup_out(a4_wr[1908]), .rdlo_out(a4_wr[2036]));
			radix2 #(.width(width)) rd_st3_1909  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1909]), .rdlo_in(a3_wr[2037]),  .coef_in(coef[936]), .rdup_out(a4_wr[1909]), .rdlo_out(a4_wr[2037]));
			radix2 #(.width(width)) rd_st3_1910  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1910]), .rdlo_in(a3_wr[2038]),  .coef_in(coef[944]), .rdup_out(a4_wr[1910]), .rdlo_out(a4_wr[2038]));
			radix2 #(.width(width)) rd_st3_1911  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1911]), .rdlo_in(a3_wr[2039]),  .coef_in(coef[952]), .rdup_out(a4_wr[1911]), .rdlo_out(a4_wr[2039]));
			radix2 #(.width(width)) rd_st3_1912  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1912]), .rdlo_in(a3_wr[2040]),  .coef_in(coef[960]), .rdup_out(a4_wr[1912]), .rdlo_out(a4_wr[2040]));
			radix2 #(.width(width)) rd_st3_1913  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1913]), .rdlo_in(a3_wr[2041]),  .coef_in(coef[968]), .rdup_out(a4_wr[1913]), .rdlo_out(a4_wr[2041]));
			radix2 #(.width(width)) rd_st3_1914  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1914]), .rdlo_in(a3_wr[2042]),  .coef_in(coef[976]), .rdup_out(a4_wr[1914]), .rdlo_out(a4_wr[2042]));
			radix2 #(.width(width)) rd_st3_1915  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1915]), .rdlo_in(a3_wr[2043]),  .coef_in(coef[984]), .rdup_out(a4_wr[1915]), .rdlo_out(a4_wr[2043]));
			radix2 #(.width(width)) rd_st3_1916  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1916]), .rdlo_in(a3_wr[2044]),  .coef_in(coef[992]), .rdup_out(a4_wr[1916]), .rdlo_out(a4_wr[2044]));
			radix2 #(.width(width)) rd_st3_1917  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1917]), .rdlo_in(a3_wr[2045]),  .coef_in(coef[1000]), .rdup_out(a4_wr[1917]), .rdlo_out(a4_wr[2045]));
			radix2 #(.width(width)) rd_st3_1918  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1918]), .rdlo_in(a3_wr[2046]),  .coef_in(coef[1008]), .rdup_out(a4_wr[1918]), .rdlo_out(a4_wr[2046]));
			radix2 #(.width(width)) rd_st3_1919  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a3_wr[1919]), .rdlo_in(a3_wr[2047]),  .coef_in(coef[1016]), .rdup_out(a4_wr[1919]), .rdlo_out(a4_wr[2047]));

		//--- radix stage 4
			radix2 #(.width(width)) rd_st4_0   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[0]), .rdlo_in(a4_wr[64]),  .coef_in(coef[0]), .rdup_out(a5_wr[0]), .rdlo_out(a5_wr[64]));
			radix2 #(.width(width)) rd_st4_1   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1]), .rdlo_in(a4_wr[65]),  .coef_in(coef[16]), .rdup_out(a5_wr[1]), .rdlo_out(a5_wr[65]));
			radix2 #(.width(width)) rd_st4_2   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[2]), .rdlo_in(a4_wr[66]),  .coef_in(coef[32]), .rdup_out(a5_wr[2]), .rdlo_out(a5_wr[66]));
			radix2 #(.width(width)) rd_st4_3   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[3]), .rdlo_in(a4_wr[67]),  .coef_in(coef[48]), .rdup_out(a5_wr[3]), .rdlo_out(a5_wr[67]));
			radix2 #(.width(width)) rd_st4_4   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[4]), .rdlo_in(a4_wr[68]),  .coef_in(coef[64]), .rdup_out(a5_wr[4]), .rdlo_out(a5_wr[68]));
			radix2 #(.width(width)) rd_st4_5   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[5]), .rdlo_in(a4_wr[69]),  .coef_in(coef[80]), .rdup_out(a5_wr[5]), .rdlo_out(a5_wr[69]));
			radix2 #(.width(width)) rd_st4_6   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[6]), .rdlo_in(a4_wr[70]),  .coef_in(coef[96]), .rdup_out(a5_wr[6]), .rdlo_out(a5_wr[70]));
			radix2 #(.width(width)) rd_st4_7   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[7]), .rdlo_in(a4_wr[71]),  .coef_in(coef[112]), .rdup_out(a5_wr[7]), .rdlo_out(a5_wr[71]));
			radix2 #(.width(width)) rd_st4_8   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[8]), .rdlo_in(a4_wr[72]),  .coef_in(coef[128]), .rdup_out(a5_wr[8]), .rdlo_out(a5_wr[72]));
			radix2 #(.width(width)) rd_st4_9   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[9]), .rdlo_in(a4_wr[73]),  .coef_in(coef[144]), .rdup_out(a5_wr[9]), .rdlo_out(a5_wr[73]));
			radix2 #(.width(width)) rd_st4_10  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[10]), .rdlo_in(a4_wr[74]),  .coef_in(coef[160]), .rdup_out(a5_wr[10]), .rdlo_out(a5_wr[74]));
			radix2 #(.width(width)) rd_st4_11  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[11]), .rdlo_in(a4_wr[75]),  .coef_in(coef[176]), .rdup_out(a5_wr[11]), .rdlo_out(a5_wr[75]));
			radix2 #(.width(width)) rd_st4_12  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[12]), .rdlo_in(a4_wr[76]),  .coef_in(coef[192]), .rdup_out(a5_wr[12]), .rdlo_out(a5_wr[76]));
			radix2 #(.width(width)) rd_st4_13  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[13]), .rdlo_in(a4_wr[77]),  .coef_in(coef[208]), .rdup_out(a5_wr[13]), .rdlo_out(a5_wr[77]));
			radix2 #(.width(width)) rd_st4_14  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[14]), .rdlo_in(a4_wr[78]),  .coef_in(coef[224]), .rdup_out(a5_wr[14]), .rdlo_out(a5_wr[78]));
			radix2 #(.width(width)) rd_st4_15  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[15]), .rdlo_in(a4_wr[79]),  .coef_in(coef[240]), .rdup_out(a5_wr[15]), .rdlo_out(a5_wr[79]));
			radix2 #(.width(width)) rd_st4_16  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[16]), .rdlo_in(a4_wr[80]),  .coef_in(coef[256]), .rdup_out(a5_wr[16]), .rdlo_out(a5_wr[80]));
			radix2 #(.width(width)) rd_st4_17  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[17]), .rdlo_in(a4_wr[81]),  .coef_in(coef[272]), .rdup_out(a5_wr[17]), .rdlo_out(a5_wr[81]));
			radix2 #(.width(width)) rd_st4_18  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[18]), .rdlo_in(a4_wr[82]),  .coef_in(coef[288]), .rdup_out(a5_wr[18]), .rdlo_out(a5_wr[82]));
			radix2 #(.width(width)) rd_st4_19  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[19]), .rdlo_in(a4_wr[83]),  .coef_in(coef[304]), .rdup_out(a5_wr[19]), .rdlo_out(a5_wr[83]));
			radix2 #(.width(width)) rd_st4_20  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[20]), .rdlo_in(a4_wr[84]),  .coef_in(coef[320]), .rdup_out(a5_wr[20]), .rdlo_out(a5_wr[84]));
			radix2 #(.width(width)) rd_st4_21  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[21]), .rdlo_in(a4_wr[85]),  .coef_in(coef[336]), .rdup_out(a5_wr[21]), .rdlo_out(a5_wr[85]));
			radix2 #(.width(width)) rd_st4_22  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[22]), .rdlo_in(a4_wr[86]),  .coef_in(coef[352]), .rdup_out(a5_wr[22]), .rdlo_out(a5_wr[86]));
			radix2 #(.width(width)) rd_st4_23  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[23]), .rdlo_in(a4_wr[87]),  .coef_in(coef[368]), .rdup_out(a5_wr[23]), .rdlo_out(a5_wr[87]));
			radix2 #(.width(width)) rd_st4_24  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[24]), .rdlo_in(a4_wr[88]),  .coef_in(coef[384]), .rdup_out(a5_wr[24]), .rdlo_out(a5_wr[88]));
			radix2 #(.width(width)) rd_st4_25  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[25]), .rdlo_in(a4_wr[89]),  .coef_in(coef[400]), .rdup_out(a5_wr[25]), .rdlo_out(a5_wr[89]));
			radix2 #(.width(width)) rd_st4_26  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[26]), .rdlo_in(a4_wr[90]),  .coef_in(coef[416]), .rdup_out(a5_wr[26]), .rdlo_out(a5_wr[90]));
			radix2 #(.width(width)) rd_st4_27  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[27]), .rdlo_in(a4_wr[91]),  .coef_in(coef[432]), .rdup_out(a5_wr[27]), .rdlo_out(a5_wr[91]));
			radix2 #(.width(width)) rd_st4_28  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[28]), .rdlo_in(a4_wr[92]),  .coef_in(coef[448]), .rdup_out(a5_wr[28]), .rdlo_out(a5_wr[92]));
			radix2 #(.width(width)) rd_st4_29  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[29]), .rdlo_in(a4_wr[93]),  .coef_in(coef[464]), .rdup_out(a5_wr[29]), .rdlo_out(a5_wr[93]));
			radix2 #(.width(width)) rd_st4_30  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[30]), .rdlo_in(a4_wr[94]),  .coef_in(coef[480]), .rdup_out(a5_wr[30]), .rdlo_out(a5_wr[94]));
			radix2 #(.width(width)) rd_st4_31  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[31]), .rdlo_in(a4_wr[95]),  .coef_in(coef[496]), .rdup_out(a5_wr[31]), .rdlo_out(a5_wr[95]));
			radix2 #(.width(width)) rd_st4_32  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[32]), .rdlo_in(a4_wr[96]),  .coef_in(coef[512]), .rdup_out(a5_wr[32]), .rdlo_out(a5_wr[96]));
			radix2 #(.width(width)) rd_st4_33  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[33]), .rdlo_in(a4_wr[97]),  .coef_in(coef[528]), .rdup_out(a5_wr[33]), .rdlo_out(a5_wr[97]));
			radix2 #(.width(width)) rd_st4_34  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[34]), .rdlo_in(a4_wr[98]),  .coef_in(coef[544]), .rdup_out(a5_wr[34]), .rdlo_out(a5_wr[98]));
			radix2 #(.width(width)) rd_st4_35  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[35]), .rdlo_in(a4_wr[99]),  .coef_in(coef[560]), .rdup_out(a5_wr[35]), .rdlo_out(a5_wr[99]));
			radix2 #(.width(width)) rd_st4_36  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[36]), .rdlo_in(a4_wr[100]),  .coef_in(coef[576]), .rdup_out(a5_wr[36]), .rdlo_out(a5_wr[100]));
			radix2 #(.width(width)) rd_st4_37  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[37]), .rdlo_in(a4_wr[101]),  .coef_in(coef[592]), .rdup_out(a5_wr[37]), .rdlo_out(a5_wr[101]));
			radix2 #(.width(width)) rd_st4_38  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[38]), .rdlo_in(a4_wr[102]),  .coef_in(coef[608]), .rdup_out(a5_wr[38]), .rdlo_out(a5_wr[102]));
			radix2 #(.width(width)) rd_st4_39  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[39]), .rdlo_in(a4_wr[103]),  .coef_in(coef[624]), .rdup_out(a5_wr[39]), .rdlo_out(a5_wr[103]));
			radix2 #(.width(width)) rd_st4_40  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[40]), .rdlo_in(a4_wr[104]),  .coef_in(coef[640]), .rdup_out(a5_wr[40]), .rdlo_out(a5_wr[104]));
			radix2 #(.width(width)) rd_st4_41  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[41]), .rdlo_in(a4_wr[105]),  .coef_in(coef[656]), .rdup_out(a5_wr[41]), .rdlo_out(a5_wr[105]));
			radix2 #(.width(width)) rd_st4_42  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[42]), .rdlo_in(a4_wr[106]),  .coef_in(coef[672]), .rdup_out(a5_wr[42]), .rdlo_out(a5_wr[106]));
			radix2 #(.width(width)) rd_st4_43  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[43]), .rdlo_in(a4_wr[107]),  .coef_in(coef[688]), .rdup_out(a5_wr[43]), .rdlo_out(a5_wr[107]));
			radix2 #(.width(width)) rd_st4_44  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[44]), .rdlo_in(a4_wr[108]),  .coef_in(coef[704]), .rdup_out(a5_wr[44]), .rdlo_out(a5_wr[108]));
			radix2 #(.width(width)) rd_st4_45  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[45]), .rdlo_in(a4_wr[109]),  .coef_in(coef[720]), .rdup_out(a5_wr[45]), .rdlo_out(a5_wr[109]));
			radix2 #(.width(width)) rd_st4_46  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[46]), .rdlo_in(a4_wr[110]),  .coef_in(coef[736]), .rdup_out(a5_wr[46]), .rdlo_out(a5_wr[110]));
			radix2 #(.width(width)) rd_st4_47  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[47]), .rdlo_in(a4_wr[111]),  .coef_in(coef[752]), .rdup_out(a5_wr[47]), .rdlo_out(a5_wr[111]));
			radix2 #(.width(width)) rd_st4_48  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[48]), .rdlo_in(a4_wr[112]),  .coef_in(coef[768]), .rdup_out(a5_wr[48]), .rdlo_out(a5_wr[112]));
			radix2 #(.width(width)) rd_st4_49  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[49]), .rdlo_in(a4_wr[113]),  .coef_in(coef[784]), .rdup_out(a5_wr[49]), .rdlo_out(a5_wr[113]));
			radix2 #(.width(width)) rd_st4_50  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[50]), .rdlo_in(a4_wr[114]),  .coef_in(coef[800]), .rdup_out(a5_wr[50]), .rdlo_out(a5_wr[114]));
			radix2 #(.width(width)) rd_st4_51  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[51]), .rdlo_in(a4_wr[115]),  .coef_in(coef[816]), .rdup_out(a5_wr[51]), .rdlo_out(a5_wr[115]));
			radix2 #(.width(width)) rd_st4_52  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[52]), .rdlo_in(a4_wr[116]),  .coef_in(coef[832]), .rdup_out(a5_wr[52]), .rdlo_out(a5_wr[116]));
			radix2 #(.width(width)) rd_st4_53  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[53]), .rdlo_in(a4_wr[117]),  .coef_in(coef[848]), .rdup_out(a5_wr[53]), .rdlo_out(a5_wr[117]));
			radix2 #(.width(width)) rd_st4_54  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[54]), .rdlo_in(a4_wr[118]),  .coef_in(coef[864]), .rdup_out(a5_wr[54]), .rdlo_out(a5_wr[118]));
			radix2 #(.width(width)) rd_st4_55  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[55]), .rdlo_in(a4_wr[119]),  .coef_in(coef[880]), .rdup_out(a5_wr[55]), .rdlo_out(a5_wr[119]));
			radix2 #(.width(width)) rd_st4_56  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[56]), .rdlo_in(a4_wr[120]),  .coef_in(coef[896]), .rdup_out(a5_wr[56]), .rdlo_out(a5_wr[120]));
			radix2 #(.width(width)) rd_st4_57  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[57]), .rdlo_in(a4_wr[121]),  .coef_in(coef[912]), .rdup_out(a5_wr[57]), .rdlo_out(a5_wr[121]));
			radix2 #(.width(width)) rd_st4_58  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[58]), .rdlo_in(a4_wr[122]),  .coef_in(coef[928]), .rdup_out(a5_wr[58]), .rdlo_out(a5_wr[122]));
			radix2 #(.width(width)) rd_st4_59  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[59]), .rdlo_in(a4_wr[123]),  .coef_in(coef[944]), .rdup_out(a5_wr[59]), .rdlo_out(a5_wr[123]));
			radix2 #(.width(width)) rd_st4_60  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[60]), .rdlo_in(a4_wr[124]),  .coef_in(coef[960]), .rdup_out(a5_wr[60]), .rdlo_out(a5_wr[124]));
			radix2 #(.width(width)) rd_st4_61  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[61]), .rdlo_in(a4_wr[125]),  .coef_in(coef[976]), .rdup_out(a5_wr[61]), .rdlo_out(a5_wr[125]));
			radix2 #(.width(width)) rd_st4_62  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[62]), .rdlo_in(a4_wr[126]),  .coef_in(coef[992]), .rdup_out(a5_wr[62]), .rdlo_out(a5_wr[126]));
			radix2 #(.width(width)) rd_st4_63  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[63]), .rdlo_in(a4_wr[127]),  .coef_in(coef[1008]), .rdup_out(a5_wr[63]), .rdlo_out(a5_wr[127]));
			radix2 #(.width(width)) rd_st4_128  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[128]), .rdlo_in(a4_wr[192]),  .coef_in(coef[0]), .rdup_out(a5_wr[128]), .rdlo_out(a5_wr[192]));
			radix2 #(.width(width)) rd_st4_129  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[129]), .rdlo_in(a4_wr[193]),  .coef_in(coef[16]), .rdup_out(a5_wr[129]), .rdlo_out(a5_wr[193]));
			radix2 #(.width(width)) rd_st4_130  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[130]), .rdlo_in(a4_wr[194]),  .coef_in(coef[32]), .rdup_out(a5_wr[130]), .rdlo_out(a5_wr[194]));
			radix2 #(.width(width)) rd_st4_131  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[131]), .rdlo_in(a4_wr[195]),  .coef_in(coef[48]), .rdup_out(a5_wr[131]), .rdlo_out(a5_wr[195]));
			radix2 #(.width(width)) rd_st4_132  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[132]), .rdlo_in(a4_wr[196]),  .coef_in(coef[64]), .rdup_out(a5_wr[132]), .rdlo_out(a5_wr[196]));
			radix2 #(.width(width)) rd_st4_133  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[133]), .rdlo_in(a4_wr[197]),  .coef_in(coef[80]), .rdup_out(a5_wr[133]), .rdlo_out(a5_wr[197]));
			radix2 #(.width(width)) rd_st4_134  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[134]), .rdlo_in(a4_wr[198]),  .coef_in(coef[96]), .rdup_out(a5_wr[134]), .rdlo_out(a5_wr[198]));
			radix2 #(.width(width)) rd_st4_135  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[135]), .rdlo_in(a4_wr[199]),  .coef_in(coef[112]), .rdup_out(a5_wr[135]), .rdlo_out(a5_wr[199]));
			radix2 #(.width(width)) rd_st4_136  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[136]), .rdlo_in(a4_wr[200]),  .coef_in(coef[128]), .rdup_out(a5_wr[136]), .rdlo_out(a5_wr[200]));
			radix2 #(.width(width)) rd_st4_137  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[137]), .rdlo_in(a4_wr[201]),  .coef_in(coef[144]), .rdup_out(a5_wr[137]), .rdlo_out(a5_wr[201]));
			radix2 #(.width(width)) rd_st4_138  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[138]), .rdlo_in(a4_wr[202]),  .coef_in(coef[160]), .rdup_out(a5_wr[138]), .rdlo_out(a5_wr[202]));
			radix2 #(.width(width)) rd_st4_139  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[139]), .rdlo_in(a4_wr[203]),  .coef_in(coef[176]), .rdup_out(a5_wr[139]), .rdlo_out(a5_wr[203]));
			radix2 #(.width(width)) rd_st4_140  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[140]), .rdlo_in(a4_wr[204]),  .coef_in(coef[192]), .rdup_out(a5_wr[140]), .rdlo_out(a5_wr[204]));
			radix2 #(.width(width)) rd_st4_141  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[141]), .rdlo_in(a4_wr[205]),  .coef_in(coef[208]), .rdup_out(a5_wr[141]), .rdlo_out(a5_wr[205]));
			radix2 #(.width(width)) rd_st4_142  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[142]), .rdlo_in(a4_wr[206]),  .coef_in(coef[224]), .rdup_out(a5_wr[142]), .rdlo_out(a5_wr[206]));
			radix2 #(.width(width)) rd_st4_143  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[143]), .rdlo_in(a4_wr[207]),  .coef_in(coef[240]), .rdup_out(a5_wr[143]), .rdlo_out(a5_wr[207]));
			radix2 #(.width(width)) rd_st4_144  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[144]), .rdlo_in(a4_wr[208]),  .coef_in(coef[256]), .rdup_out(a5_wr[144]), .rdlo_out(a5_wr[208]));
			radix2 #(.width(width)) rd_st4_145  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[145]), .rdlo_in(a4_wr[209]),  .coef_in(coef[272]), .rdup_out(a5_wr[145]), .rdlo_out(a5_wr[209]));
			radix2 #(.width(width)) rd_st4_146  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[146]), .rdlo_in(a4_wr[210]),  .coef_in(coef[288]), .rdup_out(a5_wr[146]), .rdlo_out(a5_wr[210]));
			radix2 #(.width(width)) rd_st4_147  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[147]), .rdlo_in(a4_wr[211]),  .coef_in(coef[304]), .rdup_out(a5_wr[147]), .rdlo_out(a5_wr[211]));
			radix2 #(.width(width)) rd_st4_148  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[148]), .rdlo_in(a4_wr[212]),  .coef_in(coef[320]), .rdup_out(a5_wr[148]), .rdlo_out(a5_wr[212]));
			radix2 #(.width(width)) rd_st4_149  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[149]), .rdlo_in(a4_wr[213]),  .coef_in(coef[336]), .rdup_out(a5_wr[149]), .rdlo_out(a5_wr[213]));
			radix2 #(.width(width)) rd_st4_150  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[150]), .rdlo_in(a4_wr[214]),  .coef_in(coef[352]), .rdup_out(a5_wr[150]), .rdlo_out(a5_wr[214]));
			radix2 #(.width(width)) rd_st4_151  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[151]), .rdlo_in(a4_wr[215]),  .coef_in(coef[368]), .rdup_out(a5_wr[151]), .rdlo_out(a5_wr[215]));
			radix2 #(.width(width)) rd_st4_152  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[152]), .rdlo_in(a4_wr[216]),  .coef_in(coef[384]), .rdup_out(a5_wr[152]), .rdlo_out(a5_wr[216]));
			radix2 #(.width(width)) rd_st4_153  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[153]), .rdlo_in(a4_wr[217]),  .coef_in(coef[400]), .rdup_out(a5_wr[153]), .rdlo_out(a5_wr[217]));
			radix2 #(.width(width)) rd_st4_154  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[154]), .rdlo_in(a4_wr[218]),  .coef_in(coef[416]), .rdup_out(a5_wr[154]), .rdlo_out(a5_wr[218]));
			radix2 #(.width(width)) rd_st4_155  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[155]), .rdlo_in(a4_wr[219]),  .coef_in(coef[432]), .rdup_out(a5_wr[155]), .rdlo_out(a5_wr[219]));
			radix2 #(.width(width)) rd_st4_156  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[156]), .rdlo_in(a4_wr[220]),  .coef_in(coef[448]), .rdup_out(a5_wr[156]), .rdlo_out(a5_wr[220]));
			radix2 #(.width(width)) rd_st4_157  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[157]), .rdlo_in(a4_wr[221]),  .coef_in(coef[464]), .rdup_out(a5_wr[157]), .rdlo_out(a5_wr[221]));
			radix2 #(.width(width)) rd_st4_158  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[158]), .rdlo_in(a4_wr[222]),  .coef_in(coef[480]), .rdup_out(a5_wr[158]), .rdlo_out(a5_wr[222]));
			radix2 #(.width(width)) rd_st4_159  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[159]), .rdlo_in(a4_wr[223]),  .coef_in(coef[496]), .rdup_out(a5_wr[159]), .rdlo_out(a5_wr[223]));
			radix2 #(.width(width)) rd_st4_160  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[160]), .rdlo_in(a4_wr[224]),  .coef_in(coef[512]), .rdup_out(a5_wr[160]), .rdlo_out(a5_wr[224]));
			radix2 #(.width(width)) rd_st4_161  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[161]), .rdlo_in(a4_wr[225]),  .coef_in(coef[528]), .rdup_out(a5_wr[161]), .rdlo_out(a5_wr[225]));
			radix2 #(.width(width)) rd_st4_162  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[162]), .rdlo_in(a4_wr[226]),  .coef_in(coef[544]), .rdup_out(a5_wr[162]), .rdlo_out(a5_wr[226]));
			radix2 #(.width(width)) rd_st4_163  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[163]), .rdlo_in(a4_wr[227]),  .coef_in(coef[560]), .rdup_out(a5_wr[163]), .rdlo_out(a5_wr[227]));
			radix2 #(.width(width)) rd_st4_164  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[164]), .rdlo_in(a4_wr[228]),  .coef_in(coef[576]), .rdup_out(a5_wr[164]), .rdlo_out(a5_wr[228]));
			radix2 #(.width(width)) rd_st4_165  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[165]), .rdlo_in(a4_wr[229]),  .coef_in(coef[592]), .rdup_out(a5_wr[165]), .rdlo_out(a5_wr[229]));
			radix2 #(.width(width)) rd_st4_166  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[166]), .rdlo_in(a4_wr[230]),  .coef_in(coef[608]), .rdup_out(a5_wr[166]), .rdlo_out(a5_wr[230]));
			radix2 #(.width(width)) rd_st4_167  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[167]), .rdlo_in(a4_wr[231]),  .coef_in(coef[624]), .rdup_out(a5_wr[167]), .rdlo_out(a5_wr[231]));
			radix2 #(.width(width)) rd_st4_168  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[168]), .rdlo_in(a4_wr[232]),  .coef_in(coef[640]), .rdup_out(a5_wr[168]), .rdlo_out(a5_wr[232]));
			radix2 #(.width(width)) rd_st4_169  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[169]), .rdlo_in(a4_wr[233]),  .coef_in(coef[656]), .rdup_out(a5_wr[169]), .rdlo_out(a5_wr[233]));
			radix2 #(.width(width)) rd_st4_170  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[170]), .rdlo_in(a4_wr[234]),  .coef_in(coef[672]), .rdup_out(a5_wr[170]), .rdlo_out(a5_wr[234]));
			radix2 #(.width(width)) rd_st4_171  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[171]), .rdlo_in(a4_wr[235]),  .coef_in(coef[688]), .rdup_out(a5_wr[171]), .rdlo_out(a5_wr[235]));
			radix2 #(.width(width)) rd_st4_172  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[172]), .rdlo_in(a4_wr[236]),  .coef_in(coef[704]), .rdup_out(a5_wr[172]), .rdlo_out(a5_wr[236]));
			radix2 #(.width(width)) rd_st4_173  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[173]), .rdlo_in(a4_wr[237]),  .coef_in(coef[720]), .rdup_out(a5_wr[173]), .rdlo_out(a5_wr[237]));
			radix2 #(.width(width)) rd_st4_174  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[174]), .rdlo_in(a4_wr[238]),  .coef_in(coef[736]), .rdup_out(a5_wr[174]), .rdlo_out(a5_wr[238]));
			radix2 #(.width(width)) rd_st4_175  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[175]), .rdlo_in(a4_wr[239]),  .coef_in(coef[752]), .rdup_out(a5_wr[175]), .rdlo_out(a5_wr[239]));
			radix2 #(.width(width)) rd_st4_176  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[176]), .rdlo_in(a4_wr[240]),  .coef_in(coef[768]), .rdup_out(a5_wr[176]), .rdlo_out(a5_wr[240]));
			radix2 #(.width(width)) rd_st4_177  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[177]), .rdlo_in(a4_wr[241]),  .coef_in(coef[784]), .rdup_out(a5_wr[177]), .rdlo_out(a5_wr[241]));
			radix2 #(.width(width)) rd_st4_178  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[178]), .rdlo_in(a4_wr[242]),  .coef_in(coef[800]), .rdup_out(a5_wr[178]), .rdlo_out(a5_wr[242]));
			radix2 #(.width(width)) rd_st4_179  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[179]), .rdlo_in(a4_wr[243]),  .coef_in(coef[816]), .rdup_out(a5_wr[179]), .rdlo_out(a5_wr[243]));
			radix2 #(.width(width)) rd_st4_180  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[180]), .rdlo_in(a4_wr[244]),  .coef_in(coef[832]), .rdup_out(a5_wr[180]), .rdlo_out(a5_wr[244]));
			radix2 #(.width(width)) rd_st4_181  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[181]), .rdlo_in(a4_wr[245]),  .coef_in(coef[848]), .rdup_out(a5_wr[181]), .rdlo_out(a5_wr[245]));
			radix2 #(.width(width)) rd_st4_182  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[182]), .rdlo_in(a4_wr[246]),  .coef_in(coef[864]), .rdup_out(a5_wr[182]), .rdlo_out(a5_wr[246]));
			radix2 #(.width(width)) rd_st4_183  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[183]), .rdlo_in(a4_wr[247]),  .coef_in(coef[880]), .rdup_out(a5_wr[183]), .rdlo_out(a5_wr[247]));
			radix2 #(.width(width)) rd_st4_184  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[184]), .rdlo_in(a4_wr[248]),  .coef_in(coef[896]), .rdup_out(a5_wr[184]), .rdlo_out(a5_wr[248]));
			radix2 #(.width(width)) rd_st4_185  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[185]), .rdlo_in(a4_wr[249]),  .coef_in(coef[912]), .rdup_out(a5_wr[185]), .rdlo_out(a5_wr[249]));
			radix2 #(.width(width)) rd_st4_186  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[186]), .rdlo_in(a4_wr[250]),  .coef_in(coef[928]), .rdup_out(a5_wr[186]), .rdlo_out(a5_wr[250]));
			radix2 #(.width(width)) rd_st4_187  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[187]), .rdlo_in(a4_wr[251]),  .coef_in(coef[944]), .rdup_out(a5_wr[187]), .rdlo_out(a5_wr[251]));
			radix2 #(.width(width)) rd_st4_188  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[188]), .rdlo_in(a4_wr[252]),  .coef_in(coef[960]), .rdup_out(a5_wr[188]), .rdlo_out(a5_wr[252]));
			radix2 #(.width(width)) rd_st4_189  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[189]), .rdlo_in(a4_wr[253]),  .coef_in(coef[976]), .rdup_out(a5_wr[189]), .rdlo_out(a5_wr[253]));
			radix2 #(.width(width)) rd_st4_190  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[190]), .rdlo_in(a4_wr[254]),  .coef_in(coef[992]), .rdup_out(a5_wr[190]), .rdlo_out(a5_wr[254]));
			radix2 #(.width(width)) rd_st4_191  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[191]), .rdlo_in(a4_wr[255]),  .coef_in(coef[1008]), .rdup_out(a5_wr[191]), .rdlo_out(a5_wr[255]));
			radix2 #(.width(width)) rd_st4_256  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[256]), .rdlo_in(a4_wr[320]),  .coef_in(coef[0]), .rdup_out(a5_wr[256]), .rdlo_out(a5_wr[320]));
			radix2 #(.width(width)) rd_st4_257  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[257]), .rdlo_in(a4_wr[321]),  .coef_in(coef[16]), .rdup_out(a5_wr[257]), .rdlo_out(a5_wr[321]));
			radix2 #(.width(width)) rd_st4_258  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[258]), .rdlo_in(a4_wr[322]),  .coef_in(coef[32]), .rdup_out(a5_wr[258]), .rdlo_out(a5_wr[322]));
			radix2 #(.width(width)) rd_st4_259  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[259]), .rdlo_in(a4_wr[323]),  .coef_in(coef[48]), .rdup_out(a5_wr[259]), .rdlo_out(a5_wr[323]));
			radix2 #(.width(width)) rd_st4_260  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[260]), .rdlo_in(a4_wr[324]),  .coef_in(coef[64]), .rdup_out(a5_wr[260]), .rdlo_out(a5_wr[324]));
			radix2 #(.width(width)) rd_st4_261  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[261]), .rdlo_in(a4_wr[325]),  .coef_in(coef[80]), .rdup_out(a5_wr[261]), .rdlo_out(a5_wr[325]));
			radix2 #(.width(width)) rd_st4_262  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[262]), .rdlo_in(a4_wr[326]),  .coef_in(coef[96]), .rdup_out(a5_wr[262]), .rdlo_out(a5_wr[326]));
			radix2 #(.width(width)) rd_st4_263  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[263]), .rdlo_in(a4_wr[327]),  .coef_in(coef[112]), .rdup_out(a5_wr[263]), .rdlo_out(a5_wr[327]));
			radix2 #(.width(width)) rd_st4_264  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[264]), .rdlo_in(a4_wr[328]),  .coef_in(coef[128]), .rdup_out(a5_wr[264]), .rdlo_out(a5_wr[328]));
			radix2 #(.width(width)) rd_st4_265  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[265]), .rdlo_in(a4_wr[329]),  .coef_in(coef[144]), .rdup_out(a5_wr[265]), .rdlo_out(a5_wr[329]));
			radix2 #(.width(width)) rd_st4_266  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[266]), .rdlo_in(a4_wr[330]),  .coef_in(coef[160]), .rdup_out(a5_wr[266]), .rdlo_out(a5_wr[330]));
			radix2 #(.width(width)) rd_st4_267  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[267]), .rdlo_in(a4_wr[331]),  .coef_in(coef[176]), .rdup_out(a5_wr[267]), .rdlo_out(a5_wr[331]));
			radix2 #(.width(width)) rd_st4_268  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[268]), .rdlo_in(a4_wr[332]),  .coef_in(coef[192]), .rdup_out(a5_wr[268]), .rdlo_out(a5_wr[332]));
			radix2 #(.width(width)) rd_st4_269  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[269]), .rdlo_in(a4_wr[333]),  .coef_in(coef[208]), .rdup_out(a5_wr[269]), .rdlo_out(a5_wr[333]));
			radix2 #(.width(width)) rd_st4_270  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[270]), .rdlo_in(a4_wr[334]),  .coef_in(coef[224]), .rdup_out(a5_wr[270]), .rdlo_out(a5_wr[334]));
			radix2 #(.width(width)) rd_st4_271  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[271]), .rdlo_in(a4_wr[335]),  .coef_in(coef[240]), .rdup_out(a5_wr[271]), .rdlo_out(a5_wr[335]));
			radix2 #(.width(width)) rd_st4_272  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[272]), .rdlo_in(a4_wr[336]),  .coef_in(coef[256]), .rdup_out(a5_wr[272]), .rdlo_out(a5_wr[336]));
			radix2 #(.width(width)) rd_st4_273  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[273]), .rdlo_in(a4_wr[337]),  .coef_in(coef[272]), .rdup_out(a5_wr[273]), .rdlo_out(a5_wr[337]));
			radix2 #(.width(width)) rd_st4_274  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[274]), .rdlo_in(a4_wr[338]),  .coef_in(coef[288]), .rdup_out(a5_wr[274]), .rdlo_out(a5_wr[338]));
			radix2 #(.width(width)) rd_st4_275  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[275]), .rdlo_in(a4_wr[339]),  .coef_in(coef[304]), .rdup_out(a5_wr[275]), .rdlo_out(a5_wr[339]));
			radix2 #(.width(width)) rd_st4_276  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[276]), .rdlo_in(a4_wr[340]),  .coef_in(coef[320]), .rdup_out(a5_wr[276]), .rdlo_out(a5_wr[340]));
			radix2 #(.width(width)) rd_st4_277  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[277]), .rdlo_in(a4_wr[341]),  .coef_in(coef[336]), .rdup_out(a5_wr[277]), .rdlo_out(a5_wr[341]));
			radix2 #(.width(width)) rd_st4_278  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[278]), .rdlo_in(a4_wr[342]),  .coef_in(coef[352]), .rdup_out(a5_wr[278]), .rdlo_out(a5_wr[342]));
			radix2 #(.width(width)) rd_st4_279  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[279]), .rdlo_in(a4_wr[343]),  .coef_in(coef[368]), .rdup_out(a5_wr[279]), .rdlo_out(a5_wr[343]));
			radix2 #(.width(width)) rd_st4_280  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[280]), .rdlo_in(a4_wr[344]),  .coef_in(coef[384]), .rdup_out(a5_wr[280]), .rdlo_out(a5_wr[344]));
			radix2 #(.width(width)) rd_st4_281  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[281]), .rdlo_in(a4_wr[345]),  .coef_in(coef[400]), .rdup_out(a5_wr[281]), .rdlo_out(a5_wr[345]));
			radix2 #(.width(width)) rd_st4_282  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[282]), .rdlo_in(a4_wr[346]),  .coef_in(coef[416]), .rdup_out(a5_wr[282]), .rdlo_out(a5_wr[346]));
			radix2 #(.width(width)) rd_st4_283  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[283]), .rdlo_in(a4_wr[347]),  .coef_in(coef[432]), .rdup_out(a5_wr[283]), .rdlo_out(a5_wr[347]));
			radix2 #(.width(width)) rd_st4_284  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[284]), .rdlo_in(a4_wr[348]),  .coef_in(coef[448]), .rdup_out(a5_wr[284]), .rdlo_out(a5_wr[348]));
			radix2 #(.width(width)) rd_st4_285  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[285]), .rdlo_in(a4_wr[349]),  .coef_in(coef[464]), .rdup_out(a5_wr[285]), .rdlo_out(a5_wr[349]));
			radix2 #(.width(width)) rd_st4_286  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[286]), .rdlo_in(a4_wr[350]),  .coef_in(coef[480]), .rdup_out(a5_wr[286]), .rdlo_out(a5_wr[350]));
			radix2 #(.width(width)) rd_st4_287  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[287]), .rdlo_in(a4_wr[351]),  .coef_in(coef[496]), .rdup_out(a5_wr[287]), .rdlo_out(a5_wr[351]));
			radix2 #(.width(width)) rd_st4_288  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[288]), .rdlo_in(a4_wr[352]),  .coef_in(coef[512]), .rdup_out(a5_wr[288]), .rdlo_out(a5_wr[352]));
			radix2 #(.width(width)) rd_st4_289  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[289]), .rdlo_in(a4_wr[353]),  .coef_in(coef[528]), .rdup_out(a5_wr[289]), .rdlo_out(a5_wr[353]));
			radix2 #(.width(width)) rd_st4_290  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[290]), .rdlo_in(a4_wr[354]),  .coef_in(coef[544]), .rdup_out(a5_wr[290]), .rdlo_out(a5_wr[354]));
			radix2 #(.width(width)) rd_st4_291  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[291]), .rdlo_in(a4_wr[355]),  .coef_in(coef[560]), .rdup_out(a5_wr[291]), .rdlo_out(a5_wr[355]));
			radix2 #(.width(width)) rd_st4_292  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[292]), .rdlo_in(a4_wr[356]),  .coef_in(coef[576]), .rdup_out(a5_wr[292]), .rdlo_out(a5_wr[356]));
			radix2 #(.width(width)) rd_st4_293  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[293]), .rdlo_in(a4_wr[357]),  .coef_in(coef[592]), .rdup_out(a5_wr[293]), .rdlo_out(a5_wr[357]));
			radix2 #(.width(width)) rd_st4_294  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[294]), .rdlo_in(a4_wr[358]),  .coef_in(coef[608]), .rdup_out(a5_wr[294]), .rdlo_out(a5_wr[358]));
			radix2 #(.width(width)) rd_st4_295  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[295]), .rdlo_in(a4_wr[359]),  .coef_in(coef[624]), .rdup_out(a5_wr[295]), .rdlo_out(a5_wr[359]));
			radix2 #(.width(width)) rd_st4_296  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[296]), .rdlo_in(a4_wr[360]),  .coef_in(coef[640]), .rdup_out(a5_wr[296]), .rdlo_out(a5_wr[360]));
			radix2 #(.width(width)) rd_st4_297  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[297]), .rdlo_in(a4_wr[361]),  .coef_in(coef[656]), .rdup_out(a5_wr[297]), .rdlo_out(a5_wr[361]));
			radix2 #(.width(width)) rd_st4_298  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[298]), .rdlo_in(a4_wr[362]),  .coef_in(coef[672]), .rdup_out(a5_wr[298]), .rdlo_out(a5_wr[362]));
			radix2 #(.width(width)) rd_st4_299  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[299]), .rdlo_in(a4_wr[363]),  .coef_in(coef[688]), .rdup_out(a5_wr[299]), .rdlo_out(a5_wr[363]));
			radix2 #(.width(width)) rd_st4_300  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[300]), .rdlo_in(a4_wr[364]),  .coef_in(coef[704]), .rdup_out(a5_wr[300]), .rdlo_out(a5_wr[364]));
			radix2 #(.width(width)) rd_st4_301  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[301]), .rdlo_in(a4_wr[365]),  .coef_in(coef[720]), .rdup_out(a5_wr[301]), .rdlo_out(a5_wr[365]));
			radix2 #(.width(width)) rd_st4_302  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[302]), .rdlo_in(a4_wr[366]),  .coef_in(coef[736]), .rdup_out(a5_wr[302]), .rdlo_out(a5_wr[366]));
			radix2 #(.width(width)) rd_st4_303  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[303]), .rdlo_in(a4_wr[367]),  .coef_in(coef[752]), .rdup_out(a5_wr[303]), .rdlo_out(a5_wr[367]));
			radix2 #(.width(width)) rd_st4_304  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[304]), .rdlo_in(a4_wr[368]),  .coef_in(coef[768]), .rdup_out(a5_wr[304]), .rdlo_out(a5_wr[368]));
			radix2 #(.width(width)) rd_st4_305  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[305]), .rdlo_in(a4_wr[369]),  .coef_in(coef[784]), .rdup_out(a5_wr[305]), .rdlo_out(a5_wr[369]));
			radix2 #(.width(width)) rd_st4_306  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[306]), .rdlo_in(a4_wr[370]),  .coef_in(coef[800]), .rdup_out(a5_wr[306]), .rdlo_out(a5_wr[370]));
			radix2 #(.width(width)) rd_st4_307  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[307]), .rdlo_in(a4_wr[371]),  .coef_in(coef[816]), .rdup_out(a5_wr[307]), .rdlo_out(a5_wr[371]));
			radix2 #(.width(width)) rd_st4_308  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[308]), .rdlo_in(a4_wr[372]),  .coef_in(coef[832]), .rdup_out(a5_wr[308]), .rdlo_out(a5_wr[372]));
			radix2 #(.width(width)) rd_st4_309  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[309]), .rdlo_in(a4_wr[373]),  .coef_in(coef[848]), .rdup_out(a5_wr[309]), .rdlo_out(a5_wr[373]));
			radix2 #(.width(width)) rd_st4_310  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[310]), .rdlo_in(a4_wr[374]),  .coef_in(coef[864]), .rdup_out(a5_wr[310]), .rdlo_out(a5_wr[374]));
			radix2 #(.width(width)) rd_st4_311  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[311]), .rdlo_in(a4_wr[375]),  .coef_in(coef[880]), .rdup_out(a5_wr[311]), .rdlo_out(a5_wr[375]));
			radix2 #(.width(width)) rd_st4_312  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[312]), .rdlo_in(a4_wr[376]),  .coef_in(coef[896]), .rdup_out(a5_wr[312]), .rdlo_out(a5_wr[376]));
			radix2 #(.width(width)) rd_st4_313  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[313]), .rdlo_in(a4_wr[377]),  .coef_in(coef[912]), .rdup_out(a5_wr[313]), .rdlo_out(a5_wr[377]));
			radix2 #(.width(width)) rd_st4_314  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[314]), .rdlo_in(a4_wr[378]),  .coef_in(coef[928]), .rdup_out(a5_wr[314]), .rdlo_out(a5_wr[378]));
			radix2 #(.width(width)) rd_st4_315  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[315]), .rdlo_in(a4_wr[379]),  .coef_in(coef[944]), .rdup_out(a5_wr[315]), .rdlo_out(a5_wr[379]));
			radix2 #(.width(width)) rd_st4_316  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[316]), .rdlo_in(a4_wr[380]),  .coef_in(coef[960]), .rdup_out(a5_wr[316]), .rdlo_out(a5_wr[380]));
			radix2 #(.width(width)) rd_st4_317  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[317]), .rdlo_in(a4_wr[381]),  .coef_in(coef[976]), .rdup_out(a5_wr[317]), .rdlo_out(a5_wr[381]));
			radix2 #(.width(width)) rd_st4_318  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[318]), .rdlo_in(a4_wr[382]),  .coef_in(coef[992]), .rdup_out(a5_wr[318]), .rdlo_out(a5_wr[382]));
			radix2 #(.width(width)) rd_st4_319  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[319]), .rdlo_in(a4_wr[383]),  .coef_in(coef[1008]), .rdup_out(a5_wr[319]), .rdlo_out(a5_wr[383]));
			radix2 #(.width(width)) rd_st4_384  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[384]), .rdlo_in(a4_wr[448]),  .coef_in(coef[0]), .rdup_out(a5_wr[384]), .rdlo_out(a5_wr[448]));
			radix2 #(.width(width)) rd_st4_385  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[385]), .rdlo_in(a4_wr[449]),  .coef_in(coef[16]), .rdup_out(a5_wr[385]), .rdlo_out(a5_wr[449]));
			radix2 #(.width(width)) rd_st4_386  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[386]), .rdlo_in(a4_wr[450]),  .coef_in(coef[32]), .rdup_out(a5_wr[386]), .rdlo_out(a5_wr[450]));
			radix2 #(.width(width)) rd_st4_387  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[387]), .rdlo_in(a4_wr[451]),  .coef_in(coef[48]), .rdup_out(a5_wr[387]), .rdlo_out(a5_wr[451]));
			radix2 #(.width(width)) rd_st4_388  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[388]), .rdlo_in(a4_wr[452]),  .coef_in(coef[64]), .rdup_out(a5_wr[388]), .rdlo_out(a5_wr[452]));
			radix2 #(.width(width)) rd_st4_389  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[389]), .rdlo_in(a4_wr[453]),  .coef_in(coef[80]), .rdup_out(a5_wr[389]), .rdlo_out(a5_wr[453]));
			radix2 #(.width(width)) rd_st4_390  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[390]), .rdlo_in(a4_wr[454]),  .coef_in(coef[96]), .rdup_out(a5_wr[390]), .rdlo_out(a5_wr[454]));
			radix2 #(.width(width)) rd_st4_391  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[391]), .rdlo_in(a4_wr[455]),  .coef_in(coef[112]), .rdup_out(a5_wr[391]), .rdlo_out(a5_wr[455]));
			radix2 #(.width(width)) rd_st4_392  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[392]), .rdlo_in(a4_wr[456]),  .coef_in(coef[128]), .rdup_out(a5_wr[392]), .rdlo_out(a5_wr[456]));
			radix2 #(.width(width)) rd_st4_393  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[393]), .rdlo_in(a4_wr[457]),  .coef_in(coef[144]), .rdup_out(a5_wr[393]), .rdlo_out(a5_wr[457]));
			radix2 #(.width(width)) rd_st4_394  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[394]), .rdlo_in(a4_wr[458]),  .coef_in(coef[160]), .rdup_out(a5_wr[394]), .rdlo_out(a5_wr[458]));
			radix2 #(.width(width)) rd_st4_395  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[395]), .rdlo_in(a4_wr[459]),  .coef_in(coef[176]), .rdup_out(a5_wr[395]), .rdlo_out(a5_wr[459]));
			radix2 #(.width(width)) rd_st4_396  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[396]), .rdlo_in(a4_wr[460]),  .coef_in(coef[192]), .rdup_out(a5_wr[396]), .rdlo_out(a5_wr[460]));
			radix2 #(.width(width)) rd_st4_397  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[397]), .rdlo_in(a4_wr[461]),  .coef_in(coef[208]), .rdup_out(a5_wr[397]), .rdlo_out(a5_wr[461]));
			radix2 #(.width(width)) rd_st4_398  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[398]), .rdlo_in(a4_wr[462]),  .coef_in(coef[224]), .rdup_out(a5_wr[398]), .rdlo_out(a5_wr[462]));
			radix2 #(.width(width)) rd_st4_399  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[399]), .rdlo_in(a4_wr[463]),  .coef_in(coef[240]), .rdup_out(a5_wr[399]), .rdlo_out(a5_wr[463]));
			radix2 #(.width(width)) rd_st4_400  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[400]), .rdlo_in(a4_wr[464]),  .coef_in(coef[256]), .rdup_out(a5_wr[400]), .rdlo_out(a5_wr[464]));
			radix2 #(.width(width)) rd_st4_401  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[401]), .rdlo_in(a4_wr[465]),  .coef_in(coef[272]), .rdup_out(a5_wr[401]), .rdlo_out(a5_wr[465]));
			radix2 #(.width(width)) rd_st4_402  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[402]), .rdlo_in(a4_wr[466]),  .coef_in(coef[288]), .rdup_out(a5_wr[402]), .rdlo_out(a5_wr[466]));
			radix2 #(.width(width)) rd_st4_403  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[403]), .rdlo_in(a4_wr[467]),  .coef_in(coef[304]), .rdup_out(a5_wr[403]), .rdlo_out(a5_wr[467]));
			radix2 #(.width(width)) rd_st4_404  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[404]), .rdlo_in(a4_wr[468]),  .coef_in(coef[320]), .rdup_out(a5_wr[404]), .rdlo_out(a5_wr[468]));
			radix2 #(.width(width)) rd_st4_405  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[405]), .rdlo_in(a4_wr[469]),  .coef_in(coef[336]), .rdup_out(a5_wr[405]), .rdlo_out(a5_wr[469]));
			radix2 #(.width(width)) rd_st4_406  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[406]), .rdlo_in(a4_wr[470]),  .coef_in(coef[352]), .rdup_out(a5_wr[406]), .rdlo_out(a5_wr[470]));
			radix2 #(.width(width)) rd_st4_407  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[407]), .rdlo_in(a4_wr[471]),  .coef_in(coef[368]), .rdup_out(a5_wr[407]), .rdlo_out(a5_wr[471]));
			radix2 #(.width(width)) rd_st4_408  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[408]), .rdlo_in(a4_wr[472]),  .coef_in(coef[384]), .rdup_out(a5_wr[408]), .rdlo_out(a5_wr[472]));
			radix2 #(.width(width)) rd_st4_409  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[409]), .rdlo_in(a4_wr[473]),  .coef_in(coef[400]), .rdup_out(a5_wr[409]), .rdlo_out(a5_wr[473]));
			radix2 #(.width(width)) rd_st4_410  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[410]), .rdlo_in(a4_wr[474]),  .coef_in(coef[416]), .rdup_out(a5_wr[410]), .rdlo_out(a5_wr[474]));
			radix2 #(.width(width)) rd_st4_411  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[411]), .rdlo_in(a4_wr[475]),  .coef_in(coef[432]), .rdup_out(a5_wr[411]), .rdlo_out(a5_wr[475]));
			radix2 #(.width(width)) rd_st4_412  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[412]), .rdlo_in(a4_wr[476]),  .coef_in(coef[448]), .rdup_out(a5_wr[412]), .rdlo_out(a5_wr[476]));
			radix2 #(.width(width)) rd_st4_413  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[413]), .rdlo_in(a4_wr[477]),  .coef_in(coef[464]), .rdup_out(a5_wr[413]), .rdlo_out(a5_wr[477]));
			radix2 #(.width(width)) rd_st4_414  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[414]), .rdlo_in(a4_wr[478]),  .coef_in(coef[480]), .rdup_out(a5_wr[414]), .rdlo_out(a5_wr[478]));
			radix2 #(.width(width)) rd_st4_415  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[415]), .rdlo_in(a4_wr[479]),  .coef_in(coef[496]), .rdup_out(a5_wr[415]), .rdlo_out(a5_wr[479]));
			radix2 #(.width(width)) rd_st4_416  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[416]), .rdlo_in(a4_wr[480]),  .coef_in(coef[512]), .rdup_out(a5_wr[416]), .rdlo_out(a5_wr[480]));
			radix2 #(.width(width)) rd_st4_417  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[417]), .rdlo_in(a4_wr[481]),  .coef_in(coef[528]), .rdup_out(a5_wr[417]), .rdlo_out(a5_wr[481]));
			radix2 #(.width(width)) rd_st4_418  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[418]), .rdlo_in(a4_wr[482]),  .coef_in(coef[544]), .rdup_out(a5_wr[418]), .rdlo_out(a5_wr[482]));
			radix2 #(.width(width)) rd_st4_419  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[419]), .rdlo_in(a4_wr[483]),  .coef_in(coef[560]), .rdup_out(a5_wr[419]), .rdlo_out(a5_wr[483]));
			radix2 #(.width(width)) rd_st4_420  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[420]), .rdlo_in(a4_wr[484]),  .coef_in(coef[576]), .rdup_out(a5_wr[420]), .rdlo_out(a5_wr[484]));
			radix2 #(.width(width)) rd_st4_421  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[421]), .rdlo_in(a4_wr[485]),  .coef_in(coef[592]), .rdup_out(a5_wr[421]), .rdlo_out(a5_wr[485]));
			radix2 #(.width(width)) rd_st4_422  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[422]), .rdlo_in(a4_wr[486]),  .coef_in(coef[608]), .rdup_out(a5_wr[422]), .rdlo_out(a5_wr[486]));
			radix2 #(.width(width)) rd_st4_423  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[423]), .rdlo_in(a4_wr[487]),  .coef_in(coef[624]), .rdup_out(a5_wr[423]), .rdlo_out(a5_wr[487]));
			radix2 #(.width(width)) rd_st4_424  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[424]), .rdlo_in(a4_wr[488]),  .coef_in(coef[640]), .rdup_out(a5_wr[424]), .rdlo_out(a5_wr[488]));
			radix2 #(.width(width)) rd_st4_425  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[425]), .rdlo_in(a4_wr[489]),  .coef_in(coef[656]), .rdup_out(a5_wr[425]), .rdlo_out(a5_wr[489]));
			radix2 #(.width(width)) rd_st4_426  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[426]), .rdlo_in(a4_wr[490]),  .coef_in(coef[672]), .rdup_out(a5_wr[426]), .rdlo_out(a5_wr[490]));
			radix2 #(.width(width)) rd_st4_427  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[427]), .rdlo_in(a4_wr[491]),  .coef_in(coef[688]), .rdup_out(a5_wr[427]), .rdlo_out(a5_wr[491]));
			radix2 #(.width(width)) rd_st4_428  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[428]), .rdlo_in(a4_wr[492]),  .coef_in(coef[704]), .rdup_out(a5_wr[428]), .rdlo_out(a5_wr[492]));
			radix2 #(.width(width)) rd_st4_429  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[429]), .rdlo_in(a4_wr[493]),  .coef_in(coef[720]), .rdup_out(a5_wr[429]), .rdlo_out(a5_wr[493]));
			radix2 #(.width(width)) rd_st4_430  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[430]), .rdlo_in(a4_wr[494]),  .coef_in(coef[736]), .rdup_out(a5_wr[430]), .rdlo_out(a5_wr[494]));
			radix2 #(.width(width)) rd_st4_431  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[431]), .rdlo_in(a4_wr[495]),  .coef_in(coef[752]), .rdup_out(a5_wr[431]), .rdlo_out(a5_wr[495]));
			radix2 #(.width(width)) rd_st4_432  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[432]), .rdlo_in(a4_wr[496]),  .coef_in(coef[768]), .rdup_out(a5_wr[432]), .rdlo_out(a5_wr[496]));
			radix2 #(.width(width)) rd_st4_433  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[433]), .rdlo_in(a4_wr[497]),  .coef_in(coef[784]), .rdup_out(a5_wr[433]), .rdlo_out(a5_wr[497]));
			radix2 #(.width(width)) rd_st4_434  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[434]), .rdlo_in(a4_wr[498]),  .coef_in(coef[800]), .rdup_out(a5_wr[434]), .rdlo_out(a5_wr[498]));
			radix2 #(.width(width)) rd_st4_435  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[435]), .rdlo_in(a4_wr[499]),  .coef_in(coef[816]), .rdup_out(a5_wr[435]), .rdlo_out(a5_wr[499]));
			radix2 #(.width(width)) rd_st4_436  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[436]), .rdlo_in(a4_wr[500]),  .coef_in(coef[832]), .rdup_out(a5_wr[436]), .rdlo_out(a5_wr[500]));
			radix2 #(.width(width)) rd_st4_437  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[437]), .rdlo_in(a4_wr[501]),  .coef_in(coef[848]), .rdup_out(a5_wr[437]), .rdlo_out(a5_wr[501]));
			radix2 #(.width(width)) rd_st4_438  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[438]), .rdlo_in(a4_wr[502]),  .coef_in(coef[864]), .rdup_out(a5_wr[438]), .rdlo_out(a5_wr[502]));
			radix2 #(.width(width)) rd_st4_439  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[439]), .rdlo_in(a4_wr[503]),  .coef_in(coef[880]), .rdup_out(a5_wr[439]), .rdlo_out(a5_wr[503]));
			radix2 #(.width(width)) rd_st4_440  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[440]), .rdlo_in(a4_wr[504]),  .coef_in(coef[896]), .rdup_out(a5_wr[440]), .rdlo_out(a5_wr[504]));
			radix2 #(.width(width)) rd_st4_441  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[441]), .rdlo_in(a4_wr[505]),  .coef_in(coef[912]), .rdup_out(a5_wr[441]), .rdlo_out(a5_wr[505]));
			radix2 #(.width(width)) rd_st4_442  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[442]), .rdlo_in(a4_wr[506]),  .coef_in(coef[928]), .rdup_out(a5_wr[442]), .rdlo_out(a5_wr[506]));
			radix2 #(.width(width)) rd_st4_443  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[443]), .rdlo_in(a4_wr[507]),  .coef_in(coef[944]), .rdup_out(a5_wr[443]), .rdlo_out(a5_wr[507]));
			radix2 #(.width(width)) rd_st4_444  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[444]), .rdlo_in(a4_wr[508]),  .coef_in(coef[960]), .rdup_out(a5_wr[444]), .rdlo_out(a5_wr[508]));
			radix2 #(.width(width)) rd_st4_445  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[445]), .rdlo_in(a4_wr[509]),  .coef_in(coef[976]), .rdup_out(a5_wr[445]), .rdlo_out(a5_wr[509]));
			radix2 #(.width(width)) rd_st4_446  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[446]), .rdlo_in(a4_wr[510]),  .coef_in(coef[992]), .rdup_out(a5_wr[446]), .rdlo_out(a5_wr[510]));
			radix2 #(.width(width)) rd_st4_447  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[447]), .rdlo_in(a4_wr[511]),  .coef_in(coef[1008]), .rdup_out(a5_wr[447]), .rdlo_out(a5_wr[511]));
			radix2 #(.width(width)) rd_st4_512  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[512]), .rdlo_in(a4_wr[576]),  .coef_in(coef[0]), .rdup_out(a5_wr[512]), .rdlo_out(a5_wr[576]));
			radix2 #(.width(width)) rd_st4_513  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[513]), .rdlo_in(a4_wr[577]),  .coef_in(coef[16]), .rdup_out(a5_wr[513]), .rdlo_out(a5_wr[577]));
			radix2 #(.width(width)) rd_st4_514  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[514]), .rdlo_in(a4_wr[578]),  .coef_in(coef[32]), .rdup_out(a5_wr[514]), .rdlo_out(a5_wr[578]));
			radix2 #(.width(width)) rd_st4_515  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[515]), .rdlo_in(a4_wr[579]),  .coef_in(coef[48]), .rdup_out(a5_wr[515]), .rdlo_out(a5_wr[579]));
			radix2 #(.width(width)) rd_st4_516  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[516]), .rdlo_in(a4_wr[580]),  .coef_in(coef[64]), .rdup_out(a5_wr[516]), .rdlo_out(a5_wr[580]));
			radix2 #(.width(width)) rd_st4_517  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[517]), .rdlo_in(a4_wr[581]),  .coef_in(coef[80]), .rdup_out(a5_wr[517]), .rdlo_out(a5_wr[581]));
			radix2 #(.width(width)) rd_st4_518  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[518]), .rdlo_in(a4_wr[582]),  .coef_in(coef[96]), .rdup_out(a5_wr[518]), .rdlo_out(a5_wr[582]));
			radix2 #(.width(width)) rd_st4_519  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[519]), .rdlo_in(a4_wr[583]),  .coef_in(coef[112]), .rdup_out(a5_wr[519]), .rdlo_out(a5_wr[583]));
			radix2 #(.width(width)) rd_st4_520  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[520]), .rdlo_in(a4_wr[584]),  .coef_in(coef[128]), .rdup_out(a5_wr[520]), .rdlo_out(a5_wr[584]));
			radix2 #(.width(width)) rd_st4_521  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[521]), .rdlo_in(a4_wr[585]),  .coef_in(coef[144]), .rdup_out(a5_wr[521]), .rdlo_out(a5_wr[585]));
			radix2 #(.width(width)) rd_st4_522  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[522]), .rdlo_in(a4_wr[586]),  .coef_in(coef[160]), .rdup_out(a5_wr[522]), .rdlo_out(a5_wr[586]));
			radix2 #(.width(width)) rd_st4_523  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[523]), .rdlo_in(a4_wr[587]),  .coef_in(coef[176]), .rdup_out(a5_wr[523]), .rdlo_out(a5_wr[587]));
			radix2 #(.width(width)) rd_st4_524  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[524]), .rdlo_in(a4_wr[588]),  .coef_in(coef[192]), .rdup_out(a5_wr[524]), .rdlo_out(a5_wr[588]));
			radix2 #(.width(width)) rd_st4_525  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[525]), .rdlo_in(a4_wr[589]),  .coef_in(coef[208]), .rdup_out(a5_wr[525]), .rdlo_out(a5_wr[589]));
			radix2 #(.width(width)) rd_st4_526  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[526]), .rdlo_in(a4_wr[590]),  .coef_in(coef[224]), .rdup_out(a5_wr[526]), .rdlo_out(a5_wr[590]));
			radix2 #(.width(width)) rd_st4_527  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[527]), .rdlo_in(a4_wr[591]),  .coef_in(coef[240]), .rdup_out(a5_wr[527]), .rdlo_out(a5_wr[591]));
			radix2 #(.width(width)) rd_st4_528  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[528]), .rdlo_in(a4_wr[592]),  .coef_in(coef[256]), .rdup_out(a5_wr[528]), .rdlo_out(a5_wr[592]));
			radix2 #(.width(width)) rd_st4_529  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[529]), .rdlo_in(a4_wr[593]),  .coef_in(coef[272]), .rdup_out(a5_wr[529]), .rdlo_out(a5_wr[593]));
			radix2 #(.width(width)) rd_st4_530  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[530]), .rdlo_in(a4_wr[594]),  .coef_in(coef[288]), .rdup_out(a5_wr[530]), .rdlo_out(a5_wr[594]));
			radix2 #(.width(width)) rd_st4_531  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[531]), .rdlo_in(a4_wr[595]),  .coef_in(coef[304]), .rdup_out(a5_wr[531]), .rdlo_out(a5_wr[595]));
			radix2 #(.width(width)) rd_st4_532  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[532]), .rdlo_in(a4_wr[596]),  .coef_in(coef[320]), .rdup_out(a5_wr[532]), .rdlo_out(a5_wr[596]));
			radix2 #(.width(width)) rd_st4_533  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[533]), .rdlo_in(a4_wr[597]),  .coef_in(coef[336]), .rdup_out(a5_wr[533]), .rdlo_out(a5_wr[597]));
			radix2 #(.width(width)) rd_st4_534  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[534]), .rdlo_in(a4_wr[598]),  .coef_in(coef[352]), .rdup_out(a5_wr[534]), .rdlo_out(a5_wr[598]));
			radix2 #(.width(width)) rd_st4_535  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[535]), .rdlo_in(a4_wr[599]),  .coef_in(coef[368]), .rdup_out(a5_wr[535]), .rdlo_out(a5_wr[599]));
			radix2 #(.width(width)) rd_st4_536  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[536]), .rdlo_in(a4_wr[600]),  .coef_in(coef[384]), .rdup_out(a5_wr[536]), .rdlo_out(a5_wr[600]));
			radix2 #(.width(width)) rd_st4_537  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[537]), .rdlo_in(a4_wr[601]),  .coef_in(coef[400]), .rdup_out(a5_wr[537]), .rdlo_out(a5_wr[601]));
			radix2 #(.width(width)) rd_st4_538  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[538]), .rdlo_in(a4_wr[602]),  .coef_in(coef[416]), .rdup_out(a5_wr[538]), .rdlo_out(a5_wr[602]));
			radix2 #(.width(width)) rd_st4_539  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[539]), .rdlo_in(a4_wr[603]),  .coef_in(coef[432]), .rdup_out(a5_wr[539]), .rdlo_out(a5_wr[603]));
			radix2 #(.width(width)) rd_st4_540  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[540]), .rdlo_in(a4_wr[604]),  .coef_in(coef[448]), .rdup_out(a5_wr[540]), .rdlo_out(a5_wr[604]));
			radix2 #(.width(width)) rd_st4_541  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[541]), .rdlo_in(a4_wr[605]),  .coef_in(coef[464]), .rdup_out(a5_wr[541]), .rdlo_out(a5_wr[605]));
			radix2 #(.width(width)) rd_st4_542  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[542]), .rdlo_in(a4_wr[606]),  .coef_in(coef[480]), .rdup_out(a5_wr[542]), .rdlo_out(a5_wr[606]));
			radix2 #(.width(width)) rd_st4_543  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[543]), .rdlo_in(a4_wr[607]),  .coef_in(coef[496]), .rdup_out(a5_wr[543]), .rdlo_out(a5_wr[607]));
			radix2 #(.width(width)) rd_st4_544  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[544]), .rdlo_in(a4_wr[608]),  .coef_in(coef[512]), .rdup_out(a5_wr[544]), .rdlo_out(a5_wr[608]));
			radix2 #(.width(width)) rd_st4_545  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[545]), .rdlo_in(a4_wr[609]),  .coef_in(coef[528]), .rdup_out(a5_wr[545]), .rdlo_out(a5_wr[609]));
			radix2 #(.width(width)) rd_st4_546  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[546]), .rdlo_in(a4_wr[610]),  .coef_in(coef[544]), .rdup_out(a5_wr[546]), .rdlo_out(a5_wr[610]));
			radix2 #(.width(width)) rd_st4_547  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[547]), .rdlo_in(a4_wr[611]),  .coef_in(coef[560]), .rdup_out(a5_wr[547]), .rdlo_out(a5_wr[611]));
			radix2 #(.width(width)) rd_st4_548  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[548]), .rdlo_in(a4_wr[612]),  .coef_in(coef[576]), .rdup_out(a5_wr[548]), .rdlo_out(a5_wr[612]));
			radix2 #(.width(width)) rd_st4_549  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[549]), .rdlo_in(a4_wr[613]),  .coef_in(coef[592]), .rdup_out(a5_wr[549]), .rdlo_out(a5_wr[613]));
			radix2 #(.width(width)) rd_st4_550  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[550]), .rdlo_in(a4_wr[614]),  .coef_in(coef[608]), .rdup_out(a5_wr[550]), .rdlo_out(a5_wr[614]));
			radix2 #(.width(width)) rd_st4_551  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[551]), .rdlo_in(a4_wr[615]),  .coef_in(coef[624]), .rdup_out(a5_wr[551]), .rdlo_out(a5_wr[615]));
			radix2 #(.width(width)) rd_st4_552  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[552]), .rdlo_in(a4_wr[616]),  .coef_in(coef[640]), .rdup_out(a5_wr[552]), .rdlo_out(a5_wr[616]));
			radix2 #(.width(width)) rd_st4_553  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[553]), .rdlo_in(a4_wr[617]),  .coef_in(coef[656]), .rdup_out(a5_wr[553]), .rdlo_out(a5_wr[617]));
			radix2 #(.width(width)) rd_st4_554  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[554]), .rdlo_in(a4_wr[618]),  .coef_in(coef[672]), .rdup_out(a5_wr[554]), .rdlo_out(a5_wr[618]));
			radix2 #(.width(width)) rd_st4_555  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[555]), .rdlo_in(a4_wr[619]),  .coef_in(coef[688]), .rdup_out(a5_wr[555]), .rdlo_out(a5_wr[619]));
			radix2 #(.width(width)) rd_st4_556  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[556]), .rdlo_in(a4_wr[620]),  .coef_in(coef[704]), .rdup_out(a5_wr[556]), .rdlo_out(a5_wr[620]));
			radix2 #(.width(width)) rd_st4_557  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[557]), .rdlo_in(a4_wr[621]),  .coef_in(coef[720]), .rdup_out(a5_wr[557]), .rdlo_out(a5_wr[621]));
			radix2 #(.width(width)) rd_st4_558  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[558]), .rdlo_in(a4_wr[622]),  .coef_in(coef[736]), .rdup_out(a5_wr[558]), .rdlo_out(a5_wr[622]));
			radix2 #(.width(width)) rd_st4_559  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[559]), .rdlo_in(a4_wr[623]),  .coef_in(coef[752]), .rdup_out(a5_wr[559]), .rdlo_out(a5_wr[623]));
			radix2 #(.width(width)) rd_st4_560  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[560]), .rdlo_in(a4_wr[624]),  .coef_in(coef[768]), .rdup_out(a5_wr[560]), .rdlo_out(a5_wr[624]));
			radix2 #(.width(width)) rd_st4_561  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[561]), .rdlo_in(a4_wr[625]),  .coef_in(coef[784]), .rdup_out(a5_wr[561]), .rdlo_out(a5_wr[625]));
			radix2 #(.width(width)) rd_st4_562  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[562]), .rdlo_in(a4_wr[626]),  .coef_in(coef[800]), .rdup_out(a5_wr[562]), .rdlo_out(a5_wr[626]));
			radix2 #(.width(width)) rd_st4_563  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[563]), .rdlo_in(a4_wr[627]),  .coef_in(coef[816]), .rdup_out(a5_wr[563]), .rdlo_out(a5_wr[627]));
			radix2 #(.width(width)) rd_st4_564  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[564]), .rdlo_in(a4_wr[628]),  .coef_in(coef[832]), .rdup_out(a5_wr[564]), .rdlo_out(a5_wr[628]));
			radix2 #(.width(width)) rd_st4_565  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[565]), .rdlo_in(a4_wr[629]),  .coef_in(coef[848]), .rdup_out(a5_wr[565]), .rdlo_out(a5_wr[629]));
			radix2 #(.width(width)) rd_st4_566  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[566]), .rdlo_in(a4_wr[630]),  .coef_in(coef[864]), .rdup_out(a5_wr[566]), .rdlo_out(a5_wr[630]));
			radix2 #(.width(width)) rd_st4_567  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[567]), .rdlo_in(a4_wr[631]),  .coef_in(coef[880]), .rdup_out(a5_wr[567]), .rdlo_out(a5_wr[631]));
			radix2 #(.width(width)) rd_st4_568  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[568]), .rdlo_in(a4_wr[632]),  .coef_in(coef[896]), .rdup_out(a5_wr[568]), .rdlo_out(a5_wr[632]));
			radix2 #(.width(width)) rd_st4_569  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[569]), .rdlo_in(a4_wr[633]),  .coef_in(coef[912]), .rdup_out(a5_wr[569]), .rdlo_out(a5_wr[633]));
			radix2 #(.width(width)) rd_st4_570  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[570]), .rdlo_in(a4_wr[634]),  .coef_in(coef[928]), .rdup_out(a5_wr[570]), .rdlo_out(a5_wr[634]));
			radix2 #(.width(width)) rd_st4_571  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[571]), .rdlo_in(a4_wr[635]),  .coef_in(coef[944]), .rdup_out(a5_wr[571]), .rdlo_out(a5_wr[635]));
			radix2 #(.width(width)) rd_st4_572  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[572]), .rdlo_in(a4_wr[636]),  .coef_in(coef[960]), .rdup_out(a5_wr[572]), .rdlo_out(a5_wr[636]));
			radix2 #(.width(width)) rd_st4_573  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[573]), .rdlo_in(a4_wr[637]),  .coef_in(coef[976]), .rdup_out(a5_wr[573]), .rdlo_out(a5_wr[637]));
			radix2 #(.width(width)) rd_st4_574  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[574]), .rdlo_in(a4_wr[638]),  .coef_in(coef[992]), .rdup_out(a5_wr[574]), .rdlo_out(a5_wr[638]));
			radix2 #(.width(width)) rd_st4_575  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[575]), .rdlo_in(a4_wr[639]),  .coef_in(coef[1008]), .rdup_out(a5_wr[575]), .rdlo_out(a5_wr[639]));
			radix2 #(.width(width)) rd_st4_640  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[640]), .rdlo_in(a4_wr[704]),  .coef_in(coef[0]), .rdup_out(a5_wr[640]), .rdlo_out(a5_wr[704]));
			radix2 #(.width(width)) rd_st4_641  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[641]), .rdlo_in(a4_wr[705]),  .coef_in(coef[16]), .rdup_out(a5_wr[641]), .rdlo_out(a5_wr[705]));
			radix2 #(.width(width)) rd_st4_642  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[642]), .rdlo_in(a4_wr[706]),  .coef_in(coef[32]), .rdup_out(a5_wr[642]), .rdlo_out(a5_wr[706]));
			radix2 #(.width(width)) rd_st4_643  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[643]), .rdlo_in(a4_wr[707]),  .coef_in(coef[48]), .rdup_out(a5_wr[643]), .rdlo_out(a5_wr[707]));
			radix2 #(.width(width)) rd_st4_644  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[644]), .rdlo_in(a4_wr[708]),  .coef_in(coef[64]), .rdup_out(a5_wr[644]), .rdlo_out(a5_wr[708]));
			radix2 #(.width(width)) rd_st4_645  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[645]), .rdlo_in(a4_wr[709]),  .coef_in(coef[80]), .rdup_out(a5_wr[645]), .rdlo_out(a5_wr[709]));
			radix2 #(.width(width)) rd_st4_646  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[646]), .rdlo_in(a4_wr[710]),  .coef_in(coef[96]), .rdup_out(a5_wr[646]), .rdlo_out(a5_wr[710]));
			radix2 #(.width(width)) rd_st4_647  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[647]), .rdlo_in(a4_wr[711]),  .coef_in(coef[112]), .rdup_out(a5_wr[647]), .rdlo_out(a5_wr[711]));
			radix2 #(.width(width)) rd_st4_648  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[648]), .rdlo_in(a4_wr[712]),  .coef_in(coef[128]), .rdup_out(a5_wr[648]), .rdlo_out(a5_wr[712]));
			radix2 #(.width(width)) rd_st4_649  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[649]), .rdlo_in(a4_wr[713]),  .coef_in(coef[144]), .rdup_out(a5_wr[649]), .rdlo_out(a5_wr[713]));
			radix2 #(.width(width)) rd_st4_650  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[650]), .rdlo_in(a4_wr[714]),  .coef_in(coef[160]), .rdup_out(a5_wr[650]), .rdlo_out(a5_wr[714]));
			radix2 #(.width(width)) rd_st4_651  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[651]), .rdlo_in(a4_wr[715]),  .coef_in(coef[176]), .rdup_out(a5_wr[651]), .rdlo_out(a5_wr[715]));
			radix2 #(.width(width)) rd_st4_652  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[652]), .rdlo_in(a4_wr[716]),  .coef_in(coef[192]), .rdup_out(a5_wr[652]), .rdlo_out(a5_wr[716]));
			radix2 #(.width(width)) rd_st4_653  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[653]), .rdlo_in(a4_wr[717]),  .coef_in(coef[208]), .rdup_out(a5_wr[653]), .rdlo_out(a5_wr[717]));
			radix2 #(.width(width)) rd_st4_654  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[654]), .rdlo_in(a4_wr[718]),  .coef_in(coef[224]), .rdup_out(a5_wr[654]), .rdlo_out(a5_wr[718]));
			radix2 #(.width(width)) rd_st4_655  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[655]), .rdlo_in(a4_wr[719]),  .coef_in(coef[240]), .rdup_out(a5_wr[655]), .rdlo_out(a5_wr[719]));
			radix2 #(.width(width)) rd_st4_656  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[656]), .rdlo_in(a4_wr[720]),  .coef_in(coef[256]), .rdup_out(a5_wr[656]), .rdlo_out(a5_wr[720]));
			radix2 #(.width(width)) rd_st4_657  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[657]), .rdlo_in(a4_wr[721]),  .coef_in(coef[272]), .rdup_out(a5_wr[657]), .rdlo_out(a5_wr[721]));
			radix2 #(.width(width)) rd_st4_658  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[658]), .rdlo_in(a4_wr[722]),  .coef_in(coef[288]), .rdup_out(a5_wr[658]), .rdlo_out(a5_wr[722]));
			radix2 #(.width(width)) rd_st4_659  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[659]), .rdlo_in(a4_wr[723]),  .coef_in(coef[304]), .rdup_out(a5_wr[659]), .rdlo_out(a5_wr[723]));
			radix2 #(.width(width)) rd_st4_660  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[660]), .rdlo_in(a4_wr[724]),  .coef_in(coef[320]), .rdup_out(a5_wr[660]), .rdlo_out(a5_wr[724]));
			radix2 #(.width(width)) rd_st4_661  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[661]), .rdlo_in(a4_wr[725]),  .coef_in(coef[336]), .rdup_out(a5_wr[661]), .rdlo_out(a5_wr[725]));
			radix2 #(.width(width)) rd_st4_662  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[662]), .rdlo_in(a4_wr[726]),  .coef_in(coef[352]), .rdup_out(a5_wr[662]), .rdlo_out(a5_wr[726]));
			radix2 #(.width(width)) rd_st4_663  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[663]), .rdlo_in(a4_wr[727]),  .coef_in(coef[368]), .rdup_out(a5_wr[663]), .rdlo_out(a5_wr[727]));
			radix2 #(.width(width)) rd_st4_664  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[664]), .rdlo_in(a4_wr[728]),  .coef_in(coef[384]), .rdup_out(a5_wr[664]), .rdlo_out(a5_wr[728]));
			radix2 #(.width(width)) rd_st4_665  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[665]), .rdlo_in(a4_wr[729]),  .coef_in(coef[400]), .rdup_out(a5_wr[665]), .rdlo_out(a5_wr[729]));
			radix2 #(.width(width)) rd_st4_666  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[666]), .rdlo_in(a4_wr[730]),  .coef_in(coef[416]), .rdup_out(a5_wr[666]), .rdlo_out(a5_wr[730]));
			radix2 #(.width(width)) rd_st4_667  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[667]), .rdlo_in(a4_wr[731]),  .coef_in(coef[432]), .rdup_out(a5_wr[667]), .rdlo_out(a5_wr[731]));
			radix2 #(.width(width)) rd_st4_668  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[668]), .rdlo_in(a4_wr[732]),  .coef_in(coef[448]), .rdup_out(a5_wr[668]), .rdlo_out(a5_wr[732]));
			radix2 #(.width(width)) rd_st4_669  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[669]), .rdlo_in(a4_wr[733]),  .coef_in(coef[464]), .rdup_out(a5_wr[669]), .rdlo_out(a5_wr[733]));
			radix2 #(.width(width)) rd_st4_670  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[670]), .rdlo_in(a4_wr[734]),  .coef_in(coef[480]), .rdup_out(a5_wr[670]), .rdlo_out(a5_wr[734]));
			radix2 #(.width(width)) rd_st4_671  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[671]), .rdlo_in(a4_wr[735]),  .coef_in(coef[496]), .rdup_out(a5_wr[671]), .rdlo_out(a5_wr[735]));
			radix2 #(.width(width)) rd_st4_672  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[672]), .rdlo_in(a4_wr[736]),  .coef_in(coef[512]), .rdup_out(a5_wr[672]), .rdlo_out(a5_wr[736]));
			radix2 #(.width(width)) rd_st4_673  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[673]), .rdlo_in(a4_wr[737]),  .coef_in(coef[528]), .rdup_out(a5_wr[673]), .rdlo_out(a5_wr[737]));
			radix2 #(.width(width)) rd_st4_674  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[674]), .rdlo_in(a4_wr[738]),  .coef_in(coef[544]), .rdup_out(a5_wr[674]), .rdlo_out(a5_wr[738]));
			radix2 #(.width(width)) rd_st4_675  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[675]), .rdlo_in(a4_wr[739]),  .coef_in(coef[560]), .rdup_out(a5_wr[675]), .rdlo_out(a5_wr[739]));
			radix2 #(.width(width)) rd_st4_676  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[676]), .rdlo_in(a4_wr[740]),  .coef_in(coef[576]), .rdup_out(a5_wr[676]), .rdlo_out(a5_wr[740]));
			radix2 #(.width(width)) rd_st4_677  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[677]), .rdlo_in(a4_wr[741]),  .coef_in(coef[592]), .rdup_out(a5_wr[677]), .rdlo_out(a5_wr[741]));
			radix2 #(.width(width)) rd_st4_678  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[678]), .rdlo_in(a4_wr[742]),  .coef_in(coef[608]), .rdup_out(a5_wr[678]), .rdlo_out(a5_wr[742]));
			radix2 #(.width(width)) rd_st4_679  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[679]), .rdlo_in(a4_wr[743]),  .coef_in(coef[624]), .rdup_out(a5_wr[679]), .rdlo_out(a5_wr[743]));
			radix2 #(.width(width)) rd_st4_680  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[680]), .rdlo_in(a4_wr[744]),  .coef_in(coef[640]), .rdup_out(a5_wr[680]), .rdlo_out(a5_wr[744]));
			radix2 #(.width(width)) rd_st4_681  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[681]), .rdlo_in(a4_wr[745]),  .coef_in(coef[656]), .rdup_out(a5_wr[681]), .rdlo_out(a5_wr[745]));
			radix2 #(.width(width)) rd_st4_682  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[682]), .rdlo_in(a4_wr[746]),  .coef_in(coef[672]), .rdup_out(a5_wr[682]), .rdlo_out(a5_wr[746]));
			radix2 #(.width(width)) rd_st4_683  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[683]), .rdlo_in(a4_wr[747]),  .coef_in(coef[688]), .rdup_out(a5_wr[683]), .rdlo_out(a5_wr[747]));
			radix2 #(.width(width)) rd_st4_684  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[684]), .rdlo_in(a4_wr[748]),  .coef_in(coef[704]), .rdup_out(a5_wr[684]), .rdlo_out(a5_wr[748]));
			radix2 #(.width(width)) rd_st4_685  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[685]), .rdlo_in(a4_wr[749]),  .coef_in(coef[720]), .rdup_out(a5_wr[685]), .rdlo_out(a5_wr[749]));
			radix2 #(.width(width)) rd_st4_686  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[686]), .rdlo_in(a4_wr[750]),  .coef_in(coef[736]), .rdup_out(a5_wr[686]), .rdlo_out(a5_wr[750]));
			radix2 #(.width(width)) rd_st4_687  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[687]), .rdlo_in(a4_wr[751]),  .coef_in(coef[752]), .rdup_out(a5_wr[687]), .rdlo_out(a5_wr[751]));
			radix2 #(.width(width)) rd_st4_688  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[688]), .rdlo_in(a4_wr[752]),  .coef_in(coef[768]), .rdup_out(a5_wr[688]), .rdlo_out(a5_wr[752]));
			radix2 #(.width(width)) rd_st4_689  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[689]), .rdlo_in(a4_wr[753]),  .coef_in(coef[784]), .rdup_out(a5_wr[689]), .rdlo_out(a5_wr[753]));
			radix2 #(.width(width)) rd_st4_690  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[690]), .rdlo_in(a4_wr[754]),  .coef_in(coef[800]), .rdup_out(a5_wr[690]), .rdlo_out(a5_wr[754]));
			radix2 #(.width(width)) rd_st4_691  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[691]), .rdlo_in(a4_wr[755]),  .coef_in(coef[816]), .rdup_out(a5_wr[691]), .rdlo_out(a5_wr[755]));
			radix2 #(.width(width)) rd_st4_692  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[692]), .rdlo_in(a4_wr[756]),  .coef_in(coef[832]), .rdup_out(a5_wr[692]), .rdlo_out(a5_wr[756]));
			radix2 #(.width(width)) rd_st4_693  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[693]), .rdlo_in(a4_wr[757]),  .coef_in(coef[848]), .rdup_out(a5_wr[693]), .rdlo_out(a5_wr[757]));
			radix2 #(.width(width)) rd_st4_694  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[694]), .rdlo_in(a4_wr[758]),  .coef_in(coef[864]), .rdup_out(a5_wr[694]), .rdlo_out(a5_wr[758]));
			radix2 #(.width(width)) rd_st4_695  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[695]), .rdlo_in(a4_wr[759]),  .coef_in(coef[880]), .rdup_out(a5_wr[695]), .rdlo_out(a5_wr[759]));
			radix2 #(.width(width)) rd_st4_696  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[696]), .rdlo_in(a4_wr[760]),  .coef_in(coef[896]), .rdup_out(a5_wr[696]), .rdlo_out(a5_wr[760]));
			radix2 #(.width(width)) rd_st4_697  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[697]), .rdlo_in(a4_wr[761]),  .coef_in(coef[912]), .rdup_out(a5_wr[697]), .rdlo_out(a5_wr[761]));
			radix2 #(.width(width)) rd_st4_698  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[698]), .rdlo_in(a4_wr[762]),  .coef_in(coef[928]), .rdup_out(a5_wr[698]), .rdlo_out(a5_wr[762]));
			radix2 #(.width(width)) rd_st4_699  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[699]), .rdlo_in(a4_wr[763]),  .coef_in(coef[944]), .rdup_out(a5_wr[699]), .rdlo_out(a5_wr[763]));
			radix2 #(.width(width)) rd_st4_700  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[700]), .rdlo_in(a4_wr[764]),  .coef_in(coef[960]), .rdup_out(a5_wr[700]), .rdlo_out(a5_wr[764]));
			radix2 #(.width(width)) rd_st4_701  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[701]), .rdlo_in(a4_wr[765]),  .coef_in(coef[976]), .rdup_out(a5_wr[701]), .rdlo_out(a5_wr[765]));
			radix2 #(.width(width)) rd_st4_702  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[702]), .rdlo_in(a4_wr[766]),  .coef_in(coef[992]), .rdup_out(a5_wr[702]), .rdlo_out(a5_wr[766]));
			radix2 #(.width(width)) rd_st4_703  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[703]), .rdlo_in(a4_wr[767]),  .coef_in(coef[1008]), .rdup_out(a5_wr[703]), .rdlo_out(a5_wr[767]));
			radix2 #(.width(width)) rd_st4_768  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[768]), .rdlo_in(a4_wr[832]),  .coef_in(coef[0]), .rdup_out(a5_wr[768]), .rdlo_out(a5_wr[832]));
			radix2 #(.width(width)) rd_st4_769  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[769]), .rdlo_in(a4_wr[833]),  .coef_in(coef[16]), .rdup_out(a5_wr[769]), .rdlo_out(a5_wr[833]));
			radix2 #(.width(width)) rd_st4_770  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[770]), .rdlo_in(a4_wr[834]),  .coef_in(coef[32]), .rdup_out(a5_wr[770]), .rdlo_out(a5_wr[834]));
			radix2 #(.width(width)) rd_st4_771  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[771]), .rdlo_in(a4_wr[835]),  .coef_in(coef[48]), .rdup_out(a5_wr[771]), .rdlo_out(a5_wr[835]));
			radix2 #(.width(width)) rd_st4_772  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[772]), .rdlo_in(a4_wr[836]),  .coef_in(coef[64]), .rdup_out(a5_wr[772]), .rdlo_out(a5_wr[836]));
			radix2 #(.width(width)) rd_st4_773  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[773]), .rdlo_in(a4_wr[837]),  .coef_in(coef[80]), .rdup_out(a5_wr[773]), .rdlo_out(a5_wr[837]));
			radix2 #(.width(width)) rd_st4_774  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[774]), .rdlo_in(a4_wr[838]),  .coef_in(coef[96]), .rdup_out(a5_wr[774]), .rdlo_out(a5_wr[838]));
			radix2 #(.width(width)) rd_st4_775  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[775]), .rdlo_in(a4_wr[839]),  .coef_in(coef[112]), .rdup_out(a5_wr[775]), .rdlo_out(a5_wr[839]));
			radix2 #(.width(width)) rd_st4_776  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[776]), .rdlo_in(a4_wr[840]),  .coef_in(coef[128]), .rdup_out(a5_wr[776]), .rdlo_out(a5_wr[840]));
			radix2 #(.width(width)) rd_st4_777  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[777]), .rdlo_in(a4_wr[841]),  .coef_in(coef[144]), .rdup_out(a5_wr[777]), .rdlo_out(a5_wr[841]));
			radix2 #(.width(width)) rd_st4_778  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[778]), .rdlo_in(a4_wr[842]),  .coef_in(coef[160]), .rdup_out(a5_wr[778]), .rdlo_out(a5_wr[842]));
			radix2 #(.width(width)) rd_st4_779  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[779]), .rdlo_in(a4_wr[843]),  .coef_in(coef[176]), .rdup_out(a5_wr[779]), .rdlo_out(a5_wr[843]));
			radix2 #(.width(width)) rd_st4_780  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[780]), .rdlo_in(a4_wr[844]),  .coef_in(coef[192]), .rdup_out(a5_wr[780]), .rdlo_out(a5_wr[844]));
			radix2 #(.width(width)) rd_st4_781  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[781]), .rdlo_in(a4_wr[845]),  .coef_in(coef[208]), .rdup_out(a5_wr[781]), .rdlo_out(a5_wr[845]));
			radix2 #(.width(width)) rd_st4_782  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[782]), .rdlo_in(a4_wr[846]),  .coef_in(coef[224]), .rdup_out(a5_wr[782]), .rdlo_out(a5_wr[846]));
			radix2 #(.width(width)) rd_st4_783  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[783]), .rdlo_in(a4_wr[847]),  .coef_in(coef[240]), .rdup_out(a5_wr[783]), .rdlo_out(a5_wr[847]));
			radix2 #(.width(width)) rd_st4_784  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[784]), .rdlo_in(a4_wr[848]),  .coef_in(coef[256]), .rdup_out(a5_wr[784]), .rdlo_out(a5_wr[848]));
			radix2 #(.width(width)) rd_st4_785  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[785]), .rdlo_in(a4_wr[849]),  .coef_in(coef[272]), .rdup_out(a5_wr[785]), .rdlo_out(a5_wr[849]));
			radix2 #(.width(width)) rd_st4_786  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[786]), .rdlo_in(a4_wr[850]),  .coef_in(coef[288]), .rdup_out(a5_wr[786]), .rdlo_out(a5_wr[850]));
			radix2 #(.width(width)) rd_st4_787  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[787]), .rdlo_in(a4_wr[851]),  .coef_in(coef[304]), .rdup_out(a5_wr[787]), .rdlo_out(a5_wr[851]));
			radix2 #(.width(width)) rd_st4_788  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[788]), .rdlo_in(a4_wr[852]),  .coef_in(coef[320]), .rdup_out(a5_wr[788]), .rdlo_out(a5_wr[852]));
			radix2 #(.width(width)) rd_st4_789  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[789]), .rdlo_in(a4_wr[853]),  .coef_in(coef[336]), .rdup_out(a5_wr[789]), .rdlo_out(a5_wr[853]));
			radix2 #(.width(width)) rd_st4_790  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[790]), .rdlo_in(a4_wr[854]),  .coef_in(coef[352]), .rdup_out(a5_wr[790]), .rdlo_out(a5_wr[854]));
			radix2 #(.width(width)) rd_st4_791  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[791]), .rdlo_in(a4_wr[855]),  .coef_in(coef[368]), .rdup_out(a5_wr[791]), .rdlo_out(a5_wr[855]));
			radix2 #(.width(width)) rd_st4_792  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[792]), .rdlo_in(a4_wr[856]),  .coef_in(coef[384]), .rdup_out(a5_wr[792]), .rdlo_out(a5_wr[856]));
			radix2 #(.width(width)) rd_st4_793  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[793]), .rdlo_in(a4_wr[857]),  .coef_in(coef[400]), .rdup_out(a5_wr[793]), .rdlo_out(a5_wr[857]));
			radix2 #(.width(width)) rd_st4_794  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[794]), .rdlo_in(a4_wr[858]),  .coef_in(coef[416]), .rdup_out(a5_wr[794]), .rdlo_out(a5_wr[858]));
			radix2 #(.width(width)) rd_st4_795  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[795]), .rdlo_in(a4_wr[859]),  .coef_in(coef[432]), .rdup_out(a5_wr[795]), .rdlo_out(a5_wr[859]));
			radix2 #(.width(width)) rd_st4_796  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[796]), .rdlo_in(a4_wr[860]),  .coef_in(coef[448]), .rdup_out(a5_wr[796]), .rdlo_out(a5_wr[860]));
			radix2 #(.width(width)) rd_st4_797  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[797]), .rdlo_in(a4_wr[861]),  .coef_in(coef[464]), .rdup_out(a5_wr[797]), .rdlo_out(a5_wr[861]));
			radix2 #(.width(width)) rd_st4_798  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[798]), .rdlo_in(a4_wr[862]),  .coef_in(coef[480]), .rdup_out(a5_wr[798]), .rdlo_out(a5_wr[862]));
			radix2 #(.width(width)) rd_st4_799  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[799]), .rdlo_in(a4_wr[863]),  .coef_in(coef[496]), .rdup_out(a5_wr[799]), .rdlo_out(a5_wr[863]));
			radix2 #(.width(width)) rd_st4_800  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[800]), .rdlo_in(a4_wr[864]),  .coef_in(coef[512]), .rdup_out(a5_wr[800]), .rdlo_out(a5_wr[864]));
			radix2 #(.width(width)) rd_st4_801  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[801]), .rdlo_in(a4_wr[865]),  .coef_in(coef[528]), .rdup_out(a5_wr[801]), .rdlo_out(a5_wr[865]));
			radix2 #(.width(width)) rd_st4_802  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[802]), .rdlo_in(a4_wr[866]),  .coef_in(coef[544]), .rdup_out(a5_wr[802]), .rdlo_out(a5_wr[866]));
			radix2 #(.width(width)) rd_st4_803  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[803]), .rdlo_in(a4_wr[867]),  .coef_in(coef[560]), .rdup_out(a5_wr[803]), .rdlo_out(a5_wr[867]));
			radix2 #(.width(width)) rd_st4_804  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[804]), .rdlo_in(a4_wr[868]),  .coef_in(coef[576]), .rdup_out(a5_wr[804]), .rdlo_out(a5_wr[868]));
			radix2 #(.width(width)) rd_st4_805  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[805]), .rdlo_in(a4_wr[869]),  .coef_in(coef[592]), .rdup_out(a5_wr[805]), .rdlo_out(a5_wr[869]));
			radix2 #(.width(width)) rd_st4_806  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[806]), .rdlo_in(a4_wr[870]),  .coef_in(coef[608]), .rdup_out(a5_wr[806]), .rdlo_out(a5_wr[870]));
			radix2 #(.width(width)) rd_st4_807  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[807]), .rdlo_in(a4_wr[871]),  .coef_in(coef[624]), .rdup_out(a5_wr[807]), .rdlo_out(a5_wr[871]));
			radix2 #(.width(width)) rd_st4_808  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[808]), .rdlo_in(a4_wr[872]),  .coef_in(coef[640]), .rdup_out(a5_wr[808]), .rdlo_out(a5_wr[872]));
			radix2 #(.width(width)) rd_st4_809  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[809]), .rdlo_in(a4_wr[873]),  .coef_in(coef[656]), .rdup_out(a5_wr[809]), .rdlo_out(a5_wr[873]));
			radix2 #(.width(width)) rd_st4_810  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[810]), .rdlo_in(a4_wr[874]),  .coef_in(coef[672]), .rdup_out(a5_wr[810]), .rdlo_out(a5_wr[874]));
			radix2 #(.width(width)) rd_st4_811  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[811]), .rdlo_in(a4_wr[875]),  .coef_in(coef[688]), .rdup_out(a5_wr[811]), .rdlo_out(a5_wr[875]));
			radix2 #(.width(width)) rd_st4_812  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[812]), .rdlo_in(a4_wr[876]),  .coef_in(coef[704]), .rdup_out(a5_wr[812]), .rdlo_out(a5_wr[876]));
			radix2 #(.width(width)) rd_st4_813  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[813]), .rdlo_in(a4_wr[877]),  .coef_in(coef[720]), .rdup_out(a5_wr[813]), .rdlo_out(a5_wr[877]));
			radix2 #(.width(width)) rd_st4_814  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[814]), .rdlo_in(a4_wr[878]),  .coef_in(coef[736]), .rdup_out(a5_wr[814]), .rdlo_out(a5_wr[878]));
			radix2 #(.width(width)) rd_st4_815  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[815]), .rdlo_in(a4_wr[879]),  .coef_in(coef[752]), .rdup_out(a5_wr[815]), .rdlo_out(a5_wr[879]));
			radix2 #(.width(width)) rd_st4_816  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[816]), .rdlo_in(a4_wr[880]),  .coef_in(coef[768]), .rdup_out(a5_wr[816]), .rdlo_out(a5_wr[880]));
			radix2 #(.width(width)) rd_st4_817  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[817]), .rdlo_in(a4_wr[881]),  .coef_in(coef[784]), .rdup_out(a5_wr[817]), .rdlo_out(a5_wr[881]));
			radix2 #(.width(width)) rd_st4_818  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[818]), .rdlo_in(a4_wr[882]),  .coef_in(coef[800]), .rdup_out(a5_wr[818]), .rdlo_out(a5_wr[882]));
			radix2 #(.width(width)) rd_st4_819  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[819]), .rdlo_in(a4_wr[883]),  .coef_in(coef[816]), .rdup_out(a5_wr[819]), .rdlo_out(a5_wr[883]));
			radix2 #(.width(width)) rd_st4_820  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[820]), .rdlo_in(a4_wr[884]),  .coef_in(coef[832]), .rdup_out(a5_wr[820]), .rdlo_out(a5_wr[884]));
			radix2 #(.width(width)) rd_st4_821  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[821]), .rdlo_in(a4_wr[885]),  .coef_in(coef[848]), .rdup_out(a5_wr[821]), .rdlo_out(a5_wr[885]));
			radix2 #(.width(width)) rd_st4_822  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[822]), .rdlo_in(a4_wr[886]),  .coef_in(coef[864]), .rdup_out(a5_wr[822]), .rdlo_out(a5_wr[886]));
			radix2 #(.width(width)) rd_st4_823  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[823]), .rdlo_in(a4_wr[887]),  .coef_in(coef[880]), .rdup_out(a5_wr[823]), .rdlo_out(a5_wr[887]));
			radix2 #(.width(width)) rd_st4_824  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[824]), .rdlo_in(a4_wr[888]),  .coef_in(coef[896]), .rdup_out(a5_wr[824]), .rdlo_out(a5_wr[888]));
			radix2 #(.width(width)) rd_st4_825  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[825]), .rdlo_in(a4_wr[889]),  .coef_in(coef[912]), .rdup_out(a5_wr[825]), .rdlo_out(a5_wr[889]));
			radix2 #(.width(width)) rd_st4_826  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[826]), .rdlo_in(a4_wr[890]),  .coef_in(coef[928]), .rdup_out(a5_wr[826]), .rdlo_out(a5_wr[890]));
			radix2 #(.width(width)) rd_st4_827  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[827]), .rdlo_in(a4_wr[891]),  .coef_in(coef[944]), .rdup_out(a5_wr[827]), .rdlo_out(a5_wr[891]));
			radix2 #(.width(width)) rd_st4_828  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[828]), .rdlo_in(a4_wr[892]),  .coef_in(coef[960]), .rdup_out(a5_wr[828]), .rdlo_out(a5_wr[892]));
			radix2 #(.width(width)) rd_st4_829  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[829]), .rdlo_in(a4_wr[893]),  .coef_in(coef[976]), .rdup_out(a5_wr[829]), .rdlo_out(a5_wr[893]));
			radix2 #(.width(width)) rd_st4_830  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[830]), .rdlo_in(a4_wr[894]),  .coef_in(coef[992]), .rdup_out(a5_wr[830]), .rdlo_out(a5_wr[894]));
			radix2 #(.width(width)) rd_st4_831  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[831]), .rdlo_in(a4_wr[895]),  .coef_in(coef[1008]), .rdup_out(a5_wr[831]), .rdlo_out(a5_wr[895]));
			radix2 #(.width(width)) rd_st4_896  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[896]), .rdlo_in(a4_wr[960]),  .coef_in(coef[0]), .rdup_out(a5_wr[896]), .rdlo_out(a5_wr[960]));
			radix2 #(.width(width)) rd_st4_897  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[897]), .rdlo_in(a4_wr[961]),  .coef_in(coef[16]), .rdup_out(a5_wr[897]), .rdlo_out(a5_wr[961]));
			radix2 #(.width(width)) rd_st4_898  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[898]), .rdlo_in(a4_wr[962]),  .coef_in(coef[32]), .rdup_out(a5_wr[898]), .rdlo_out(a5_wr[962]));
			radix2 #(.width(width)) rd_st4_899  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[899]), .rdlo_in(a4_wr[963]),  .coef_in(coef[48]), .rdup_out(a5_wr[899]), .rdlo_out(a5_wr[963]));
			radix2 #(.width(width)) rd_st4_900  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[900]), .rdlo_in(a4_wr[964]),  .coef_in(coef[64]), .rdup_out(a5_wr[900]), .rdlo_out(a5_wr[964]));
			radix2 #(.width(width)) rd_st4_901  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[901]), .rdlo_in(a4_wr[965]),  .coef_in(coef[80]), .rdup_out(a5_wr[901]), .rdlo_out(a5_wr[965]));
			radix2 #(.width(width)) rd_st4_902  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[902]), .rdlo_in(a4_wr[966]),  .coef_in(coef[96]), .rdup_out(a5_wr[902]), .rdlo_out(a5_wr[966]));
			radix2 #(.width(width)) rd_st4_903  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[903]), .rdlo_in(a4_wr[967]),  .coef_in(coef[112]), .rdup_out(a5_wr[903]), .rdlo_out(a5_wr[967]));
			radix2 #(.width(width)) rd_st4_904  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[904]), .rdlo_in(a4_wr[968]),  .coef_in(coef[128]), .rdup_out(a5_wr[904]), .rdlo_out(a5_wr[968]));
			radix2 #(.width(width)) rd_st4_905  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[905]), .rdlo_in(a4_wr[969]),  .coef_in(coef[144]), .rdup_out(a5_wr[905]), .rdlo_out(a5_wr[969]));
			radix2 #(.width(width)) rd_st4_906  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[906]), .rdlo_in(a4_wr[970]),  .coef_in(coef[160]), .rdup_out(a5_wr[906]), .rdlo_out(a5_wr[970]));
			radix2 #(.width(width)) rd_st4_907  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[907]), .rdlo_in(a4_wr[971]),  .coef_in(coef[176]), .rdup_out(a5_wr[907]), .rdlo_out(a5_wr[971]));
			radix2 #(.width(width)) rd_st4_908  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[908]), .rdlo_in(a4_wr[972]),  .coef_in(coef[192]), .rdup_out(a5_wr[908]), .rdlo_out(a5_wr[972]));
			radix2 #(.width(width)) rd_st4_909  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[909]), .rdlo_in(a4_wr[973]),  .coef_in(coef[208]), .rdup_out(a5_wr[909]), .rdlo_out(a5_wr[973]));
			radix2 #(.width(width)) rd_st4_910  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[910]), .rdlo_in(a4_wr[974]),  .coef_in(coef[224]), .rdup_out(a5_wr[910]), .rdlo_out(a5_wr[974]));
			radix2 #(.width(width)) rd_st4_911  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[911]), .rdlo_in(a4_wr[975]),  .coef_in(coef[240]), .rdup_out(a5_wr[911]), .rdlo_out(a5_wr[975]));
			radix2 #(.width(width)) rd_st4_912  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[912]), .rdlo_in(a4_wr[976]),  .coef_in(coef[256]), .rdup_out(a5_wr[912]), .rdlo_out(a5_wr[976]));
			radix2 #(.width(width)) rd_st4_913  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[913]), .rdlo_in(a4_wr[977]),  .coef_in(coef[272]), .rdup_out(a5_wr[913]), .rdlo_out(a5_wr[977]));
			radix2 #(.width(width)) rd_st4_914  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[914]), .rdlo_in(a4_wr[978]),  .coef_in(coef[288]), .rdup_out(a5_wr[914]), .rdlo_out(a5_wr[978]));
			radix2 #(.width(width)) rd_st4_915  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[915]), .rdlo_in(a4_wr[979]),  .coef_in(coef[304]), .rdup_out(a5_wr[915]), .rdlo_out(a5_wr[979]));
			radix2 #(.width(width)) rd_st4_916  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[916]), .rdlo_in(a4_wr[980]),  .coef_in(coef[320]), .rdup_out(a5_wr[916]), .rdlo_out(a5_wr[980]));
			radix2 #(.width(width)) rd_st4_917  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[917]), .rdlo_in(a4_wr[981]),  .coef_in(coef[336]), .rdup_out(a5_wr[917]), .rdlo_out(a5_wr[981]));
			radix2 #(.width(width)) rd_st4_918  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[918]), .rdlo_in(a4_wr[982]),  .coef_in(coef[352]), .rdup_out(a5_wr[918]), .rdlo_out(a5_wr[982]));
			radix2 #(.width(width)) rd_st4_919  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[919]), .rdlo_in(a4_wr[983]),  .coef_in(coef[368]), .rdup_out(a5_wr[919]), .rdlo_out(a5_wr[983]));
			radix2 #(.width(width)) rd_st4_920  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[920]), .rdlo_in(a4_wr[984]),  .coef_in(coef[384]), .rdup_out(a5_wr[920]), .rdlo_out(a5_wr[984]));
			radix2 #(.width(width)) rd_st4_921  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[921]), .rdlo_in(a4_wr[985]),  .coef_in(coef[400]), .rdup_out(a5_wr[921]), .rdlo_out(a5_wr[985]));
			radix2 #(.width(width)) rd_st4_922  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[922]), .rdlo_in(a4_wr[986]),  .coef_in(coef[416]), .rdup_out(a5_wr[922]), .rdlo_out(a5_wr[986]));
			radix2 #(.width(width)) rd_st4_923  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[923]), .rdlo_in(a4_wr[987]),  .coef_in(coef[432]), .rdup_out(a5_wr[923]), .rdlo_out(a5_wr[987]));
			radix2 #(.width(width)) rd_st4_924  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[924]), .rdlo_in(a4_wr[988]),  .coef_in(coef[448]), .rdup_out(a5_wr[924]), .rdlo_out(a5_wr[988]));
			radix2 #(.width(width)) rd_st4_925  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[925]), .rdlo_in(a4_wr[989]),  .coef_in(coef[464]), .rdup_out(a5_wr[925]), .rdlo_out(a5_wr[989]));
			radix2 #(.width(width)) rd_st4_926  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[926]), .rdlo_in(a4_wr[990]),  .coef_in(coef[480]), .rdup_out(a5_wr[926]), .rdlo_out(a5_wr[990]));
			radix2 #(.width(width)) rd_st4_927  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[927]), .rdlo_in(a4_wr[991]),  .coef_in(coef[496]), .rdup_out(a5_wr[927]), .rdlo_out(a5_wr[991]));
			radix2 #(.width(width)) rd_st4_928  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[928]), .rdlo_in(a4_wr[992]),  .coef_in(coef[512]), .rdup_out(a5_wr[928]), .rdlo_out(a5_wr[992]));
			radix2 #(.width(width)) rd_st4_929  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[929]), .rdlo_in(a4_wr[993]),  .coef_in(coef[528]), .rdup_out(a5_wr[929]), .rdlo_out(a5_wr[993]));
			radix2 #(.width(width)) rd_st4_930  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[930]), .rdlo_in(a4_wr[994]),  .coef_in(coef[544]), .rdup_out(a5_wr[930]), .rdlo_out(a5_wr[994]));
			radix2 #(.width(width)) rd_st4_931  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[931]), .rdlo_in(a4_wr[995]),  .coef_in(coef[560]), .rdup_out(a5_wr[931]), .rdlo_out(a5_wr[995]));
			radix2 #(.width(width)) rd_st4_932  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[932]), .rdlo_in(a4_wr[996]),  .coef_in(coef[576]), .rdup_out(a5_wr[932]), .rdlo_out(a5_wr[996]));
			radix2 #(.width(width)) rd_st4_933  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[933]), .rdlo_in(a4_wr[997]),  .coef_in(coef[592]), .rdup_out(a5_wr[933]), .rdlo_out(a5_wr[997]));
			radix2 #(.width(width)) rd_st4_934  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[934]), .rdlo_in(a4_wr[998]),  .coef_in(coef[608]), .rdup_out(a5_wr[934]), .rdlo_out(a5_wr[998]));
			radix2 #(.width(width)) rd_st4_935  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[935]), .rdlo_in(a4_wr[999]),  .coef_in(coef[624]), .rdup_out(a5_wr[935]), .rdlo_out(a5_wr[999]));
			radix2 #(.width(width)) rd_st4_936  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[936]), .rdlo_in(a4_wr[1000]),  .coef_in(coef[640]), .rdup_out(a5_wr[936]), .rdlo_out(a5_wr[1000]));
			radix2 #(.width(width)) rd_st4_937  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[937]), .rdlo_in(a4_wr[1001]),  .coef_in(coef[656]), .rdup_out(a5_wr[937]), .rdlo_out(a5_wr[1001]));
			radix2 #(.width(width)) rd_st4_938  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[938]), .rdlo_in(a4_wr[1002]),  .coef_in(coef[672]), .rdup_out(a5_wr[938]), .rdlo_out(a5_wr[1002]));
			radix2 #(.width(width)) rd_st4_939  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[939]), .rdlo_in(a4_wr[1003]),  .coef_in(coef[688]), .rdup_out(a5_wr[939]), .rdlo_out(a5_wr[1003]));
			radix2 #(.width(width)) rd_st4_940  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[940]), .rdlo_in(a4_wr[1004]),  .coef_in(coef[704]), .rdup_out(a5_wr[940]), .rdlo_out(a5_wr[1004]));
			radix2 #(.width(width)) rd_st4_941  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[941]), .rdlo_in(a4_wr[1005]),  .coef_in(coef[720]), .rdup_out(a5_wr[941]), .rdlo_out(a5_wr[1005]));
			radix2 #(.width(width)) rd_st4_942  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[942]), .rdlo_in(a4_wr[1006]),  .coef_in(coef[736]), .rdup_out(a5_wr[942]), .rdlo_out(a5_wr[1006]));
			radix2 #(.width(width)) rd_st4_943  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[943]), .rdlo_in(a4_wr[1007]),  .coef_in(coef[752]), .rdup_out(a5_wr[943]), .rdlo_out(a5_wr[1007]));
			radix2 #(.width(width)) rd_st4_944  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[944]), .rdlo_in(a4_wr[1008]),  .coef_in(coef[768]), .rdup_out(a5_wr[944]), .rdlo_out(a5_wr[1008]));
			radix2 #(.width(width)) rd_st4_945  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[945]), .rdlo_in(a4_wr[1009]),  .coef_in(coef[784]), .rdup_out(a5_wr[945]), .rdlo_out(a5_wr[1009]));
			radix2 #(.width(width)) rd_st4_946  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[946]), .rdlo_in(a4_wr[1010]),  .coef_in(coef[800]), .rdup_out(a5_wr[946]), .rdlo_out(a5_wr[1010]));
			radix2 #(.width(width)) rd_st4_947  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[947]), .rdlo_in(a4_wr[1011]),  .coef_in(coef[816]), .rdup_out(a5_wr[947]), .rdlo_out(a5_wr[1011]));
			radix2 #(.width(width)) rd_st4_948  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[948]), .rdlo_in(a4_wr[1012]),  .coef_in(coef[832]), .rdup_out(a5_wr[948]), .rdlo_out(a5_wr[1012]));
			radix2 #(.width(width)) rd_st4_949  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[949]), .rdlo_in(a4_wr[1013]),  .coef_in(coef[848]), .rdup_out(a5_wr[949]), .rdlo_out(a5_wr[1013]));
			radix2 #(.width(width)) rd_st4_950  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[950]), .rdlo_in(a4_wr[1014]),  .coef_in(coef[864]), .rdup_out(a5_wr[950]), .rdlo_out(a5_wr[1014]));
			radix2 #(.width(width)) rd_st4_951  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[951]), .rdlo_in(a4_wr[1015]),  .coef_in(coef[880]), .rdup_out(a5_wr[951]), .rdlo_out(a5_wr[1015]));
			radix2 #(.width(width)) rd_st4_952  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[952]), .rdlo_in(a4_wr[1016]),  .coef_in(coef[896]), .rdup_out(a5_wr[952]), .rdlo_out(a5_wr[1016]));
			radix2 #(.width(width)) rd_st4_953  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[953]), .rdlo_in(a4_wr[1017]),  .coef_in(coef[912]), .rdup_out(a5_wr[953]), .rdlo_out(a5_wr[1017]));
			radix2 #(.width(width)) rd_st4_954  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[954]), .rdlo_in(a4_wr[1018]),  .coef_in(coef[928]), .rdup_out(a5_wr[954]), .rdlo_out(a5_wr[1018]));
			radix2 #(.width(width)) rd_st4_955  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[955]), .rdlo_in(a4_wr[1019]),  .coef_in(coef[944]), .rdup_out(a5_wr[955]), .rdlo_out(a5_wr[1019]));
			radix2 #(.width(width)) rd_st4_956  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[956]), .rdlo_in(a4_wr[1020]),  .coef_in(coef[960]), .rdup_out(a5_wr[956]), .rdlo_out(a5_wr[1020]));
			radix2 #(.width(width)) rd_st4_957  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[957]), .rdlo_in(a4_wr[1021]),  .coef_in(coef[976]), .rdup_out(a5_wr[957]), .rdlo_out(a5_wr[1021]));
			radix2 #(.width(width)) rd_st4_958  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[958]), .rdlo_in(a4_wr[1022]),  .coef_in(coef[992]), .rdup_out(a5_wr[958]), .rdlo_out(a5_wr[1022]));
			radix2 #(.width(width)) rd_st4_959  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[959]), .rdlo_in(a4_wr[1023]),  .coef_in(coef[1008]), .rdup_out(a5_wr[959]), .rdlo_out(a5_wr[1023]));
			radix2 #(.width(width)) rd_st4_1024  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1024]), .rdlo_in(a4_wr[1088]),  .coef_in(coef[0]), .rdup_out(a5_wr[1024]), .rdlo_out(a5_wr[1088]));
			radix2 #(.width(width)) rd_st4_1025  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1025]), .rdlo_in(a4_wr[1089]),  .coef_in(coef[16]), .rdup_out(a5_wr[1025]), .rdlo_out(a5_wr[1089]));
			radix2 #(.width(width)) rd_st4_1026  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1026]), .rdlo_in(a4_wr[1090]),  .coef_in(coef[32]), .rdup_out(a5_wr[1026]), .rdlo_out(a5_wr[1090]));
			radix2 #(.width(width)) rd_st4_1027  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1027]), .rdlo_in(a4_wr[1091]),  .coef_in(coef[48]), .rdup_out(a5_wr[1027]), .rdlo_out(a5_wr[1091]));
			radix2 #(.width(width)) rd_st4_1028  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1028]), .rdlo_in(a4_wr[1092]),  .coef_in(coef[64]), .rdup_out(a5_wr[1028]), .rdlo_out(a5_wr[1092]));
			radix2 #(.width(width)) rd_st4_1029  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1029]), .rdlo_in(a4_wr[1093]),  .coef_in(coef[80]), .rdup_out(a5_wr[1029]), .rdlo_out(a5_wr[1093]));
			radix2 #(.width(width)) rd_st4_1030  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1030]), .rdlo_in(a4_wr[1094]),  .coef_in(coef[96]), .rdup_out(a5_wr[1030]), .rdlo_out(a5_wr[1094]));
			radix2 #(.width(width)) rd_st4_1031  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1031]), .rdlo_in(a4_wr[1095]),  .coef_in(coef[112]), .rdup_out(a5_wr[1031]), .rdlo_out(a5_wr[1095]));
			radix2 #(.width(width)) rd_st4_1032  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1032]), .rdlo_in(a4_wr[1096]),  .coef_in(coef[128]), .rdup_out(a5_wr[1032]), .rdlo_out(a5_wr[1096]));
			radix2 #(.width(width)) rd_st4_1033  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1033]), .rdlo_in(a4_wr[1097]),  .coef_in(coef[144]), .rdup_out(a5_wr[1033]), .rdlo_out(a5_wr[1097]));
			radix2 #(.width(width)) rd_st4_1034  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1034]), .rdlo_in(a4_wr[1098]),  .coef_in(coef[160]), .rdup_out(a5_wr[1034]), .rdlo_out(a5_wr[1098]));
			radix2 #(.width(width)) rd_st4_1035  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1035]), .rdlo_in(a4_wr[1099]),  .coef_in(coef[176]), .rdup_out(a5_wr[1035]), .rdlo_out(a5_wr[1099]));
			radix2 #(.width(width)) rd_st4_1036  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1036]), .rdlo_in(a4_wr[1100]),  .coef_in(coef[192]), .rdup_out(a5_wr[1036]), .rdlo_out(a5_wr[1100]));
			radix2 #(.width(width)) rd_st4_1037  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1037]), .rdlo_in(a4_wr[1101]),  .coef_in(coef[208]), .rdup_out(a5_wr[1037]), .rdlo_out(a5_wr[1101]));
			radix2 #(.width(width)) rd_st4_1038  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1038]), .rdlo_in(a4_wr[1102]),  .coef_in(coef[224]), .rdup_out(a5_wr[1038]), .rdlo_out(a5_wr[1102]));
			radix2 #(.width(width)) rd_st4_1039  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1039]), .rdlo_in(a4_wr[1103]),  .coef_in(coef[240]), .rdup_out(a5_wr[1039]), .rdlo_out(a5_wr[1103]));
			radix2 #(.width(width)) rd_st4_1040  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1040]), .rdlo_in(a4_wr[1104]),  .coef_in(coef[256]), .rdup_out(a5_wr[1040]), .rdlo_out(a5_wr[1104]));
			radix2 #(.width(width)) rd_st4_1041  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1041]), .rdlo_in(a4_wr[1105]),  .coef_in(coef[272]), .rdup_out(a5_wr[1041]), .rdlo_out(a5_wr[1105]));
			radix2 #(.width(width)) rd_st4_1042  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1042]), .rdlo_in(a4_wr[1106]),  .coef_in(coef[288]), .rdup_out(a5_wr[1042]), .rdlo_out(a5_wr[1106]));
			radix2 #(.width(width)) rd_st4_1043  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1043]), .rdlo_in(a4_wr[1107]),  .coef_in(coef[304]), .rdup_out(a5_wr[1043]), .rdlo_out(a5_wr[1107]));
			radix2 #(.width(width)) rd_st4_1044  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1044]), .rdlo_in(a4_wr[1108]),  .coef_in(coef[320]), .rdup_out(a5_wr[1044]), .rdlo_out(a5_wr[1108]));
			radix2 #(.width(width)) rd_st4_1045  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1045]), .rdlo_in(a4_wr[1109]),  .coef_in(coef[336]), .rdup_out(a5_wr[1045]), .rdlo_out(a5_wr[1109]));
			radix2 #(.width(width)) rd_st4_1046  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1046]), .rdlo_in(a4_wr[1110]),  .coef_in(coef[352]), .rdup_out(a5_wr[1046]), .rdlo_out(a5_wr[1110]));
			radix2 #(.width(width)) rd_st4_1047  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1047]), .rdlo_in(a4_wr[1111]),  .coef_in(coef[368]), .rdup_out(a5_wr[1047]), .rdlo_out(a5_wr[1111]));
			radix2 #(.width(width)) rd_st4_1048  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1048]), .rdlo_in(a4_wr[1112]),  .coef_in(coef[384]), .rdup_out(a5_wr[1048]), .rdlo_out(a5_wr[1112]));
			radix2 #(.width(width)) rd_st4_1049  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1049]), .rdlo_in(a4_wr[1113]),  .coef_in(coef[400]), .rdup_out(a5_wr[1049]), .rdlo_out(a5_wr[1113]));
			radix2 #(.width(width)) rd_st4_1050  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1050]), .rdlo_in(a4_wr[1114]),  .coef_in(coef[416]), .rdup_out(a5_wr[1050]), .rdlo_out(a5_wr[1114]));
			radix2 #(.width(width)) rd_st4_1051  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1051]), .rdlo_in(a4_wr[1115]),  .coef_in(coef[432]), .rdup_out(a5_wr[1051]), .rdlo_out(a5_wr[1115]));
			radix2 #(.width(width)) rd_st4_1052  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1052]), .rdlo_in(a4_wr[1116]),  .coef_in(coef[448]), .rdup_out(a5_wr[1052]), .rdlo_out(a5_wr[1116]));
			radix2 #(.width(width)) rd_st4_1053  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1053]), .rdlo_in(a4_wr[1117]),  .coef_in(coef[464]), .rdup_out(a5_wr[1053]), .rdlo_out(a5_wr[1117]));
			radix2 #(.width(width)) rd_st4_1054  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1054]), .rdlo_in(a4_wr[1118]),  .coef_in(coef[480]), .rdup_out(a5_wr[1054]), .rdlo_out(a5_wr[1118]));
			radix2 #(.width(width)) rd_st4_1055  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1055]), .rdlo_in(a4_wr[1119]),  .coef_in(coef[496]), .rdup_out(a5_wr[1055]), .rdlo_out(a5_wr[1119]));
			radix2 #(.width(width)) rd_st4_1056  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1056]), .rdlo_in(a4_wr[1120]),  .coef_in(coef[512]), .rdup_out(a5_wr[1056]), .rdlo_out(a5_wr[1120]));
			radix2 #(.width(width)) rd_st4_1057  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1057]), .rdlo_in(a4_wr[1121]),  .coef_in(coef[528]), .rdup_out(a5_wr[1057]), .rdlo_out(a5_wr[1121]));
			radix2 #(.width(width)) rd_st4_1058  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1058]), .rdlo_in(a4_wr[1122]),  .coef_in(coef[544]), .rdup_out(a5_wr[1058]), .rdlo_out(a5_wr[1122]));
			radix2 #(.width(width)) rd_st4_1059  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1059]), .rdlo_in(a4_wr[1123]),  .coef_in(coef[560]), .rdup_out(a5_wr[1059]), .rdlo_out(a5_wr[1123]));
			radix2 #(.width(width)) rd_st4_1060  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1060]), .rdlo_in(a4_wr[1124]),  .coef_in(coef[576]), .rdup_out(a5_wr[1060]), .rdlo_out(a5_wr[1124]));
			radix2 #(.width(width)) rd_st4_1061  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1061]), .rdlo_in(a4_wr[1125]),  .coef_in(coef[592]), .rdup_out(a5_wr[1061]), .rdlo_out(a5_wr[1125]));
			radix2 #(.width(width)) rd_st4_1062  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1062]), .rdlo_in(a4_wr[1126]),  .coef_in(coef[608]), .rdup_out(a5_wr[1062]), .rdlo_out(a5_wr[1126]));
			radix2 #(.width(width)) rd_st4_1063  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1063]), .rdlo_in(a4_wr[1127]),  .coef_in(coef[624]), .rdup_out(a5_wr[1063]), .rdlo_out(a5_wr[1127]));
			radix2 #(.width(width)) rd_st4_1064  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1064]), .rdlo_in(a4_wr[1128]),  .coef_in(coef[640]), .rdup_out(a5_wr[1064]), .rdlo_out(a5_wr[1128]));
			radix2 #(.width(width)) rd_st4_1065  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1065]), .rdlo_in(a4_wr[1129]),  .coef_in(coef[656]), .rdup_out(a5_wr[1065]), .rdlo_out(a5_wr[1129]));
			radix2 #(.width(width)) rd_st4_1066  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1066]), .rdlo_in(a4_wr[1130]),  .coef_in(coef[672]), .rdup_out(a5_wr[1066]), .rdlo_out(a5_wr[1130]));
			radix2 #(.width(width)) rd_st4_1067  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1067]), .rdlo_in(a4_wr[1131]),  .coef_in(coef[688]), .rdup_out(a5_wr[1067]), .rdlo_out(a5_wr[1131]));
			radix2 #(.width(width)) rd_st4_1068  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1068]), .rdlo_in(a4_wr[1132]),  .coef_in(coef[704]), .rdup_out(a5_wr[1068]), .rdlo_out(a5_wr[1132]));
			radix2 #(.width(width)) rd_st4_1069  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1069]), .rdlo_in(a4_wr[1133]),  .coef_in(coef[720]), .rdup_out(a5_wr[1069]), .rdlo_out(a5_wr[1133]));
			radix2 #(.width(width)) rd_st4_1070  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1070]), .rdlo_in(a4_wr[1134]),  .coef_in(coef[736]), .rdup_out(a5_wr[1070]), .rdlo_out(a5_wr[1134]));
			radix2 #(.width(width)) rd_st4_1071  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1071]), .rdlo_in(a4_wr[1135]),  .coef_in(coef[752]), .rdup_out(a5_wr[1071]), .rdlo_out(a5_wr[1135]));
			radix2 #(.width(width)) rd_st4_1072  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1072]), .rdlo_in(a4_wr[1136]),  .coef_in(coef[768]), .rdup_out(a5_wr[1072]), .rdlo_out(a5_wr[1136]));
			radix2 #(.width(width)) rd_st4_1073  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1073]), .rdlo_in(a4_wr[1137]),  .coef_in(coef[784]), .rdup_out(a5_wr[1073]), .rdlo_out(a5_wr[1137]));
			radix2 #(.width(width)) rd_st4_1074  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1074]), .rdlo_in(a4_wr[1138]),  .coef_in(coef[800]), .rdup_out(a5_wr[1074]), .rdlo_out(a5_wr[1138]));
			radix2 #(.width(width)) rd_st4_1075  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1075]), .rdlo_in(a4_wr[1139]),  .coef_in(coef[816]), .rdup_out(a5_wr[1075]), .rdlo_out(a5_wr[1139]));
			radix2 #(.width(width)) rd_st4_1076  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1076]), .rdlo_in(a4_wr[1140]),  .coef_in(coef[832]), .rdup_out(a5_wr[1076]), .rdlo_out(a5_wr[1140]));
			radix2 #(.width(width)) rd_st4_1077  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1077]), .rdlo_in(a4_wr[1141]),  .coef_in(coef[848]), .rdup_out(a5_wr[1077]), .rdlo_out(a5_wr[1141]));
			radix2 #(.width(width)) rd_st4_1078  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1078]), .rdlo_in(a4_wr[1142]),  .coef_in(coef[864]), .rdup_out(a5_wr[1078]), .rdlo_out(a5_wr[1142]));
			radix2 #(.width(width)) rd_st4_1079  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1079]), .rdlo_in(a4_wr[1143]),  .coef_in(coef[880]), .rdup_out(a5_wr[1079]), .rdlo_out(a5_wr[1143]));
			radix2 #(.width(width)) rd_st4_1080  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1080]), .rdlo_in(a4_wr[1144]),  .coef_in(coef[896]), .rdup_out(a5_wr[1080]), .rdlo_out(a5_wr[1144]));
			radix2 #(.width(width)) rd_st4_1081  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1081]), .rdlo_in(a4_wr[1145]),  .coef_in(coef[912]), .rdup_out(a5_wr[1081]), .rdlo_out(a5_wr[1145]));
			radix2 #(.width(width)) rd_st4_1082  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1082]), .rdlo_in(a4_wr[1146]),  .coef_in(coef[928]), .rdup_out(a5_wr[1082]), .rdlo_out(a5_wr[1146]));
			radix2 #(.width(width)) rd_st4_1083  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1083]), .rdlo_in(a4_wr[1147]),  .coef_in(coef[944]), .rdup_out(a5_wr[1083]), .rdlo_out(a5_wr[1147]));
			radix2 #(.width(width)) rd_st4_1084  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1084]), .rdlo_in(a4_wr[1148]),  .coef_in(coef[960]), .rdup_out(a5_wr[1084]), .rdlo_out(a5_wr[1148]));
			radix2 #(.width(width)) rd_st4_1085  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1085]), .rdlo_in(a4_wr[1149]),  .coef_in(coef[976]), .rdup_out(a5_wr[1085]), .rdlo_out(a5_wr[1149]));
			radix2 #(.width(width)) rd_st4_1086  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1086]), .rdlo_in(a4_wr[1150]),  .coef_in(coef[992]), .rdup_out(a5_wr[1086]), .rdlo_out(a5_wr[1150]));
			radix2 #(.width(width)) rd_st4_1087  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1087]), .rdlo_in(a4_wr[1151]),  .coef_in(coef[1008]), .rdup_out(a5_wr[1087]), .rdlo_out(a5_wr[1151]));
			radix2 #(.width(width)) rd_st4_1152  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1152]), .rdlo_in(a4_wr[1216]),  .coef_in(coef[0]), .rdup_out(a5_wr[1152]), .rdlo_out(a5_wr[1216]));
			radix2 #(.width(width)) rd_st4_1153  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1153]), .rdlo_in(a4_wr[1217]),  .coef_in(coef[16]), .rdup_out(a5_wr[1153]), .rdlo_out(a5_wr[1217]));
			radix2 #(.width(width)) rd_st4_1154  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1154]), .rdlo_in(a4_wr[1218]),  .coef_in(coef[32]), .rdup_out(a5_wr[1154]), .rdlo_out(a5_wr[1218]));
			radix2 #(.width(width)) rd_st4_1155  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1155]), .rdlo_in(a4_wr[1219]),  .coef_in(coef[48]), .rdup_out(a5_wr[1155]), .rdlo_out(a5_wr[1219]));
			radix2 #(.width(width)) rd_st4_1156  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1156]), .rdlo_in(a4_wr[1220]),  .coef_in(coef[64]), .rdup_out(a5_wr[1156]), .rdlo_out(a5_wr[1220]));
			radix2 #(.width(width)) rd_st4_1157  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1157]), .rdlo_in(a4_wr[1221]),  .coef_in(coef[80]), .rdup_out(a5_wr[1157]), .rdlo_out(a5_wr[1221]));
			radix2 #(.width(width)) rd_st4_1158  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1158]), .rdlo_in(a4_wr[1222]),  .coef_in(coef[96]), .rdup_out(a5_wr[1158]), .rdlo_out(a5_wr[1222]));
			radix2 #(.width(width)) rd_st4_1159  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1159]), .rdlo_in(a4_wr[1223]),  .coef_in(coef[112]), .rdup_out(a5_wr[1159]), .rdlo_out(a5_wr[1223]));
			radix2 #(.width(width)) rd_st4_1160  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1160]), .rdlo_in(a4_wr[1224]),  .coef_in(coef[128]), .rdup_out(a5_wr[1160]), .rdlo_out(a5_wr[1224]));
			radix2 #(.width(width)) rd_st4_1161  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1161]), .rdlo_in(a4_wr[1225]),  .coef_in(coef[144]), .rdup_out(a5_wr[1161]), .rdlo_out(a5_wr[1225]));
			radix2 #(.width(width)) rd_st4_1162  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1162]), .rdlo_in(a4_wr[1226]),  .coef_in(coef[160]), .rdup_out(a5_wr[1162]), .rdlo_out(a5_wr[1226]));
			radix2 #(.width(width)) rd_st4_1163  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1163]), .rdlo_in(a4_wr[1227]),  .coef_in(coef[176]), .rdup_out(a5_wr[1163]), .rdlo_out(a5_wr[1227]));
			radix2 #(.width(width)) rd_st4_1164  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1164]), .rdlo_in(a4_wr[1228]),  .coef_in(coef[192]), .rdup_out(a5_wr[1164]), .rdlo_out(a5_wr[1228]));
			radix2 #(.width(width)) rd_st4_1165  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1165]), .rdlo_in(a4_wr[1229]),  .coef_in(coef[208]), .rdup_out(a5_wr[1165]), .rdlo_out(a5_wr[1229]));
			radix2 #(.width(width)) rd_st4_1166  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1166]), .rdlo_in(a4_wr[1230]),  .coef_in(coef[224]), .rdup_out(a5_wr[1166]), .rdlo_out(a5_wr[1230]));
			radix2 #(.width(width)) rd_st4_1167  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1167]), .rdlo_in(a4_wr[1231]),  .coef_in(coef[240]), .rdup_out(a5_wr[1167]), .rdlo_out(a5_wr[1231]));
			radix2 #(.width(width)) rd_st4_1168  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1168]), .rdlo_in(a4_wr[1232]),  .coef_in(coef[256]), .rdup_out(a5_wr[1168]), .rdlo_out(a5_wr[1232]));
			radix2 #(.width(width)) rd_st4_1169  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1169]), .rdlo_in(a4_wr[1233]),  .coef_in(coef[272]), .rdup_out(a5_wr[1169]), .rdlo_out(a5_wr[1233]));
			radix2 #(.width(width)) rd_st4_1170  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1170]), .rdlo_in(a4_wr[1234]),  .coef_in(coef[288]), .rdup_out(a5_wr[1170]), .rdlo_out(a5_wr[1234]));
			radix2 #(.width(width)) rd_st4_1171  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1171]), .rdlo_in(a4_wr[1235]),  .coef_in(coef[304]), .rdup_out(a5_wr[1171]), .rdlo_out(a5_wr[1235]));
			radix2 #(.width(width)) rd_st4_1172  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1172]), .rdlo_in(a4_wr[1236]),  .coef_in(coef[320]), .rdup_out(a5_wr[1172]), .rdlo_out(a5_wr[1236]));
			radix2 #(.width(width)) rd_st4_1173  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1173]), .rdlo_in(a4_wr[1237]),  .coef_in(coef[336]), .rdup_out(a5_wr[1173]), .rdlo_out(a5_wr[1237]));
			radix2 #(.width(width)) rd_st4_1174  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1174]), .rdlo_in(a4_wr[1238]),  .coef_in(coef[352]), .rdup_out(a5_wr[1174]), .rdlo_out(a5_wr[1238]));
			radix2 #(.width(width)) rd_st4_1175  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1175]), .rdlo_in(a4_wr[1239]),  .coef_in(coef[368]), .rdup_out(a5_wr[1175]), .rdlo_out(a5_wr[1239]));
			radix2 #(.width(width)) rd_st4_1176  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1176]), .rdlo_in(a4_wr[1240]),  .coef_in(coef[384]), .rdup_out(a5_wr[1176]), .rdlo_out(a5_wr[1240]));
			radix2 #(.width(width)) rd_st4_1177  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1177]), .rdlo_in(a4_wr[1241]),  .coef_in(coef[400]), .rdup_out(a5_wr[1177]), .rdlo_out(a5_wr[1241]));
			radix2 #(.width(width)) rd_st4_1178  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1178]), .rdlo_in(a4_wr[1242]),  .coef_in(coef[416]), .rdup_out(a5_wr[1178]), .rdlo_out(a5_wr[1242]));
			radix2 #(.width(width)) rd_st4_1179  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1179]), .rdlo_in(a4_wr[1243]),  .coef_in(coef[432]), .rdup_out(a5_wr[1179]), .rdlo_out(a5_wr[1243]));
			radix2 #(.width(width)) rd_st4_1180  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1180]), .rdlo_in(a4_wr[1244]),  .coef_in(coef[448]), .rdup_out(a5_wr[1180]), .rdlo_out(a5_wr[1244]));
			radix2 #(.width(width)) rd_st4_1181  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1181]), .rdlo_in(a4_wr[1245]),  .coef_in(coef[464]), .rdup_out(a5_wr[1181]), .rdlo_out(a5_wr[1245]));
			radix2 #(.width(width)) rd_st4_1182  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1182]), .rdlo_in(a4_wr[1246]),  .coef_in(coef[480]), .rdup_out(a5_wr[1182]), .rdlo_out(a5_wr[1246]));
			radix2 #(.width(width)) rd_st4_1183  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1183]), .rdlo_in(a4_wr[1247]),  .coef_in(coef[496]), .rdup_out(a5_wr[1183]), .rdlo_out(a5_wr[1247]));
			radix2 #(.width(width)) rd_st4_1184  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1184]), .rdlo_in(a4_wr[1248]),  .coef_in(coef[512]), .rdup_out(a5_wr[1184]), .rdlo_out(a5_wr[1248]));
			radix2 #(.width(width)) rd_st4_1185  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1185]), .rdlo_in(a4_wr[1249]),  .coef_in(coef[528]), .rdup_out(a5_wr[1185]), .rdlo_out(a5_wr[1249]));
			radix2 #(.width(width)) rd_st4_1186  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1186]), .rdlo_in(a4_wr[1250]),  .coef_in(coef[544]), .rdup_out(a5_wr[1186]), .rdlo_out(a5_wr[1250]));
			radix2 #(.width(width)) rd_st4_1187  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1187]), .rdlo_in(a4_wr[1251]),  .coef_in(coef[560]), .rdup_out(a5_wr[1187]), .rdlo_out(a5_wr[1251]));
			radix2 #(.width(width)) rd_st4_1188  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1188]), .rdlo_in(a4_wr[1252]),  .coef_in(coef[576]), .rdup_out(a5_wr[1188]), .rdlo_out(a5_wr[1252]));
			radix2 #(.width(width)) rd_st4_1189  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1189]), .rdlo_in(a4_wr[1253]),  .coef_in(coef[592]), .rdup_out(a5_wr[1189]), .rdlo_out(a5_wr[1253]));
			radix2 #(.width(width)) rd_st4_1190  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1190]), .rdlo_in(a4_wr[1254]),  .coef_in(coef[608]), .rdup_out(a5_wr[1190]), .rdlo_out(a5_wr[1254]));
			radix2 #(.width(width)) rd_st4_1191  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1191]), .rdlo_in(a4_wr[1255]),  .coef_in(coef[624]), .rdup_out(a5_wr[1191]), .rdlo_out(a5_wr[1255]));
			radix2 #(.width(width)) rd_st4_1192  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1192]), .rdlo_in(a4_wr[1256]),  .coef_in(coef[640]), .rdup_out(a5_wr[1192]), .rdlo_out(a5_wr[1256]));
			radix2 #(.width(width)) rd_st4_1193  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1193]), .rdlo_in(a4_wr[1257]),  .coef_in(coef[656]), .rdup_out(a5_wr[1193]), .rdlo_out(a5_wr[1257]));
			radix2 #(.width(width)) rd_st4_1194  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1194]), .rdlo_in(a4_wr[1258]),  .coef_in(coef[672]), .rdup_out(a5_wr[1194]), .rdlo_out(a5_wr[1258]));
			radix2 #(.width(width)) rd_st4_1195  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1195]), .rdlo_in(a4_wr[1259]),  .coef_in(coef[688]), .rdup_out(a5_wr[1195]), .rdlo_out(a5_wr[1259]));
			radix2 #(.width(width)) rd_st4_1196  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1196]), .rdlo_in(a4_wr[1260]),  .coef_in(coef[704]), .rdup_out(a5_wr[1196]), .rdlo_out(a5_wr[1260]));
			radix2 #(.width(width)) rd_st4_1197  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1197]), .rdlo_in(a4_wr[1261]),  .coef_in(coef[720]), .rdup_out(a5_wr[1197]), .rdlo_out(a5_wr[1261]));
			radix2 #(.width(width)) rd_st4_1198  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1198]), .rdlo_in(a4_wr[1262]),  .coef_in(coef[736]), .rdup_out(a5_wr[1198]), .rdlo_out(a5_wr[1262]));
			radix2 #(.width(width)) rd_st4_1199  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1199]), .rdlo_in(a4_wr[1263]),  .coef_in(coef[752]), .rdup_out(a5_wr[1199]), .rdlo_out(a5_wr[1263]));
			radix2 #(.width(width)) rd_st4_1200  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1200]), .rdlo_in(a4_wr[1264]),  .coef_in(coef[768]), .rdup_out(a5_wr[1200]), .rdlo_out(a5_wr[1264]));
			radix2 #(.width(width)) rd_st4_1201  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1201]), .rdlo_in(a4_wr[1265]),  .coef_in(coef[784]), .rdup_out(a5_wr[1201]), .rdlo_out(a5_wr[1265]));
			radix2 #(.width(width)) rd_st4_1202  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1202]), .rdlo_in(a4_wr[1266]),  .coef_in(coef[800]), .rdup_out(a5_wr[1202]), .rdlo_out(a5_wr[1266]));
			radix2 #(.width(width)) rd_st4_1203  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1203]), .rdlo_in(a4_wr[1267]),  .coef_in(coef[816]), .rdup_out(a5_wr[1203]), .rdlo_out(a5_wr[1267]));
			radix2 #(.width(width)) rd_st4_1204  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1204]), .rdlo_in(a4_wr[1268]),  .coef_in(coef[832]), .rdup_out(a5_wr[1204]), .rdlo_out(a5_wr[1268]));
			radix2 #(.width(width)) rd_st4_1205  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1205]), .rdlo_in(a4_wr[1269]),  .coef_in(coef[848]), .rdup_out(a5_wr[1205]), .rdlo_out(a5_wr[1269]));
			radix2 #(.width(width)) rd_st4_1206  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1206]), .rdlo_in(a4_wr[1270]),  .coef_in(coef[864]), .rdup_out(a5_wr[1206]), .rdlo_out(a5_wr[1270]));
			radix2 #(.width(width)) rd_st4_1207  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1207]), .rdlo_in(a4_wr[1271]),  .coef_in(coef[880]), .rdup_out(a5_wr[1207]), .rdlo_out(a5_wr[1271]));
			radix2 #(.width(width)) rd_st4_1208  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1208]), .rdlo_in(a4_wr[1272]),  .coef_in(coef[896]), .rdup_out(a5_wr[1208]), .rdlo_out(a5_wr[1272]));
			radix2 #(.width(width)) rd_st4_1209  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1209]), .rdlo_in(a4_wr[1273]),  .coef_in(coef[912]), .rdup_out(a5_wr[1209]), .rdlo_out(a5_wr[1273]));
			radix2 #(.width(width)) rd_st4_1210  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1210]), .rdlo_in(a4_wr[1274]),  .coef_in(coef[928]), .rdup_out(a5_wr[1210]), .rdlo_out(a5_wr[1274]));
			radix2 #(.width(width)) rd_st4_1211  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1211]), .rdlo_in(a4_wr[1275]),  .coef_in(coef[944]), .rdup_out(a5_wr[1211]), .rdlo_out(a5_wr[1275]));
			radix2 #(.width(width)) rd_st4_1212  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1212]), .rdlo_in(a4_wr[1276]),  .coef_in(coef[960]), .rdup_out(a5_wr[1212]), .rdlo_out(a5_wr[1276]));
			radix2 #(.width(width)) rd_st4_1213  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1213]), .rdlo_in(a4_wr[1277]),  .coef_in(coef[976]), .rdup_out(a5_wr[1213]), .rdlo_out(a5_wr[1277]));
			radix2 #(.width(width)) rd_st4_1214  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1214]), .rdlo_in(a4_wr[1278]),  .coef_in(coef[992]), .rdup_out(a5_wr[1214]), .rdlo_out(a5_wr[1278]));
			radix2 #(.width(width)) rd_st4_1215  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1215]), .rdlo_in(a4_wr[1279]),  .coef_in(coef[1008]), .rdup_out(a5_wr[1215]), .rdlo_out(a5_wr[1279]));
			radix2 #(.width(width)) rd_st4_1280  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1280]), .rdlo_in(a4_wr[1344]),  .coef_in(coef[0]), .rdup_out(a5_wr[1280]), .rdlo_out(a5_wr[1344]));
			radix2 #(.width(width)) rd_st4_1281  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1281]), .rdlo_in(a4_wr[1345]),  .coef_in(coef[16]), .rdup_out(a5_wr[1281]), .rdlo_out(a5_wr[1345]));
			radix2 #(.width(width)) rd_st4_1282  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1282]), .rdlo_in(a4_wr[1346]),  .coef_in(coef[32]), .rdup_out(a5_wr[1282]), .rdlo_out(a5_wr[1346]));
			radix2 #(.width(width)) rd_st4_1283  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1283]), .rdlo_in(a4_wr[1347]),  .coef_in(coef[48]), .rdup_out(a5_wr[1283]), .rdlo_out(a5_wr[1347]));
			radix2 #(.width(width)) rd_st4_1284  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1284]), .rdlo_in(a4_wr[1348]),  .coef_in(coef[64]), .rdup_out(a5_wr[1284]), .rdlo_out(a5_wr[1348]));
			radix2 #(.width(width)) rd_st4_1285  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1285]), .rdlo_in(a4_wr[1349]),  .coef_in(coef[80]), .rdup_out(a5_wr[1285]), .rdlo_out(a5_wr[1349]));
			radix2 #(.width(width)) rd_st4_1286  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1286]), .rdlo_in(a4_wr[1350]),  .coef_in(coef[96]), .rdup_out(a5_wr[1286]), .rdlo_out(a5_wr[1350]));
			radix2 #(.width(width)) rd_st4_1287  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1287]), .rdlo_in(a4_wr[1351]),  .coef_in(coef[112]), .rdup_out(a5_wr[1287]), .rdlo_out(a5_wr[1351]));
			radix2 #(.width(width)) rd_st4_1288  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1288]), .rdlo_in(a4_wr[1352]),  .coef_in(coef[128]), .rdup_out(a5_wr[1288]), .rdlo_out(a5_wr[1352]));
			radix2 #(.width(width)) rd_st4_1289  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1289]), .rdlo_in(a4_wr[1353]),  .coef_in(coef[144]), .rdup_out(a5_wr[1289]), .rdlo_out(a5_wr[1353]));
			radix2 #(.width(width)) rd_st4_1290  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1290]), .rdlo_in(a4_wr[1354]),  .coef_in(coef[160]), .rdup_out(a5_wr[1290]), .rdlo_out(a5_wr[1354]));
			radix2 #(.width(width)) rd_st4_1291  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1291]), .rdlo_in(a4_wr[1355]),  .coef_in(coef[176]), .rdup_out(a5_wr[1291]), .rdlo_out(a5_wr[1355]));
			radix2 #(.width(width)) rd_st4_1292  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1292]), .rdlo_in(a4_wr[1356]),  .coef_in(coef[192]), .rdup_out(a5_wr[1292]), .rdlo_out(a5_wr[1356]));
			radix2 #(.width(width)) rd_st4_1293  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1293]), .rdlo_in(a4_wr[1357]),  .coef_in(coef[208]), .rdup_out(a5_wr[1293]), .rdlo_out(a5_wr[1357]));
			radix2 #(.width(width)) rd_st4_1294  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1294]), .rdlo_in(a4_wr[1358]),  .coef_in(coef[224]), .rdup_out(a5_wr[1294]), .rdlo_out(a5_wr[1358]));
			radix2 #(.width(width)) rd_st4_1295  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1295]), .rdlo_in(a4_wr[1359]),  .coef_in(coef[240]), .rdup_out(a5_wr[1295]), .rdlo_out(a5_wr[1359]));
			radix2 #(.width(width)) rd_st4_1296  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1296]), .rdlo_in(a4_wr[1360]),  .coef_in(coef[256]), .rdup_out(a5_wr[1296]), .rdlo_out(a5_wr[1360]));
			radix2 #(.width(width)) rd_st4_1297  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1297]), .rdlo_in(a4_wr[1361]),  .coef_in(coef[272]), .rdup_out(a5_wr[1297]), .rdlo_out(a5_wr[1361]));
			radix2 #(.width(width)) rd_st4_1298  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1298]), .rdlo_in(a4_wr[1362]),  .coef_in(coef[288]), .rdup_out(a5_wr[1298]), .rdlo_out(a5_wr[1362]));
			radix2 #(.width(width)) rd_st4_1299  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1299]), .rdlo_in(a4_wr[1363]),  .coef_in(coef[304]), .rdup_out(a5_wr[1299]), .rdlo_out(a5_wr[1363]));
			radix2 #(.width(width)) rd_st4_1300  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1300]), .rdlo_in(a4_wr[1364]),  .coef_in(coef[320]), .rdup_out(a5_wr[1300]), .rdlo_out(a5_wr[1364]));
			radix2 #(.width(width)) rd_st4_1301  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1301]), .rdlo_in(a4_wr[1365]),  .coef_in(coef[336]), .rdup_out(a5_wr[1301]), .rdlo_out(a5_wr[1365]));
			radix2 #(.width(width)) rd_st4_1302  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1302]), .rdlo_in(a4_wr[1366]),  .coef_in(coef[352]), .rdup_out(a5_wr[1302]), .rdlo_out(a5_wr[1366]));
			radix2 #(.width(width)) rd_st4_1303  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1303]), .rdlo_in(a4_wr[1367]),  .coef_in(coef[368]), .rdup_out(a5_wr[1303]), .rdlo_out(a5_wr[1367]));
			radix2 #(.width(width)) rd_st4_1304  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1304]), .rdlo_in(a4_wr[1368]),  .coef_in(coef[384]), .rdup_out(a5_wr[1304]), .rdlo_out(a5_wr[1368]));
			radix2 #(.width(width)) rd_st4_1305  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1305]), .rdlo_in(a4_wr[1369]),  .coef_in(coef[400]), .rdup_out(a5_wr[1305]), .rdlo_out(a5_wr[1369]));
			radix2 #(.width(width)) rd_st4_1306  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1306]), .rdlo_in(a4_wr[1370]),  .coef_in(coef[416]), .rdup_out(a5_wr[1306]), .rdlo_out(a5_wr[1370]));
			radix2 #(.width(width)) rd_st4_1307  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1307]), .rdlo_in(a4_wr[1371]),  .coef_in(coef[432]), .rdup_out(a5_wr[1307]), .rdlo_out(a5_wr[1371]));
			radix2 #(.width(width)) rd_st4_1308  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1308]), .rdlo_in(a4_wr[1372]),  .coef_in(coef[448]), .rdup_out(a5_wr[1308]), .rdlo_out(a5_wr[1372]));
			radix2 #(.width(width)) rd_st4_1309  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1309]), .rdlo_in(a4_wr[1373]),  .coef_in(coef[464]), .rdup_out(a5_wr[1309]), .rdlo_out(a5_wr[1373]));
			radix2 #(.width(width)) rd_st4_1310  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1310]), .rdlo_in(a4_wr[1374]),  .coef_in(coef[480]), .rdup_out(a5_wr[1310]), .rdlo_out(a5_wr[1374]));
			radix2 #(.width(width)) rd_st4_1311  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1311]), .rdlo_in(a4_wr[1375]),  .coef_in(coef[496]), .rdup_out(a5_wr[1311]), .rdlo_out(a5_wr[1375]));
			radix2 #(.width(width)) rd_st4_1312  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1312]), .rdlo_in(a4_wr[1376]),  .coef_in(coef[512]), .rdup_out(a5_wr[1312]), .rdlo_out(a5_wr[1376]));
			radix2 #(.width(width)) rd_st4_1313  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1313]), .rdlo_in(a4_wr[1377]),  .coef_in(coef[528]), .rdup_out(a5_wr[1313]), .rdlo_out(a5_wr[1377]));
			radix2 #(.width(width)) rd_st4_1314  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1314]), .rdlo_in(a4_wr[1378]),  .coef_in(coef[544]), .rdup_out(a5_wr[1314]), .rdlo_out(a5_wr[1378]));
			radix2 #(.width(width)) rd_st4_1315  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1315]), .rdlo_in(a4_wr[1379]),  .coef_in(coef[560]), .rdup_out(a5_wr[1315]), .rdlo_out(a5_wr[1379]));
			radix2 #(.width(width)) rd_st4_1316  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1316]), .rdlo_in(a4_wr[1380]),  .coef_in(coef[576]), .rdup_out(a5_wr[1316]), .rdlo_out(a5_wr[1380]));
			radix2 #(.width(width)) rd_st4_1317  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1317]), .rdlo_in(a4_wr[1381]),  .coef_in(coef[592]), .rdup_out(a5_wr[1317]), .rdlo_out(a5_wr[1381]));
			radix2 #(.width(width)) rd_st4_1318  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1318]), .rdlo_in(a4_wr[1382]),  .coef_in(coef[608]), .rdup_out(a5_wr[1318]), .rdlo_out(a5_wr[1382]));
			radix2 #(.width(width)) rd_st4_1319  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1319]), .rdlo_in(a4_wr[1383]),  .coef_in(coef[624]), .rdup_out(a5_wr[1319]), .rdlo_out(a5_wr[1383]));
			radix2 #(.width(width)) rd_st4_1320  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1320]), .rdlo_in(a4_wr[1384]),  .coef_in(coef[640]), .rdup_out(a5_wr[1320]), .rdlo_out(a5_wr[1384]));
			radix2 #(.width(width)) rd_st4_1321  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1321]), .rdlo_in(a4_wr[1385]),  .coef_in(coef[656]), .rdup_out(a5_wr[1321]), .rdlo_out(a5_wr[1385]));
			radix2 #(.width(width)) rd_st4_1322  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1322]), .rdlo_in(a4_wr[1386]),  .coef_in(coef[672]), .rdup_out(a5_wr[1322]), .rdlo_out(a5_wr[1386]));
			radix2 #(.width(width)) rd_st4_1323  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1323]), .rdlo_in(a4_wr[1387]),  .coef_in(coef[688]), .rdup_out(a5_wr[1323]), .rdlo_out(a5_wr[1387]));
			radix2 #(.width(width)) rd_st4_1324  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1324]), .rdlo_in(a4_wr[1388]),  .coef_in(coef[704]), .rdup_out(a5_wr[1324]), .rdlo_out(a5_wr[1388]));
			radix2 #(.width(width)) rd_st4_1325  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1325]), .rdlo_in(a4_wr[1389]),  .coef_in(coef[720]), .rdup_out(a5_wr[1325]), .rdlo_out(a5_wr[1389]));
			radix2 #(.width(width)) rd_st4_1326  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1326]), .rdlo_in(a4_wr[1390]),  .coef_in(coef[736]), .rdup_out(a5_wr[1326]), .rdlo_out(a5_wr[1390]));
			radix2 #(.width(width)) rd_st4_1327  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1327]), .rdlo_in(a4_wr[1391]),  .coef_in(coef[752]), .rdup_out(a5_wr[1327]), .rdlo_out(a5_wr[1391]));
			radix2 #(.width(width)) rd_st4_1328  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1328]), .rdlo_in(a4_wr[1392]),  .coef_in(coef[768]), .rdup_out(a5_wr[1328]), .rdlo_out(a5_wr[1392]));
			radix2 #(.width(width)) rd_st4_1329  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1329]), .rdlo_in(a4_wr[1393]),  .coef_in(coef[784]), .rdup_out(a5_wr[1329]), .rdlo_out(a5_wr[1393]));
			radix2 #(.width(width)) rd_st4_1330  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1330]), .rdlo_in(a4_wr[1394]),  .coef_in(coef[800]), .rdup_out(a5_wr[1330]), .rdlo_out(a5_wr[1394]));
			radix2 #(.width(width)) rd_st4_1331  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1331]), .rdlo_in(a4_wr[1395]),  .coef_in(coef[816]), .rdup_out(a5_wr[1331]), .rdlo_out(a5_wr[1395]));
			radix2 #(.width(width)) rd_st4_1332  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1332]), .rdlo_in(a4_wr[1396]),  .coef_in(coef[832]), .rdup_out(a5_wr[1332]), .rdlo_out(a5_wr[1396]));
			radix2 #(.width(width)) rd_st4_1333  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1333]), .rdlo_in(a4_wr[1397]),  .coef_in(coef[848]), .rdup_out(a5_wr[1333]), .rdlo_out(a5_wr[1397]));
			radix2 #(.width(width)) rd_st4_1334  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1334]), .rdlo_in(a4_wr[1398]),  .coef_in(coef[864]), .rdup_out(a5_wr[1334]), .rdlo_out(a5_wr[1398]));
			radix2 #(.width(width)) rd_st4_1335  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1335]), .rdlo_in(a4_wr[1399]),  .coef_in(coef[880]), .rdup_out(a5_wr[1335]), .rdlo_out(a5_wr[1399]));
			radix2 #(.width(width)) rd_st4_1336  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1336]), .rdlo_in(a4_wr[1400]),  .coef_in(coef[896]), .rdup_out(a5_wr[1336]), .rdlo_out(a5_wr[1400]));
			radix2 #(.width(width)) rd_st4_1337  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1337]), .rdlo_in(a4_wr[1401]),  .coef_in(coef[912]), .rdup_out(a5_wr[1337]), .rdlo_out(a5_wr[1401]));
			radix2 #(.width(width)) rd_st4_1338  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1338]), .rdlo_in(a4_wr[1402]),  .coef_in(coef[928]), .rdup_out(a5_wr[1338]), .rdlo_out(a5_wr[1402]));
			radix2 #(.width(width)) rd_st4_1339  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1339]), .rdlo_in(a4_wr[1403]),  .coef_in(coef[944]), .rdup_out(a5_wr[1339]), .rdlo_out(a5_wr[1403]));
			radix2 #(.width(width)) rd_st4_1340  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1340]), .rdlo_in(a4_wr[1404]),  .coef_in(coef[960]), .rdup_out(a5_wr[1340]), .rdlo_out(a5_wr[1404]));
			radix2 #(.width(width)) rd_st4_1341  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1341]), .rdlo_in(a4_wr[1405]),  .coef_in(coef[976]), .rdup_out(a5_wr[1341]), .rdlo_out(a5_wr[1405]));
			radix2 #(.width(width)) rd_st4_1342  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1342]), .rdlo_in(a4_wr[1406]),  .coef_in(coef[992]), .rdup_out(a5_wr[1342]), .rdlo_out(a5_wr[1406]));
			radix2 #(.width(width)) rd_st4_1343  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1343]), .rdlo_in(a4_wr[1407]),  .coef_in(coef[1008]), .rdup_out(a5_wr[1343]), .rdlo_out(a5_wr[1407]));
			radix2 #(.width(width)) rd_st4_1408  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1408]), .rdlo_in(a4_wr[1472]),  .coef_in(coef[0]), .rdup_out(a5_wr[1408]), .rdlo_out(a5_wr[1472]));
			radix2 #(.width(width)) rd_st4_1409  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1409]), .rdlo_in(a4_wr[1473]),  .coef_in(coef[16]), .rdup_out(a5_wr[1409]), .rdlo_out(a5_wr[1473]));
			radix2 #(.width(width)) rd_st4_1410  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1410]), .rdlo_in(a4_wr[1474]),  .coef_in(coef[32]), .rdup_out(a5_wr[1410]), .rdlo_out(a5_wr[1474]));
			radix2 #(.width(width)) rd_st4_1411  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1411]), .rdlo_in(a4_wr[1475]),  .coef_in(coef[48]), .rdup_out(a5_wr[1411]), .rdlo_out(a5_wr[1475]));
			radix2 #(.width(width)) rd_st4_1412  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1412]), .rdlo_in(a4_wr[1476]),  .coef_in(coef[64]), .rdup_out(a5_wr[1412]), .rdlo_out(a5_wr[1476]));
			radix2 #(.width(width)) rd_st4_1413  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1413]), .rdlo_in(a4_wr[1477]),  .coef_in(coef[80]), .rdup_out(a5_wr[1413]), .rdlo_out(a5_wr[1477]));
			radix2 #(.width(width)) rd_st4_1414  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1414]), .rdlo_in(a4_wr[1478]),  .coef_in(coef[96]), .rdup_out(a5_wr[1414]), .rdlo_out(a5_wr[1478]));
			radix2 #(.width(width)) rd_st4_1415  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1415]), .rdlo_in(a4_wr[1479]),  .coef_in(coef[112]), .rdup_out(a5_wr[1415]), .rdlo_out(a5_wr[1479]));
			radix2 #(.width(width)) rd_st4_1416  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1416]), .rdlo_in(a4_wr[1480]),  .coef_in(coef[128]), .rdup_out(a5_wr[1416]), .rdlo_out(a5_wr[1480]));
			radix2 #(.width(width)) rd_st4_1417  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1417]), .rdlo_in(a4_wr[1481]),  .coef_in(coef[144]), .rdup_out(a5_wr[1417]), .rdlo_out(a5_wr[1481]));
			radix2 #(.width(width)) rd_st4_1418  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1418]), .rdlo_in(a4_wr[1482]),  .coef_in(coef[160]), .rdup_out(a5_wr[1418]), .rdlo_out(a5_wr[1482]));
			radix2 #(.width(width)) rd_st4_1419  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1419]), .rdlo_in(a4_wr[1483]),  .coef_in(coef[176]), .rdup_out(a5_wr[1419]), .rdlo_out(a5_wr[1483]));
			radix2 #(.width(width)) rd_st4_1420  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1420]), .rdlo_in(a4_wr[1484]),  .coef_in(coef[192]), .rdup_out(a5_wr[1420]), .rdlo_out(a5_wr[1484]));
			radix2 #(.width(width)) rd_st4_1421  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1421]), .rdlo_in(a4_wr[1485]),  .coef_in(coef[208]), .rdup_out(a5_wr[1421]), .rdlo_out(a5_wr[1485]));
			radix2 #(.width(width)) rd_st4_1422  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1422]), .rdlo_in(a4_wr[1486]),  .coef_in(coef[224]), .rdup_out(a5_wr[1422]), .rdlo_out(a5_wr[1486]));
			radix2 #(.width(width)) rd_st4_1423  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1423]), .rdlo_in(a4_wr[1487]),  .coef_in(coef[240]), .rdup_out(a5_wr[1423]), .rdlo_out(a5_wr[1487]));
			radix2 #(.width(width)) rd_st4_1424  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1424]), .rdlo_in(a4_wr[1488]),  .coef_in(coef[256]), .rdup_out(a5_wr[1424]), .rdlo_out(a5_wr[1488]));
			radix2 #(.width(width)) rd_st4_1425  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1425]), .rdlo_in(a4_wr[1489]),  .coef_in(coef[272]), .rdup_out(a5_wr[1425]), .rdlo_out(a5_wr[1489]));
			radix2 #(.width(width)) rd_st4_1426  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1426]), .rdlo_in(a4_wr[1490]),  .coef_in(coef[288]), .rdup_out(a5_wr[1426]), .rdlo_out(a5_wr[1490]));
			radix2 #(.width(width)) rd_st4_1427  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1427]), .rdlo_in(a4_wr[1491]),  .coef_in(coef[304]), .rdup_out(a5_wr[1427]), .rdlo_out(a5_wr[1491]));
			radix2 #(.width(width)) rd_st4_1428  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1428]), .rdlo_in(a4_wr[1492]),  .coef_in(coef[320]), .rdup_out(a5_wr[1428]), .rdlo_out(a5_wr[1492]));
			radix2 #(.width(width)) rd_st4_1429  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1429]), .rdlo_in(a4_wr[1493]),  .coef_in(coef[336]), .rdup_out(a5_wr[1429]), .rdlo_out(a5_wr[1493]));
			radix2 #(.width(width)) rd_st4_1430  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1430]), .rdlo_in(a4_wr[1494]),  .coef_in(coef[352]), .rdup_out(a5_wr[1430]), .rdlo_out(a5_wr[1494]));
			radix2 #(.width(width)) rd_st4_1431  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1431]), .rdlo_in(a4_wr[1495]),  .coef_in(coef[368]), .rdup_out(a5_wr[1431]), .rdlo_out(a5_wr[1495]));
			radix2 #(.width(width)) rd_st4_1432  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1432]), .rdlo_in(a4_wr[1496]),  .coef_in(coef[384]), .rdup_out(a5_wr[1432]), .rdlo_out(a5_wr[1496]));
			radix2 #(.width(width)) rd_st4_1433  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1433]), .rdlo_in(a4_wr[1497]),  .coef_in(coef[400]), .rdup_out(a5_wr[1433]), .rdlo_out(a5_wr[1497]));
			radix2 #(.width(width)) rd_st4_1434  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1434]), .rdlo_in(a4_wr[1498]),  .coef_in(coef[416]), .rdup_out(a5_wr[1434]), .rdlo_out(a5_wr[1498]));
			radix2 #(.width(width)) rd_st4_1435  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1435]), .rdlo_in(a4_wr[1499]),  .coef_in(coef[432]), .rdup_out(a5_wr[1435]), .rdlo_out(a5_wr[1499]));
			radix2 #(.width(width)) rd_st4_1436  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1436]), .rdlo_in(a4_wr[1500]),  .coef_in(coef[448]), .rdup_out(a5_wr[1436]), .rdlo_out(a5_wr[1500]));
			radix2 #(.width(width)) rd_st4_1437  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1437]), .rdlo_in(a4_wr[1501]),  .coef_in(coef[464]), .rdup_out(a5_wr[1437]), .rdlo_out(a5_wr[1501]));
			radix2 #(.width(width)) rd_st4_1438  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1438]), .rdlo_in(a4_wr[1502]),  .coef_in(coef[480]), .rdup_out(a5_wr[1438]), .rdlo_out(a5_wr[1502]));
			radix2 #(.width(width)) rd_st4_1439  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1439]), .rdlo_in(a4_wr[1503]),  .coef_in(coef[496]), .rdup_out(a5_wr[1439]), .rdlo_out(a5_wr[1503]));
			radix2 #(.width(width)) rd_st4_1440  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1440]), .rdlo_in(a4_wr[1504]),  .coef_in(coef[512]), .rdup_out(a5_wr[1440]), .rdlo_out(a5_wr[1504]));
			radix2 #(.width(width)) rd_st4_1441  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1441]), .rdlo_in(a4_wr[1505]),  .coef_in(coef[528]), .rdup_out(a5_wr[1441]), .rdlo_out(a5_wr[1505]));
			radix2 #(.width(width)) rd_st4_1442  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1442]), .rdlo_in(a4_wr[1506]),  .coef_in(coef[544]), .rdup_out(a5_wr[1442]), .rdlo_out(a5_wr[1506]));
			radix2 #(.width(width)) rd_st4_1443  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1443]), .rdlo_in(a4_wr[1507]),  .coef_in(coef[560]), .rdup_out(a5_wr[1443]), .rdlo_out(a5_wr[1507]));
			radix2 #(.width(width)) rd_st4_1444  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1444]), .rdlo_in(a4_wr[1508]),  .coef_in(coef[576]), .rdup_out(a5_wr[1444]), .rdlo_out(a5_wr[1508]));
			radix2 #(.width(width)) rd_st4_1445  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1445]), .rdlo_in(a4_wr[1509]),  .coef_in(coef[592]), .rdup_out(a5_wr[1445]), .rdlo_out(a5_wr[1509]));
			radix2 #(.width(width)) rd_st4_1446  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1446]), .rdlo_in(a4_wr[1510]),  .coef_in(coef[608]), .rdup_out(a5_wr[1446]), .rdlo_out(a5_wr[1510]));
			radix2 #(.width(width)) rd_st4_1447  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1447]), .rdlo_in(a4_wr[1511]),  .coef_in(coef[624]), .rdup_out(a5_wr[1447]), .rdlo_out(a5_wr[1511]));
			radix2 #(.width(width)) rd_st4_1448  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1448]), .rdlo_in(a4_wr[1512]),  .coef_in(coef[640]), .rdup_out(a5_wr[1448]), .rdlo_out(a5_wr[1512]));
			radix2 #(.width(width)) rd_st4_1449  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1449]), .rdlo_in(a4_wr[1513]),  .coef_in(coef[656]), .rdup_out(a5_wr[1449]), .rdlo_out(a5_wr[1513]));
			radix2 #(.width(width)) rd_st4_1450  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1450]), .rdlo_in(a4_wr[1514]),  .coef_in(coef[672]), .rdup_out(a5_wr[1450]), .rdlo_out(a5_wr[1514]));
			radix2 #(.width(width)) rd_st4_1451  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1451]), .rdlo_in(a4_wr[1515]),  .coef_in(coef[688]), .rdup_out(a5_wr[1451]), .rdlo_out(a5_wr[1515]));
			radix2 #(.width(width)) rd_st4_1452  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1452]), .rdlo_in(a4_wr[1516]),  .coef_in(coef[704]), .rdup_out(a5_wr[1452]), .rdlo_out(a5_wr[1516]));
			radix2 #(.width(width)) rd_st4_1453  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1453]), .rdlo_in(a4_wr[1517]),  .coef_in(coef[720]), .rdup_out(a5_wr[1453]), .rdlo_out(a5_wr[1517]));
			radix2 #(.width(width)) rd_st4_1454  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1454]), .rdlo_in(a4_wr[1518]),  .coef_in(coef[736]), .rdup_out(a5_wr[1454]), .rdlo_out(a5_wr[1518]));
			radix2 #(.width(width)) rd_st4_1455  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1455]), .rdlo_in(a4_wr[1519]),  .coef_in(coef[752]), .rdup_out(a5_wr[1455]), .rdlo_out(a5_wr[1519]));
			radix2 #(.width(width)) rd_st4_1456  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1456]), .rdlo_in(a4_wr[1520]),  .coef_in(coef[768]), .rdup_out(a5_wr[1456]), .rdlo_out(a5_wr[1520]));
			radix2 #(.width(width)) rd_st4_1457  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1457]), .rdlo_in(a4_wr[1521]),  .coef_in(coef[784]), .rdup_out(a5_wr[1457]), .rdlo_out(a5_wr[1521]));
			radix2 #(.width(width)) rd_st4_1458  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1458]), .rdlo_in(a4_wr[1522]),  .coef_in(coef[800]), .rdup_out(a5_wr[1458]), .rdlo_out(a5_wr[1522]));
			radix2 #(.width(width)) rd_st4_1459  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1459]), .rdlo_in(a4_wr[1523]),  .coef_in(coef[816]), .rdup_out(a5_wr[1459]), .rdlo_out(a5_wr[1523]));
			radix2 #(.width(width)) rd_st4_1460  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1460]), .rdlo_in(a4_wr[1524]),  .coef_in(coef[832]), .rdup_out(a5_wr[1460]), .rdlo_out(a5_wr[1524]));
			radix2 #(.width(width)) rd_st4_1461  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1461]), .rdlo_in(a4_wr[1525]),  .coef_in(coef[848]), .rdup_out(a5_wr[1461]), .rdlo_out(a5_wr[1525]));
			radix2 #(.width(width)) rd_st4_1462  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1462]), .rdlo_in(a4_wr[1526]),  .coef_in(coef[864]), .rdup_out(a5_wr[1462]), .rdlo_out(a5_wr[1526]));
			radix2 #(.width(width)) rd_st4_1463  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1463]), .rdlo_in(a4_wr[1527]),  .coef_in(coef[880]), .rdup_out(a5_wr[1463]), .rdlo_out(a5_wr[1527]));
			radix2 #(.width(width)) rd_st4_1464  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1464]), .rdlo_in(a4_wr[1528]),  .coef_in(coef[896]), .rdup_out(a5_wr[1464]), .rdlo_out(a5_wr[1528]));
			radix2 #(.width(width)) rd_st4_1465  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1465]), .rdlo_in(a4_wr[1529]),  .coef_in(coef[912]), .rdup_out(a5_wr[1465]), .rdlo_out(a5_wr[1529]));
			radix2 #(.width(width)) rd_st4_1466  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1466]), .rdlo_in(a4_wr[1530]),  .coef_in(coef[928]), .rdup_out(a5_wr[1466]), .rdlo_out(a5_wr[1530]));
			radix2 #(.width(width)) rd_st4_1467  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1467]), .rdlo_in(a4_wr[1531]),  .coef_in(coef[944]), .rdup_out(a5_wr[1467]), .rdlo_out(a5_wr[1531]));
			radix2 #(.width(width)) rd_st4_1468  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1468]), .rdlo_in(a4_wr[1532]),  .coef_in(coef[960]), .rdup_out(a5_wr[1468]), .rdlo_out(a5_wr[1532]));
			radix2 #(.width(width)) rd_st4_1469  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1469]), .rdlo_in(a4_wr[1533]),  .coef_in(coef[976]), .rdup_out(a5_wr[1469]), .rdlo_out(a5_wr[1533]));
			radix2 #(.width(width)) rd_st4_1470  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1470]), .rdlo_in(a4_wr[1534]),  .coef_in(coef[992]), .rdup_out(a5_wr[1470]), .rdlo_out(a5_wr[1534]));
			radix2 #(.width(width)) rd_st4_1471  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1471]), .rdlo_in(a4_wr[1535]),  .coef_in(coef[1008]), .rdup_out(a5_wr[1471]), .rdlo_out(a5_wr[1535]));
			radix2 #(.width(width)) rd_st4_1536  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1536]), .rdlo_in(a4_wr[1600]),  .coef_in(coef[0]), .rdup_out(a5_wr[1536]), .rdlo_out(a5_wr[1600]));
			radix2 #(.width(width)) rd_st4_1537  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1537]), .rdlo_in(a4_wr[1601]),  .coef_in(coef[16]), .rdup_out(a5_wr[1537]), .rdlo_out(a5_wr[1601]));
			radix2 #(.width(width)) rd_st4_1538  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1538]), .rdlo_in(a4_wr[1602]),  .coef_in(coef[32]), .rdup_out(a5_wr[1538]), .rdlo_out(a5_wr[1602]));
			radix2 #(.width(width)) rd_st4_1539  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1539]), .rdlo_in(a4_wr[1603]),  .coef_in(coef[48]), .rdup_out(a5_wr[1539]), .rdlo_out(a5_wr[1603]));
			radix2 #(.width(width)) rd_st4_1540  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1540]), .rdlo_in(a4_wr[1604]),  .coef_in(coef[64]), .rdup_out(a5_wr[1540]), .rdlo_out(a5_wr[1604]));
			radix2 #(.width(width)) rd_st4_1541  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1541]), .rdlo_in(a4_wr[1605]),  .coef_in(coef[80]), .rdup_out(a5_wr[1541]), .rdlo_out(a5_wr[1605]));
			radix2 #(.width(width)) rd_st4_1542  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1542]), .rdlo_in(a4_wr[1606]),  .coef_in(coef[96]), .rdup_out(a5_wr[1542]), .rdlo_out(a5_wr[1606]));
			radix2 #(.width(width)) rd_st4_1543  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1543]), .rdlo_in(a4_wr[1607]),  .coef_in(coef[112]), .rdup_out(a5_wr[1543]), .rdlo_out(a5_wr[1607]));
			radix2 #(.width(width)) rd_st4_1544  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1544]), .rdlo_in(a4_wr[1608]),  .coef_in(coef[128]), .rdup_out(a5_wr[1544]), .rdlo_out(a5_wr[1608]));
			radix2 #(.width(width)) rd_st4_1545  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1545]), .rdlo_in(a4_wr[1609]),  .coef_in(coef[144]), .rdup_out(a5_wr[1545]), .rdlo_out(a5_wr[1609]));
			radix2 #(.width(width)) rd_st4_1546  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1546]), .rdlo_in(a4_wr[1610]),  .coef_in(coef[160]), .rdup_out(a5_wr[1546]), .rdlo_out(a5_wr[1610]));
			radix2 #(.width(width)) rd_st4_1547  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1547]), .rdlo_in(a4_wr[1611]),  .coef_in(coef[176]), .rdup_out(a5_wr[1547]), .rdlo_out(a5_wr[1611]));
			radix2 #(.width(width)) rd_st4_1548  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1548]), .rdlo_in(a4_wr[1612]),  .coef_in(coef[192]), .rdup_out(a5_wr[1548]), .rdlo_out(a5_wr[1612]));
			radix2 #(.width(width)) rd_st4_1549  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1549]), .rdlo_in(a4_wr[1613]),  .coef_in(coef[208]), .rdup_out(a5_wr[1549]), .rdlo_out(a5_wr[1613]));
			radix2 #(.width(width)) rd_st4_1550  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1550]), .rdlo_in(a4_wr[1614]),  .coef_in(coef[224]), .rdup_out(a5_wr[1550]), .rdlo_out(a5_wr[1614]));
			radix2 #(.width(width)) rd_st4_1551  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1551]), .rdlo_in(a4_wr[1615]),  .coef_in(coef[240]), .rdup_out(a5_wr[1551]), .rdlo_out(a5_wr[1615]));
			radix2 #(.width(width)) rd_st4_1552  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1552]), .rdlo_in(a4_wr[1616]),  .coef_in(coef[256]), .rdup_out(a5_wr[1552]), .rdlo_out(a5_wr[1616]));
			radix2 #(.width(width)) rd_st4_1553  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1553]), .rdlo_in(a4_wr[1617]),  .coef_in(coef[272]), .rdup_out(a5_wr[1553]), .rdlo_out(a5_wr[1617]));
			radix2 #(.width(width)) rd_st4_1554  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1554]), .rdlo_in(a4_wr[1618]),  .coef_in(coef[288]), .rdup_out(a5_wr[1554]), .rdlo_out(a5_wr[1618]));
			radix2 #(.width(width)) rd_st4_1555  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1555]), .rdlo_in(a4_wr[1619]),  .coef_in(coef[304]), .rdup_out(a5_wr[1555]), .rdlo_out(a5_wr[1619]));
			radix2 #(.width(width)) rd_st4_1556  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1556]), .rdlo_in(a4_wr[1620]),  .coef_in(coef[320]), .rdup_out(a5_wr[1556]), .rdlo_out(a5_wr[1620]));
			radix2 #(.width(width)) rd_st4_1557  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1557]), .rdlo_in(a4_wr[1621]),  .coef_in(coef[336]), .rdup_out(a5_wr[1557]), .rdlo_out(a5_wr[1621]));
			radix2 #(.width(width)) rd_st4_1558  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1558]), .rdlo_in(a4_wr[1622]),  .coef_in(coef[352]), .rdup_out(a5_wr[1558]), .rdlo_out(a5_wr[1622]));
			radix2 #(.width(width)) rd_st4_1559  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1559]), .rdlo_in(a4_wr[1623]),  .coef_in(coef[368]), .rdup_out(a5_wr[1559]), .rdlo_out(a5_wr[1623]));
			radix2 #(.width(width)) rd_st4_1560  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1560]), .rdlo_in(a4_wr[1624]),  .coef_in(coef[384]), .rdup_out(a5_wr[1560]), .rdlo_out(a5_wr[1624]));
			radix2 #(.width(width)) rd_st4_1561  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1561]), .rdlo_in(a4_wr[1625]),  .coef_in(coef[400]), .rdup_out(a5_wr[1561]), .rdlo_out(a5_wr[1625]));
			radix2 #(.width(width)) rd_st4_1562  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1562]), .rdlo_in(a4_wr[1626]),  .coef_in(coef[416]), .rdup_out(a5_wr[1562]), .rdlo_out(a5_wr[1626]));
			radix2 #(.width(width)) rd_st4_1563  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1563]), .rdlo_in(a4_wr[1627]),  .coef_in(coef[432]), .rdup_out(a5_wr[1563]), .rdlo_out(a5_wr[1627]));
			radix2 #(.width(width)) rd_st4_1564  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1564]), .rdlo_in(a4_wr[1628]),  .coef_in(coef[448]), .rdup_out(a5_wr[1564]), .rdlo_out(a5_wr[1628]));
			radix2 #(.width(width)) rd_st4_1565  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1565]), .rdlo_in(a4_wr[1629]),  .coef_in(coef[464]), .rdup_out(a5_wr[1565]), .rdlo_out(a5_wr[1629]));
			radix2 #(.width(width)) rd_st4_1566  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1566]), .rdlo_in(a4_wr[1630]),  .coef_in(coef[480]), .rdup_out(a5_wr[1566]), .rdlo_out(a5_wr[1630]));
			radix2 #(.width(width)) rd_st4_1567  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1567]), .rdlo_in(a4_wr[1631]),  .coef_in(coef[496]), .rdup_out(a5_wr[1567]), .rdlo_out(a5_wr[1631]));
			radix2 #(.width(width)) rd_st4_1568  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1568]), .rdlo_in(a4_wr[1632]),  .coef_in(coef[512]), .rdup_out(a5_wr[1568]), .rdlo_out(a5_wr[1632]));
			radix2 #(.width(width)) rd_st4_1569  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1569]), .rdlo_in(a4_wr[1633]),  .coef_in(coef[528]), .rdup_out(a5_wr[1569]), .rdlo_out(a5_wr[1633]));
			radix2 #(.width(width)) rd_st4_1570  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1570]), .rdlo_in(a4_wr[1634]),  .coef_in(coef[544]), .rdup_out(a5_wr[1570]), .rdlo_out(a5_wr[1634]));
			radix2 #(.width(width)) rd_st4_1571  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1571]), .rdlo_in(a4_wr[1635]),  .coef_in(coef[560]), .rdup_out(a5_wr[1571]), .rdlo_out(a5_wr[1635]));
			radix2 #(.width(width)) rd_st4_1572  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1572]), .rdlo_in(a4_wr[1636]),  .coef_in(coef[576]), .rdup_out(a5_wr[1572]), .rdlo_out(a5_wr[1636]));
			radix2 #(.width(width)) rd_st4_1573  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1573]), .rdlo_in(a4_wr[1637]),  .coef_in(coef[592]), .rdup_out(a5_wr[1573]), .rdlo_out(a5_wr[1637]));
			radix2 #(.width(width)) rd_st4_1574  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1574]), .rdlo_in(a4_wr[1638]),  .coef_in(coef[608]), .rdup_out(a5_wr[1574]), .rdlo_out(a5_wr[1638]));
			radix2 #(.width(width)) rd_st4_1575  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1575]), .rdlo_in(a4_wr[1639]),  .coef_in(coef[624]), .rdup_out(a5_wr[1575]), .rdlo_out(a5_wr[1639]));
			radix2 #(.width(width)) rd_st4_1576  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1576]), .rdlo_in(a4_wr[1640]),  .coef_in(coef[640]), .rdup_out(a5_wr[1576]), .rdlo_out(a5_wr[1640]));
			radix2 #(.width(width)) rd_st4_1577  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1577]), .rdlo_in(a4_wr[1641]),  .coef_in(coef[656]), .rdup_out(a5_wr[1577]), .rdlo_out(a5_wr[1641]));
			radix2 #(.width(width)) rd_st4_1578  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1578]), .rdlo_in(a4_wr[1642]),  .coef_in(coef[672]), .rdup_out(a5_wr[1578]), .rdlo_out(a5_wr[1642]));
			radix2 #(.width(width)) rd_st4_1579  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1579]), .rdlo_in(a4_wr[1643]),  .coef_in(coef[688]), .rdup_out(a5_wr[1579]), .rdlo_out(a5_wr[1643]));
			radix2 #(.width(width)) rd_st4_1580  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1580]), .rdlo_in(a4_wr[1644]),  .coef_in(coef[704]), .rdup_out(a5_wr[1580]), .rdlo_out(a5_wr[1644]));
			radix2 #(.width(width)) rd_st4_1581  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1581]), .rdlo_in(a4_wr[1645]),  .coef_in(coef[720]), .rdup_out(a5_wr[1581]), .rdlo_out(a5_wr[1645]));
			radix2 #(.width(width)) rd_st4_1582  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1582]), .rdlo_in(a4_wr[1646]),  .coef_in(coef[736]), .rdup_out(a5_wr[1582]), .rdlo_out(a5_wr[1646]));
			radix2 #(.width(width)) rd_st4_1583  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1583]), .rdlo_in(a4_wr[1647]),  .coef_in(coef[752]), .rdup_out(a5_wr[1583]), .rdlo_out(a5_wr[1647]));
			radix2 #(.width(width)) rd_st4_1584  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1584]), .rdlo_in(a4_wr[1648]),  .coef_in(coef[768]), .rdup_out(a5_wr[1584]), .rdlo_out(a5_wr[1648]));
			radix2 #(.width(width)) rd_st4_1585  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1585]), .rdlo_in(a4_wr[1649]),  .coef_in(coef[784]), .rdup_out(a5_wr[1585]), .rdlo_out(a5_wr[1649]));
			radix2 #(.width(width)) rd_st4_1586  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1586]), .rdlo_in(a4_wr[1650]),  .coef_in(coef[800]), .rdup_out(a5_wr[1586]), .rdlo_out(a5_wr[1650]));
			radix2 #(.width(width)) rd_st4_1587  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1587]), .rdlo_in(a4_wr[1651]),  .coef_in(coef[816]), .rdup_out(a5_wr[1587]), .rdlo_out(a5_wr[1651]));
			radix2 #(.width(width)) rd_st4_1588  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1588]), .rdlo_in(a4_wr[1652]),  .coef_in(coef[832]), .rdup_out(a5_wr[1588]), .rdlo_out(a5_wr[1652]));
			radix2 #(.width(width)) rd_st4_1589  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1589]), .rdlo_in(a4_wr[1653]),  .coef_in(coef[848]), .rdup_out(a5_wr[1589]), .rdlo_out(a5_wr[1653]));
			radix2 #(.width(width)) rd_st4_1590  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1590]), .rdlo_in(a4_wr[1654]),  .coef_in(coef[864]), .rdup_out(a5_wr[1590]), .rdlo_out(a5_wr[1654]));
			radix2 #(.width(width)) rd_st4_1591  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1591]), .rdlo_in(a4_wr[1655]),  .coef_in(coef[880]), .rdup_out(a5_wr[1591]), .rdlo_out(a5_wr[1655]));
			radix2 #(.width(width)) rd_st4_1592  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1592]), .rdlo_in(a4_wr[1656]),  .coef_in(coef[896]), .rdup_out(a5_wr[1592]), .rdlo_out(a5_wr[1656]));
			radix2 #(.width(width)) rd_st4_1593  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1593]), .rdlo_in(a4_wr[1657]),  .coef_in(coef[912]), .rdup_out(a5_wr[1593]), .rdlo_out(a5_wr[1657]));
			radix2 #(.width(width)) rd_st4_1594  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1594]), .rdlo_in(a4_wr[1658]),  .coef_in(coef[928]), .rdup_out(a5_wr[1594]), .rdlo_out(a5_wr[1658]));
			radix2 #(.width(width)) rd_st4_1595  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1595]), .rdlo_in(a4_wr[1659]),  .coef_in(coef[944]), .rdup_out(a5_wr[1595]), .rdlo_out(a5_wr[1659]));
			radix2 #(.width(width)) rd_st4_1596  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1596]), .rdlo_in(a4_wr[1660]),  .coef_in(coef[960]), .rdup_out(a5_wr[1596]), .rdlo_out(a5_wr[1660]));
			radix2 #(.width(width)) rd_st4_1597  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1597]), .rdlo_in(a4_wr[1661]),  .coef_in(coef[976]), .rdup_out(a5_wr[1597]), .rdlo_out(a5_wr[1661]));
			radix2 #(.width(width)) rd_st4_1598  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1598]), .rdlo_in(a4_wr[1662]),  .coef_in(coef[992]), .rdup_out(a5_wr[1598]), .rdlo_out(a5_wr[1662]));
			radix2 #(.width(width)) rd_st4_1599  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1599]), .rdlo_in(a4_wr[1663]),  .coef_in(coef[1008]), .rdup_out(a5_wr[1599]), .rdlo_out(a5_wr[1663]));
			radix2 #(.width(width)) rd_st4_1664  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1664]), .rdlo_in(a4_wr[1728]),  .coef_in(coef[0]), .rdup_out(a5_wr[1664]), .rdlo_out(a5_wr[1728]));
			radix2 #(.width(width)) rd_st4_1665  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1665]), .rdlo_in(a4_wr[1729]),  .coef_in(coef[16]), .rdup_out(a5_wr[1665]), .rdlo_out(a5_wr[1729]));
			radix2 #(.width(width)) rd_st4_1666  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1666]), .rdlo_in(a4_wr[1730]),  .coef_in(coef[32]), .rdup_out(a5_wr[1666]), .rdlo_out(a5_wr[1730]));
			radix2 #(.width(width)) rd_st4_1667  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1667]), .rdlo_in(a4_wr[1731]),  .coef_in(coef[48]), .rdup_out(a5_wr[1667]), .rdlo_out(a5_wr[1731]));
			radix2 #(.width(width)) rd_st4_1668  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1668]), .rdlo_in(a4_wr[1732]),  .coef_in(coef[64]), .rdup_out(a5_wr[1668]), .rdlo_out(a5_wr[1732]));
			radix2 #(.width(width)) rd_st4_1669  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1669]), .rdlo_in(a4_wr[1733]),  .coef_in(coef[80]), .rdup_out(a5_wr[1669]), .rdlo_out(a5_wr[1733]));
			radix2 #(.width(width)) rd_st4_1670  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1670]), .rdlo_in(a4_wr[1734]),  .coef_in(coef[96]), .rdup_out(a5_wr[1670]), .rdlo_out(a5_wr[1734]));
			radix2 #(.width(width)) rd_st4_1671  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1671]), .rdlo_in(a4_wr[1735]),  .coef_in(coef[112]), .rdup_out(a5_wr[1671]), .rdlo_out(a5_wr[1735]));
			radix2 #(.width(width)) rd_st4_1672  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1672]), .rdlo_in(a4_wr[1736]),  .coef_in(coef[128]), .rdup_out(a5_wr[1672]), .rdlo_out(a5_wr[1736]));
			radix2 #(.width(width)) rd_st4_1673  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1673]), .rdlo_in(a4_wr[1737]),  .coef_in(coef[144]), .rdup_out(a5_wr[1673]), .rdlo_out(a5_wr[1737]));
			radix2 #(.width(width)) rd_st4_1674  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1674]), .rdlo_in(a4_wr[1738]),  .coef_in(coef[160]), .rdup_out(a5_wr[1674]), .rdlo_out(a5_wr[1738]));
			radix2 #(.width(width)) rd_st4_1675  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1675]), .rdlo_in(a4_wr[1739]),  .coef_in(coef[176]), .rdup_out(a5_wr[1675]), .rdlo_out(a5_wr[1739]));
			radix2 #(.width(width)) rd_st4_1676  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1676]), .rdlo_in(a4_wr[1740]),  .coef_in(coef[192]), .rdup_out(a5_wr[1676]), .rdlo_out(a5_wr[1740]));
			radix2 #(.width(width)) rd_st4_1677  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1677]), .rdlo_in(a4_wr[1741]),  .coef_in(coef[208]), .rdup_out(a5_wr[1677]), .rdlo_out(a5_wr[1741]));
			radix2 #(.width(width)) rd_st4_1678  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1678]), .rdlo_in(a4_wr[1742]),  .coef_in(coef[224]), .rdup_out(a5_wr[1678]), .rdlo_out(a5_wr[1742]));
			radix2 #(.width(width)) rd_st4_1679  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1679]), .rdlo_in(a4_wr[1743]),  .coef_in(coef[240]), .rdup_out(a5_wr[1679]), .rdlo_out(a5_wr[1743]));
			radix2 #(.width(width)) rd_st4_1680  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1680]), .rdlo_in(a4_wr[1744]),  .coef_in(coef[256]), .rdup_out(a5_wr[1680]), .rdlo_out(a5_wr[1744]));
			radix2 #(.width(width)) rd_st4_1681  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1681]), .rdlo_in(a4_wr[1745]),  .coef_in(coef[272]), .rdup_out(a5_wr[1681]), .rdlo_out(a5_wr[1745]));
			radix2 #(.width(width)) rd_st4_1682  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1682]), .rdlo_in(a4_wr[1746]),  .coef_in(coef[288]), .rdup_out(a5_wr[1682]), .rdlo_out(a5_wr[1746]));
			radix2 #(.width(width)) rd_st4_1683  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1683]), .rdlo_in(a4_wr[1747]),  .coef_in(coef[304]), .rdup_out(a5_wr[1683]), .rdlo_out(a5_wr[1747]));
			radix2 #(.width(width)) rd_st4_1684  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1684]), .rdlo_in(a4_wr[1748]),  .coef_in(coef[320]), .rdup_out(a5_wr[1684]), .rdlo_out(a5_wr[1748]));
			radix2 #(.width(width)) rd_st4_1685  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1685]), .rdlo_in(a4_wr[1749]),  .coef_in(coef[336]), .rdup_out(a5_wr[1685]), .rdlo_out(a5_wr[1749]));
			radix2 #(.width(width)) rd_st4_1686  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1686]), .rdlo_in(a4_wr[1750]),  .coef_in(coef[352]), .rdup_out(a5_wr[1686]), .rdlo_out(a5_wr[1750]));
			radix2 #(.width(width)) rd_st4_1687  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1687]), .rdlo_in(a4_wr[1751]),  .coef_in(coef[368]), .rdup_out(a5_wr[1687]), .rdlo_out(a5_wr[1751]));
			radix2 #(.width(width)) rd_st4_1688  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1688]), .rdlo_in(a4_wr[1752]),  .coef_in(coef[384]), .rdup_out(a5_wr[1688]), .rdlo_out(a5_wr[1752]));
			radix2 #(.width(width)) rd_st4_1689  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1689]), .rdlo_in(a4_wr[1753]),  .coef_in(coef[400]), .rdup_out(a5_wr[1689]), .rdlo_out(a5_wr[1753]));
			radix2 #(.width(width)) rd_st4_1690  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1690]), .rdlo_in(a4_wr[1754]),  .coef_in(coef[416]), .rdup_out(a5_wr[1690]), .rdlo_out(a5_wr[1754]));
			radix2 #(.width(width)) rd_st4_1691  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1691]), .rdlo_in(a4_wr[1755]),  .coef_in(coef[432]), .rdup_out(a5_wr[1691]), .rdlo_out(a5_wr[1755]));
			radix2 #(.width(width)) rd_st4_1692  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1692]), .rdlo_in(a4_wr[1756]),  .coef_in(coef[448]), .rdup_out(a5_wr[1692]), .rdlo_out(a5_wr[1756]));
			radix2 #(.width(width)) rd_st4_1693  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1693]), .rdlo_in(a4_wr[1757]),  .coef_in(coef[464]), .rdup_out(a5_wr[1693]), .rdlo_out(a5_wr[1757]));
			radix2 #(.width(width)) rd_st4_1694  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1694]), .rdlo_in(a4_wr[1758]),  .coef_in(coef[480]), .rdup_out(a5_wr[1694]), .rdlo_out(a5_wr[1758]));
			radix2 #(.width(width)) rd_st4_1695  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1695]), .rdlo_in(a4_wr[1759]),  .coef_in(coef[496]), .rdup_out(a5_wr[1695]), .rdlo_out(a5_wr[1759]));
			radix2 #(.width(width)) rd_st4_1696  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1696]), .rdlo_in(a4_wr[1760]),  .coef_in(coef[512]), .rdup_out(a5_wr[1696]), .rdlo_out(a5_wr[1760]));
			radix2 #(.width(width)) rd_st4_1697  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1697]), .rdlo_in(a4_wr[1761]),  .coef_in(coef[528]), .rdup_out(a5_wr[1697]), .rdlo_out(a5_wr[1761]));
			radix2 #(.width(width)) rd_st4_1698  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1698]), .rdlo_in(a4_wr[1762]),  .coef_in(coef[544]), .rdup_out(a5_wr[1698]), .rdlo_out(a5_wr[1762]));
			radix2 #(.width(width)) rd_st4_1699  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1699]), .rdlo_in(a4_wr[1763]),  .coef_in(coef[560]), .rdup_out(a5_wr[1699]), .rdlo_out(a5_wr[1763]));
			radix2 #(.width(width)) rd_st4_1700  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1700]), .rdlo_in(a4_wr[1764]),  .coef_in(coef[576]), .rdup_out(a5_wr[1700]), .rdlo_out(a5_wr[1764]));
			radix2 #(.width(width)) rd_st4_1701  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1701]), .rdlo_in(a4_wr[1765]),  .coef_in(coef[592]), .rdup_out(a5_wr[1701]), .rdlo_out(a5_wr[1765]));
			radix2 #(.width(width)) rd_st4_1702  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1702]), .rdlo_in(a4_wr[1766]),  .coef_in(coef[608]), .rdup_out(a5_wr[1702]), .rdlo_out(a5_wr[1766]));
			radix2 #(.width(width)) rd_st4_1703  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1703]), .rdlo_in(a4_wr[1767]),  .coef_in(coef[624]), .rdup_out(a5_wr[1703]), .rdlo_out(a5_wr[1767]));
			radix2 #(.width(width)) rd_st4_1704  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1704]), .rdlo_in(a4_wr[1768]),  .coef_in(coef[640]), .rdup_out(a5_wr[1704]), .rdlo_out(a5_wr[1768]));
			radix2 #(.width(width)) rd_st4_1705  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1705]), .rdlo_in(a4_wr[1769]),  .coef_in(coef[656]), .rdup_out(a5_wr[1705]), .rdlo_out(a5_wr[1769]));
			radix2 #(.width(width)) rd_st4_1706  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1706]), .rdlo_in(a4_wr[1770]),  .coef_in(coef[672]), .rdup_out(a5_wr[1706]), .rdlo_out(a5_wr[1770]));
			radix2 #(.width(width)) rd_st4_1707  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1707]), .rdlo_in(a4_wr[1771]),  .coef_in(coef[688]), .rdup_out(a5_wr[1707]), .rdlo_out(a5_wr[1771]));
			radix2 #(.width(width)) rd_st4_1708  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1708]), .rdlo_in(a4_wr[1772]),  .coef_in(coef[704]), .rdup_out(a5_wr[1708]), .rdlo_out(a5_wr[1772]));
			radix2 #(.width(width)) rd_st4_1709  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1709]), .rdlo_in(a4_wr[1773]),  .coef_in(coef[720]), .rdup_out(a5_wr[1709]), .rdlo_out(a5_wr[1773]));
			radix2 #(.width(width)) rd_st4_1710  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1710]), .rdlo_in(a4_wr[1774]),  .coef_in(coef[736]), .rdup_out(a5_wr[1710]), .rdlo_out(a5_wr[1774]));
			radix2 #(.width(width)) rd_st4_1711  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1711]), .rdlo_in(a4_wr[1775]),  .coef_in(coef[752]), .rdup_out(a5_wr[1711]), .rdlo_out(a5_wr[1775]));
			radix2 #(.width(width)) rd_st4_1712  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1712]), .rdlo_in(a4_wr[1776]),  .coef_in(coef[768]), .rdup_out(a5_wr[1712]), .rdlo_out(a5_wr[1776]));
			radix2 #(.width(width)) rd_st4_1713  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1713]), .rdlo_in(a4_wr[1777]),  .coef_in(coef[784]), .rdup_out(a5_wr[1713]), .rdlo_out(a5_wr[1777]));
			radix2 #(.width(width)) rd_st4_1714  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1714]), .rdlo_in(a4_wr[1778]),  .coef_in(coef[800]), .rdup_out(a5_wr[1714]), .rdlo_out(a5_wr[1778]));
			radix2 #(.width(width)) rd_st4_1715  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1715]), .rdlo_in(a4_wr[1779]),  .coef_in(coef[816]), .rdup_out(a5_wr[1715]), .rdlo_out(a5_wr[1779]));
			radix2 #(.width(width)) rd_st4_1716  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1716]), .rdlo_in(a4_wr[1780]),  .coef_in(coef[832]), .rdup_out(a5_wr[1716]), .rdlo_out(a5_wr[1780]));
			radix2 #(.width(width)) rd_st4_1717  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1717]), .rdlo_in(a4_wr[1781]),  .coef_in(coef[848]), .rdup_out(a5_wr[1717]), .rdlo_out(a5_wr[1781]));
			radix2 #(.width(width)) rd_st4_1718  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1718]), .rdlo_in(a4_wr[1782]),  .coef_in(coef[864]), .rdup_out(a5_wr[1718]), .rdlo_out(a5_wr[1782]));
			radix2 #(.width(width)) rd_st4_1719  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1719]), .rdlo_in(a4_wr[1783]),  .coef_in(coef[880]), .rdup_out(a5_wr[1719]), .rdlo_out(a5_wr[1783]));
			radix2 #(.width(width)) rd_st4_1720  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1720]), .rdlo_in(a4_wr[1784]),  .coef_in(coef[896]), .rdup_out(a5_wr[1720]), .rdlo_out(a5_wr[1784]));
			radix2 #(.width(width)) rd_st4_1721  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1721]), .rdlo_in(a4_wr[1785]),  .coef_in(coef[912]), .rdup_out(a5_wr[1721]), .rdlo_out(a5_wr[1785]));
			radix2 #(.width(width)) rd_st4_1722  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1722]), .rdlo_in(a4_wr[1786]),  .coef_in(coef[928]), .rdup_out(a5_wr[1722]), .rdlo_out(a5_wr[1786]));
			radix2 #(.width(width)) rd_st4_1723  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1723]), .rdlo_in(a4_wr[1787]),  .coef_in(coef[944]), .rdup_out(a5_wr[1723]), .rdlo_out(a5_wr[1787]));
			radix2 #(.width(width)) rd_st4_1724  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1724]), .rdlo_in(a4_wr[1788]),  .coef_in(coef[960]), .rdup_out(a5_wr[1724]), .rdlo_out(a5_wr[1788]));
			radix2 #(.width(width)) rd_st4_1725  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1725]), .rdlo_in(a4_wr[1789]),  .coef_in(coef[976]), .rdup_out(a5_wr[1725]), .rdlo_out(a5_wr[1789]));
			radix2 #(.width(width)) rd_st4_1726  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1726]), .rdlo_in(a4_wr[1790]),  .coef_in(coef[992]), .rdup_out(a5_wr[1726]), .rdlo_out(a5_wr[1790]));
			radix2 #(.width(width)) rd_st4_1727  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1727]), .rdlo_in(a4_wr[1791]),  .coef_in(coef[1008]), .rdup_out(a5_wr[1727]), .rdlo_out(a5_wr[1791]));
			radix2 #(.width(width)) rd_st4_1792  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1792]), .rdlo_in(a4_wr[1856]),  .coef_in(coef[0]), .rdup_out(a5_wr[1792]), .rdlo_out(a5_wr[1856]));
			radix2 #(.width(width)) rd_st4_1793  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1793]), .rdlo_in(a4_wr[1857]),  .coef_in(coef[16]), .rdup_out(a5_wr[1793]), .rdlo_out(a5_wr[1857]));
			radix2 #(.width(width)) rd_st4_1794  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1794]), .rdlo_in(a4_wr[1858]),  .coef_in(coef[32]), .rdup_out(a5_wr[1794]), .rdlo_out(a5_wr[1858]));
			radix2 #(.width(width)) rd_st4_1795  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1795]), .rdlo_in(a4_wr[1859]),  .coef_in(coef[48]), .rdup_out(a5_wr[1795]), .rdlo_out(a5_wr[1859]));
			radix2 #(.width(width)) rd_st4_1796  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1796]), .rdlo_in(a4_wr[1860]),  .coef_in(coef[64]), .rdup_out(a5_wr[1796]), .rdlo_out(a5_wr[1860]));
			radix2 #(.width(width)) rd_st4_1797  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1797]), .rdlo_in(a4_wr[1861]),  .coef_in(coef[80]), .rdup_out(a5_wr[1797]), .rdlo_out(a5_wr[1861]));
			radix2 #(.width(width)) rd_st4_1798  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1798]), .rdlo_in(a4_wr[1862]),  .coef_in(coef[96]), .rdup_out(a5_wr[1798]), .rdlo_out(a5_wr[1862]));
			radix2 #(.width(width)) rd_st4_1799  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1799]), .rdlo_in(a4_wr[1863]),  .coef_in(coef[112]), .rdup_out(a5_wr[1799]), .rdlo_out(a5_wr[1863]));
			radix2 #(.width(width)) rd_st4_1800  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1800]), .rdlo_in(a4_wr[1864]),  .coef_in(coef[128]), .rdup_out(a5_wr[1800]), .rdlo_out(a5_wr[1864]));
			radix2 #(.width(width)) rd_st4_1801  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1801]), .rdlo_in(a4_wr[1865]),  .coef_in(coef[144]), .rdup_out(a5_wr[1801]), .rdlo_out(a5_wr[1865]));
			radix2 #(.width(width)) rd_st4_1802  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1802]), .rdlo_in(a4_wr[1866]),  .coef_in(coef[160]), .rdup_out(a5_wr[1802]), .rdlo_out(a5_wr[1866]));
			radix2 #(.width(width)) rd_st4_1803  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1803]), .rdlo_in(a4_wr[1867]),  .coef_in(coef[176]), .rdup_out(a5_wr[1803]), .rdlo_out(a5_wr[1867]));
			radix2 #(.width(width)) rd_st4_1804  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1804]), .rdlo_in(a4_wr[1868]),  .coef_in(coef[192]), .rdup_out(a5_wr[1804]), .rdlo_out(a5_wr[1868]));
			radix2 #(.width(width)) rd_st4_1805  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1805]), .rdlo_in(a4_wr[1869]),  .coef_in(coef[208]), .rdup_out(a5_wr[1805]), .rdlo_out(a5_wr[1869]));
			radix2 #(.width(width)) rd_st4_1806  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1806]), .rdlo_in(a4_wr[1870]),  .coef_in(coef[224]), .rdup_out(a5_wr[1806]), .rdlo_out(a5_wr[1870]));
			radix2 #(.width(width)) rd_st4_1807  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1807]), .rdlo_in(a4_wr[1871]),  .coef_in(coef[240]), .rdup_out(a5_wr[1807]), .rdlo_out(a5_wr[1871]));
			radix2 #(.width(width)) rd_st4_1808  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1808]), .rdlo_in(a4_wr[1872]),  .coef_in(coef[256]), .rdup_out(a5_wr[1808]), .rdlo_out(a5_wr[1872]));
			radix2 #(.width(width)) rd_st4_1809  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1809]), .rdlo_in(a4_wr[1873]),  .coef_in(coef[272]), .rdup_out(a5_wr[1809]), .rdlo_out(a5_wr[1873]));
			radix2 #(.width(width)) rd_st4_1810  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1810]), .rdlo_in(a4_wr[1874]),  .coef_in(coef[288]), .rdup_out(a5_wr[1810]), .rdlo_out(a5_wr[1874]));
			radix2 #(.width(width)) rd_st4_1811  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1811]), .rdlo_in(a4_wr[1875]),  .coef_in(coef[304]), .rdup_out(a5_wr[1811]), .rdlo_out(a5_wr[1875]));
			radix2 #(.width(width)) rd_st4_1812  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1812]), .rdlo_in(a4_wr[1876]),  .coef_in(coef[320]), .rdup_out(a5_wr[1812]), .rdlo_out(a5_wr[1876]));
			radix2 #(.width(width)) rd_st4_1813  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1813]), .rdlo_in(a4_wr[1877]),  .coef_in(coef[336]), .rdup_out(a5_wr[1813]), .rdlo_out(a5_wr[1877]));
			radix2 #(.width(width)) rd_st4_1814  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1814]), .rdlo_in(a4_wr[1878]),  .coef_in(coef[352]), .rdup_out(a5_wr[1814]), .rdlo_out(a5_wr[1878]));
			radix2 #(.width(width)) rd_st4_1815  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1815]), .rdlo_in(a4_wr[1879]),  .coef_in(coef[368]), .rdup_out(a5_wr[1815]), .rdlo_out(a5_wr[1879]));
			radix2 #(.width(width)) rd_st4_1816  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1816]), .rdlo_in(a4_wr[1880]),  .coef_in(coef[384]), .rdup_out(a5_wr[1816]), .rdlo_out(a5_wr[1880]));
			radix2 #(.width(width)) rd_st4_1817  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1817]), .rdlo_in(a4_wr[1881]),  .coef_in(coef[400]), .rdup_out(a5_wr[1817]), .rdlo_out(a5_wr[1881]));
			radix2 #(.width(width)) rd_st4_1818  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1818]), .rdlo_in(a4_wr[1882]),  .coef_in(coef[416]), .rdup_out(a5_wr[1818]), .rdlo_out(a5_wr[1882]));
			radix2 #(.width(width)) rd_st4_1819  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1819]), .rdlo_in(a4_wr[1883]),  .coef_in(coef[432]), .rdup_out(a5_wr[1819]), .rdlo_out(a5_wr[1883]));
			radix2 #(.width(width)) rd_st4_1820  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1820]), .rdlo_in(a4_wr[1884]),  .coef_in(coef[448]), .rdup_out(a5_wr[1820]), .rdlo_out(a5_wr[1884]));
			radix2 #(.width(width)) rd_st4_1821  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1821]), .rdlo_in(a4_wr[1885]),  .coef_in(coef[464]), .rdup_out(a5_wr[1821]), .rdlo_out(a5_wr[1885]));
			radix2 #(.width(width)) rd_st4_1822  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1822]), .rdlo_in(a4_wr[1886]),  .coef_in(coef[480]), .rdup_out(a5_wr[1822]), .rdlo_out(a5_wr[1886]));
			radix2 #(.width(width)) rd_st4_1823  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1823]), .rdlo_in(a4_wr[1887]),  .coef_in(coef[496]), .rdup_out(a5_wr[1823]), .rdlo_out(a5_wr[1887]));
			radix2 #(.width(width)) rd_st4_1824  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1824]), .rdlo_in(a4_wr[1888]),  .coef_in(coef[512]), .rdup_out(a5_wr[1824]), .rdlo_out(a5_wr[1888]));
			radix2 #(.width(width)) rd_st4_1825  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1825]), .rdlo_in(a4_wr[1889]),  .coef_in(coef[528]), .rdup_out(a5_wr[1825]), .rdlo_out(a5_wr[1889]));
			radix2 #(.width(width)) rd_st4_1826  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1826]), .rdlo_in(a4_wr[1890]),  .coef_in(coef[544]), .rdup_out(a5_wr[1826]), .rdlo_out(a5_wr[1890]));
			radix2 #(.width(width)) rd_st4_1827  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1827]), .rdlo_in(a4_wr[1891]),  .coef_in(coef[560]), .rdup_out(a5_wr[1827]), .rdlo_out(a5_wr[1891]));
			radix2 #(.width(width)) rd_st4_1828  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1828]), .rdlo_in(a4_wr[1892]),  .coef_in(coef[576]), .rdup_out(a5_wr[1828]), .rdlo_out(a5_wr[1892]));
			radix2 #(.width(width)) rd_st4_1829  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1829]), .rdlo_in(a4_wr[1893]),  .coef_in(coef[592]), .rdup_out(a5_wr[1829]), .rdlo_out(a5_wr[1893]));
			radix2 #(.width(width)) rd_st4_1830  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1830]), .rdlo_in(a4_wr[1894]),  .coef_in(coef[608]), .rdup_out(a5_wr[1830]), .rdlo_out(a5_wr[1894]));
			radix2 #(.width(width)) rd_st4_1831  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1831]), .rdlo_in(a4_wr[1895]),  .coef_in(coef[624]), .rdup_out(a5_wr[1831]), .rdlo_out(a5_wr[1895]));
			radix2 #(.width(width)) rd_st4_1832  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1832]), .rdlo_in(a4_wr[1896]),  .coef_in(coef[640]), .rdup_out(a5_wr[1832]), .rdlo_out(a5_wr[1896]));
			radix2 #(.width(width)) rd_st4_1833  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1833]), .rdlo_in(a4_wr[1897]),  .coef_in(coef[656]), .rdup_out(a5_wr[1833]), .rdlo_out(a5_wr[1897]));
			radix2 #(.width(width)) rd_st4_1834  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1834]), .rdlo_in(a4_wr[1898]),  .coef_in(coef[672]), .rdup_out(a5_wr[1834]), .rdlo_out(a5_wr[1898]));
			radix2 #(.width(width)) rd_st4_1835  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1835]), .rdlo_in(a4_wr[1899]),  .coef_in(coef[688]), .rdup_out(a5_wr[1835]), .rdlo_out(a5_wr[1899]));
			radix2 #(.width(width)) rd_st4_1836  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1836]), .rdlo_in(a4_wr[1900]),  .coef_in(coef[704]), .rdup_out(a5_wr[1836]), .rdlo_out(a5_wr[1900]));
			radix2 #(.width(width)) rd_st4_1837  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1837]), .rdlo_in(a4_wr[1901]),  .coef_in(coef[720]), .rdup_out(a5_wr[1837]), .rdlo_out(a5_wr[1901]));
			radix2 #(.width(width)) rd_st4_1838  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1838]), .rdlo_in(a4_wr[1902]),  .coef_in(coef[736]), .rdup_out(a5_wr[1838]), .rdlo_out(a5_wr[1902]));
			radix2 #(.width(width)) rd_st4_1839  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1839]), .rdlo_in(a4_wr[1903]),  .coef_in(coef[752]), .rdup_out(a5_wr[1839]), .rdlo_out(a5_wr[1903]));
			radix2 #(.width(width)) rd_st4_1840  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1840]), .rdlo_in(a4_wr[1904]),  .coef_in(coef[768]), .rdup_out(a5_wr[1840]), .rdlo_out(a5_wr[1904]));
			radix2 #(.width(width)) rd_st4_1841  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1841]), .rdlo_in(a4_wr[1905]),  .coef_in(coef[784]), .rdup_out(a5_wr[1841]), .rdlo_out(a5_wr[1905]));
			radix2 #(.width(width)) rd_st4_1842  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1842]), .rdlo_in(a4_wr[1906]),  .coef_in(coef[800]), .rdup_out(a5_wr[1842]), .rdlo_out(a5_wr[1906]));
			radix2 #(.width(width)) rd_st4_1843  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1843]), .rdlo_in(a4_wr[1907]),  .coef_in(coef[816]), .rdup_out(a5_wr[1843]), .rdlo_out(a5_wr[1907]));
			radix2 #(.width(width)) rd_st4_1844  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1844]), .rdlo_in(a4_wr[1908]),  .coef_in(coef[832]), .rdup_out(a5_wr[1844]), .rdlo_out(a5_wr[1908]));
			radix2 #(.width(width)) rd_st4_1845  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1845]), .rdlo_in(a4_wr[1909]),  .coef_in(coef[848]), .rdup_out(a5_wr[1845]), .rdlo_out(a5_wr[1909]));
			radix2 #(.width(width)) rd_st4_1846  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1846]), .rdlo_in(a4_wr[1910]),  .coef_in(coef[864]), .rdup_out(a5_wr[1846]), .rdlo_out(a5_wr[1910]));
			radix2 #(.width(width)) rd_st4_1847  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1847]), .rdlo_in(a4_wr[1911]),  .coef_in(coef[880]), .rdup_out(a5_wr[1847]), .rdlo_out(a5_wr[1911]));
			radix2 #(.width(width)) rd_st4_1848  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1848]), .rdlo_in(a4_wr[1912]),  .coef_in(coef[896]), .rdup_out(a5_wr[1848]), .rdlo_out(a5_wr[1912]));
			radix2 #(.width(width)) rd_st4_1849  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1849]), .rdlo_in(a4_wr[1913]),  .coef_in(coef[912]), .rdup_out(a5_wr[1849]), .rdlo_out(a5_wr[1913]));
			radix2 #(.width(width)) rd_st4_1850  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1850]), .rdlo_in(a4_wr[1914]),  .coef_in(coef[928]), .rdup_out(a5_wr[1850]), .rdlo_out(a5_wr[1914]));
			radix2 #(.width(width)) rd_st4_1851  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1851]), .rdlo_in(a4_wr[1915]),  .coef_in(coef[944]), .rdup_out(a5_wr[1851]), .rdlo_out(a5_wr[1915]));
			radix2 #(.width(width)) rd_st4_1852  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1852]), .rdlo_in(a4_wr[1916]),  .coef_in(coef[960]), .rdup_out(a5_wr[1852]), .rdlo_out(a5_wr[1916]));
			radix2 #(.width(width)) rd_st4_1853  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1853]), .rdlo_in(a4_wr[1917]),  .coef_in(coef[976]), .rdup_out(a5_wr[1853]), .rdlo_out(a5_wr[1917]));
			radix2 #(.width(width)) rd_st4_1854  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1854]), .rdlo_in(a4_wr[1918]),  .coef_in(coef[992]), .rdup_out(a5_wr[1854]), .rdlo_out(a5_wr[1918]));
			radix2 #(.width(width)) rd_st4_1855  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1855]), .rdlo_in(a4_wr[1919]),  .coef_in(coef[1008]), .rdup_out(a5_wr[1855]), .rdlo_out(a5_wr[1919]));
			radix2 #(.width(width)) rd_st4_1920  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1920]), .rdlo_in(a4_wr[1984]),  .coef_in(coef[0]), .rdup_out(a5_wr[1920]), .rdlo_out(a5_wr[1984]));
			radix2 #(.width(width)) rd_st4_1921  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1921]), .rdlo_in(a4_wr[1985]),  .coef_in(coef[16]), .rdup_out(a5_wr[1921]), .rdlo_out(a5_wr[1985]));
			radix2 #(.width(width)) rd_st4_1922  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1922]), .rdlo_in(a4_wr[1986]),  .coef_in(coef[32]), .rdup_out(a5_wr[1922]), .rdlo_out(a5_wr[1986]));
			radix2 #(.width(width)) rd_st4_1923  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1923]), .rdlo_in(a4_wr[1987]),  .coef_in(coef[48]), .rdup_out(a5_wr[1923]), .rdlo_out(a5_wr[1987]));
			radix2 #(.width(width)) rd_st4_1924  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1924]), .rdlo_in(a4_wr[1988]),  .coef_in(coef[64]), .rdup_out(a5_wr[1924]), .rdlo_out(a5_wr[1988]));
			radix2 #(.width(width)) rd_st4_1925  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1925]), .rdlo_in(a4_wr[1989]),  .coef_in(coef[80]), .rdup_out(a5_wr[1925]), .rdlo_out(a5_wr[1989]));
			radix2 #(.width(width)) rd_st4_1926  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1926]), .rdlo_in(a4_wr[1990]),  .coef_in(coef[96]), .rdup_out(a5_wr[1926]), .rdlo_out(a5_wr[1990]));
			radix2 #(.width(width)) rd_st4_1927  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1927]), .rdlo_in(a4_wr[1991]),  .coef_in(coef[112]), .rdup_out(a5_wr[1927]), .rdlo_out(a5_wr[1991]));
			radix2 #(.width(width)) rd_st4_1928  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1928]), .rdlo_in(a4_wr[1992]),  .coef_in(coef[128]), .rdup_out(a5_wr[1928]), .rdlo_out(a5_wr[1992]));
			radix2 #(.width(width)) rd_st4_1929  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1929]), .rdlo_in(a4_wr[1993]),  .coef_in(coef[144]), .rdup_out(a5_wr[1929]), .rdlo_out(a5_wr[1993]));
			radix2 #(.width(width)) rd_st4_1930  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1930]), .rdlo_in(a4_wr[1994]),  .coef_in(coef[160]), .rdup_out(a5_wr[1930]), .rdlo_out(a5_wr[1994]));
			radix2 #(.width(width)) rd_st4_1931  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1931]), .rdlo_in(a4_wr[1995]),  .coef_in(coef[176]), .rdup_out(a5_wr[1931]), .rdlo_out(a5_wr[1995]));
			radix2 #(.width(width)) rd_st4_1932  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1932]), .rdlo_in(a4_wr[1996]),  .coef_in(coef[192]), .rdup_out(a5_wr[1932]), .rdlo_out(a5_wr[1996]));
			radix2 #(.width(width)) rd_st4_1933  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1933]), .rdlo_in(a4_wr[1997]),  .coef_in(coef[208]), .rdup_out(a5_wr[1933]), .rdlo_out(a5_wr[1997]));
			radix2 #(.width(width)) rd_st4_1934  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1934]), .rdlo_in(a4_wr[1998]),  .coef_in(coef[224]), .rdup_out(a5_wr[1934]), .rdlo_out(a5_wr[1998]));
			radix2 #(.width(width)) rd_st4_1935  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1935]), .rdlo_in(a4_wr[1999]),  .coef_in(coef[240]), .rdup_out(a5_wr[1935]), .rdlo_out(a5_wr[1999]));
			radix2 #(.width(width)) rd_st4_1936  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1936]), .rdlo_in(a4_wr[2000]),  .coef_in(coef[256]), .rdup_out(a5_wr[1936]), .rdlo_out(a5_wr[2000]));
			radix2 #(.width(width)) rd_st4_1937  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1937]), .rdlo_in(a4_wr[2001]),  .coef_in(coef[272]), .rdup_out(a5_wr[1937]), .rdlo_out(a5_wr[2001]));
			radix2 #(.width(width)) rd_st4_1938  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1938]), .rdlo_in(a4_wr[2002]),  .coef_in(coef[288]), .rdup_out(a5_wr[1938]), .rdlo_out(a5_wr[2002]));
			radix2 #(.width(width)) rd_st4_1939  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1939]), .rdlo_in(a4_wr[2003]),  .coef_in(coef[304]), .rdup_out(a5_wr[1939]), .rdlo_out(a5_wr[2003]));
			radix2 #(.width(width)) rd_st4_1940  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1940]), .rdlo_in(a4_wr[2004]),  .coef_in(coef[320]), .rdup_out(a5_wr[1940]), .rdlo_out(a5_wr[2004]));
			radix2 #(.width(width)) rd_st4_1941  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1941]), .rdlo_in(a4_wr[2005]),  .coef_in(coef[336]), .rdup_out(a5_wr[1941]), .rdlo_out(a5_wr[2005]));
			radix2 #(.width(width)) rd_st4_1942  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1942]), .rdlo_in(a4_wr[2006]),  .coef_in(coef[352]), .rdup_out(a5_wr[1942]), .rdlo_out(a5_wr[2006]));
			radix2 #(.width(width)) rd_st4_1943  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1943]), .rdlo_in(a4_wr[2007]),  .coef_in(coef[368]), .rdup_out(a5_wr[1943]), .rdlo_out(a5_wr[2007]));
			radix2 #(.width(width)) rd_st4_1944  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1944]), .rdlo_in(a4_wr[2008]),  .coef_in(coef[384]), .rdup_out(a5_wr[1944]), .rdlo_out(a5_wr[2008]));
			radix2 #(.width(width)) rd_st4_1945  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1945]), .rdlo_in(a4_wr[2009]),  .coef_in(coef[400]), .rdup_out(a5_wr[1945]), .rdlo_out(a5_wr[2009]));
			radix2 #(.width(width)) rd_st4_1946  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1946]), .rdlo_in(a4_wr[2010]),  .coef_in(coef[416]), .rdup_out(a5_wr[1946]), .rdlo_out(a5_wr[2010]));
			radix2 #(.width(width)) rd_st4_1947  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1947]), .rdlo_in(a4_wr[2011]),  .coef_in(coef[432]), .rdup_out(a5_wr[1947]), .rdlo_out(a5_wr[2011]));
			radix2 #(.width(width)) rd_st4_1948  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1948]), .rdlo_in(a4_wr[2012]),  .coef_in(coef[448]), .rdup_out(a5_wr[1948]), .rdlo_out(a5_wr[2012]));
			radix2 #(.width(width)) rd_st4_1949  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1949]), .rdlo_in(a4_wr[2013]),  .coef_in(coef[464]), .rdup_out(a5_wr[1949]), .rdlo_out(a5_wr[2013]));
			radix2 #(.width(width)) rd_st4_1950  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1950]), .rdlo_in(a4_wr[2014]),  .coef_in(coef[480]), .rdup_out(a5_wr[1950]), .rdlo_out(a5_wr[2014]));
			radix2 #(.width(width)) rd_st4_1951  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1951]), .rdlo_in(a4_wr[2015]),  .coef_in(coef[496]), .rdup_out(a5_wr[1951]), .rdlo_out(a5_wr[2015]));
			radix2 #(.width(width)) rd_st4_1952  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1952]), .rdlo_in(a4_wr[2016]),  .coef_in(coef[512]), .rdup_out(a5_wr[1952]), .rdlo_out(a5_wr[2016]));
			radix2 #(.width(width)) rd_st4_1953  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1953]), .rdlo_in(a4_wr[2017]),  .coef_in(coef[528]), .rdup_out(a5_wr[1953]), .rdlo_out(a5_wr[2017]));
			radix2 #(.width(width)) rd_st4_1954  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1954]), .rdlo_in(a4_wr[2018]),  .coef_in(coef[544]), .rdup_out(a5_wr[1954]), .rdlo_out(a5_wr[2018]));
			radix2 #(.width(width)) rd_st4_1955  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1955]), .rdlo_in(a4_wr[2019]),  .coef_in(coef[560]), .rdup_out(a5_wr[1955]), .rdlo_out(a5_wr[2019]));
			radix2 #(.width(width)) rd_st4_1956  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1956]), .rdlo_in(a4_wr[2020]),  .coef_in(coef[576]), .rdup_out(a5_wr[1956]), .rdlo_out(a5_wr[2020]));
			radix2 #(.width(width)) rd_st4_1957  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1957]), .rdlo_in(a4_wr[2021]),  .coef_in(coef[592]), .rdup_out(a5_wr[1957]), .rdlo_out(a5_wr[2021]));
			radix2 #(.width(width)) rd_st4_1958  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1958]), .rdlo_in(a4_wr[2022]),  .coef_in(coef[608]), .rdup_out(a5_wr[1958]), .rdlo_out(a5_wr[2022]));
			radix2 #(.width(width)) rd_st4_1959  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1959]), .rdlo_in(a4_wr[2023]),  .coef_in(coef[624]), .rdup_out(a5_wr[1959]), .rdlo_out(a5_wr[2023]));
			radix2 #(.width(width)) rd_st4_1960  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1960]), .rdlo_in(a4_wr[2024]),  .coef_in(coef[640]), .rdup_out(a5_wr[1960]), .rdlo_out(a5_wr[2024]));
			radix2 #(.width(width)) rd_st4_1961  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1961]), .rdlo_in(a4_wr[2025]),  .coef_in(coef[656]), .rdup_out(a5_wr[1961]), .rdlo_out(a5_wr[2025]));
			radix2 #(.width(width)) rd_st4_1962  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1962]), .rdlo_in(a4_wr[2026]),  .coef_in(coef[672]), .rdup_out(a5_wr[1962]), .rdlo_out(a5_wr[2026]));
			radix2 #(.width(width)) rd_st4_1963  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1963]), .rdlo_in(a4_wr[2027]),  .coef_in(coef[688]), .rdup_out(a5_wr[1963]), .rdlo_out(a5_wr[2027]));
			radix2 #(.width(width)) rd_st4_1964  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1964]), .rdlo_in(a4_wr[2028]),  .coef_in(coef[704]), .rdup_out(a5_wr[1964]), .rdlo_out(a5_wr[2028]));
			radix2 #(.width(width)) rd_st4_1965  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1965]), .rdlo_in(a4_wr[2029]),  .coef_in(coef[720]), .rdup_out(a5_wr[1965]), .rdlo_out(a5_wr[2029]));
			radix2 #(.width(width)) rd_st4_1966  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1966]), .rdlo_in(a4_wr[2030]),  .coef_in(coef[736]), .rdup_out(a5_wr[1966]), .rdlo_out(a5_wr[2030]));
			radix2 #(.width(width)) rd_st4_1967  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1967]), .rdlo_in(a4_wr[2031]),  .coef_in(coef[752]), .rdup_out(a5_wr[1967]), .rdlo_out(a5_wr[2031]));
			radix2 #(.width(width)) rd_st4_1968  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1968]), .rdlo_in(a4_wr[2032]),  .coef_in(coef[768]), .rdup_out(a5_wr[1968]), .rdlo_out(a5_wr[2032]));
			radix2 #(.width(width)) rd_st4_1969  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1969]), .rdlo_in(a4_wr[2033]),  .coef_in(coef[784]), .rdup_out(a5_wr[1969]), .rdlo_out(a5_wr[2033]));
			radix2 #(.width(width)) rd_st4_1970  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1970]), .rdlo_in(a4_wr[2034]),  .coef_in(coef[800]), .rdup_out(a5_wr[1970]), .rdlo_out(a5_wr[2034]));
			radix2 #(.width(width)) rd_st4_1971  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1971]), .rdlo_in(a4_wr[2035]),  .coef_in(coef[816]), .rdup_out(a5_wr[1971]), .rdlo_out(a5_wr[2035]));
			radix2 #(.width(width)) rd_st4_1972  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1972]), .rdlo_in(a4_wr[2036]),  .coef_in(coef[832]), .rdup_out(a5_wr[1972]), .rdlo_out(a5_wr[2036]));
			radix2 #(.width(width)) rd_st4_1973  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1973]), .rdlo_in(a4_wr[2037]),  .coef_in(coef[848]), .rdup_out(a5_wr[1973]), .rdlo_out(a5_wr[2037]));
			radix2 #(.width(width)) rd_st4_1974  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1974]), .rdlo_in(a4_wr[2038]),  .coef_in(coef[864]), .rdup_out(a5_wr[1974]), .rdlo_out(a5_wr[2038]));
			radix2 #(.width(width)) rd_st4_1975  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1975]), .rdlo_in(a4_wr[2039]),  .coef_in(coef[880]), .rdup_out(a5_wr[1975]), .rdlo_out(a5_wr[2039]));
			radix2 #(.width(width)) rd_st4_1976  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1976]), .rdlo_in(a4_wr[2040]),  .coef_in(coef[896]), .rdup_out(a5_wr[1976]), .rdlo_out(a5_wr[2040]));
			radix2 #(.width(width)) rd_st4_1977  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1977]), .rdlo_in(a4_wr[2041]),  .coef_in(coef[912]), .rdup_out(a5_wr[1977]), .rdlo_out(a5_wr[2041]));
			radix2 #(.width(width)) rd_st4_1978  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1978]), .rdlo_in(a4_wr[2042]),  .coef_in(coef[928]), .rdup_out(a5_wr[1978]), .rdlo_out(a5_wr[2042]));
			radix2 #(.width(width)) rd_st4_1979  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1979]), .rdlo_in(a4_wr[2043]),  .coef_in(coef[944]), .rdup_out(a5_wr[1979]), .rdlo_out(a5_wr[2043]));
			radix2 #(.width(width)) rd_st4_1980  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1980]), .rdlo_in(a4_wr[2044]),  .coef_in(coef[960]), .rdup_out(a5_wr[1980]), .rdlo_out(a5_wr[2044]));
			radix2 #(.width(width)) rd_st4_1981  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1981]), .rdlo_in(a4_wr[2045]),  .coef_in(coef[976]), .rdup_out(a5_wr[1981]), .rdlo_out(a5_wr[2045]));
			radix2 #(.width(width)) rd_st4_1982  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1982]), .rdlo_in(a4_wr[2046]),  .coef_in(coef[992]), .rdup_out(a5_wr[1982]), .rdlo_out(a5_wr[2046]));
			radix2 #(.width(width)) rd_st4_1983  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a4_wr[1983]), .rdlo_in(a4_wr[2047]),  .coef_in(coef[1008]), .rdup_out(a5_wr[1983]), .rdlo_out(a5_wr[2047]));

		//--- radix stage 5
			radix2 #(.width(width)) rd_st5_0   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[0]), .rdlo_in(a5_wr[32]),  .coef_in(coef[0]), .rdup_out(a6_wr[0]), .rdlo_out(a6_wr[32]));
			radix2 #(.width(width)) rd_st5_1   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1]), .rdlo_in(a5_wr[33]),  .coef_in(coef[32]), .rdup_out(a6_wr[1]), .rdlo_out(a6_wr[33]));
			radix2 #(.width(width)) rd_st5_2   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[2]), .rdlo_in(a5_wr[34]),  .coef_in(coef[64]), .rdup_out(a6_wr[2]), .rdlo_out(a6_wr[34]));
			radix2 #(.width(width)) rd_st5_3   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[3]), .rdlo_in(a5_wr[35]),  .coef_in(coef[96]), .rdup_out(a6_wr[3]), .rdlo_out(a6_wr[35]));
			radix2 #(.width(width)) rd_st5_4   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[4]), .rdlo_in(a5_wr[36]),  .coef_in(coef[128]), .rdup_out(a6_wr[4]), .rdlo_out(a6_wr[36]));
			radix2 #(.width(width)) rd_st5_5   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[5]), .rdlo_in(a5_wr[37]),  .coef_in(coef[160]), .rdup_out(a6_wr[5]), .rdlo_out(a6_wr[37]));
			radix2 #(.width(width)) rd_st5_6   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[6]), .rdlo_in(a5_wr[38]),  .coef_in(coef[192]), .rdup_out(a6_wr[6]), .rdlo_out(a6_wr[38]));
			radix2 #(.width(width)) rd_st5_7   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[7]), .rdlo_in(a5_wr[39]),  .coef_in(coef[224]), .rdup_out(a6_wr[7]), .rdlo_out(a6_wr[39]));
			radix2 #(.width(width)) rd_st5_8   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[8]), .rdlo_in(a5_wr[40]),  .coef_in(coef[256]), .rdup_out(a6_wr[8]), .rdlo_out(a6_wr[40]));
			radix2 #(.width(width)) rd_st5_9   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[9]), .rdlo_in(a5_wr[41]),  .coef_in(coef[288]), .rdup_out(a6_wr[9]), .rdlo_out(a6_wr[41]));
			radix2 #(.width(width)) rd_st5_10  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[10]), .rdlo_in(a5_wr[42]),  .coef_in(coef[320]), .rdup_out(a6_wr[10]), .rdlo_out(a6_wr[42]));
			radix2 #(.width(width)) rd_st5_11  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[11]), .rdlo_in(a5_wr[43]),  .coef_in(coef[352]), .rdup_out(a6_wr[11]), .rdlo_out(a6_wr[43]));
			radix2 #(.width(width)) rd_st5_12  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[12]), .rdlo_in(a5_wr[44]),  .coef_in(coef[384]), .rdup_out(a6_wr[12]), .rdlo_out(a6_wr[44]));
			radix2 #(.width(width)) rd_st5_13  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[13]), .rdlo_in(a5_wr[45]),  .coef_in(coef[416]), .rdup_out(a6_wr[13]), .rdlo_out(a6_wr[45]));
			radix2 #(.width(width)) rd_st5_14  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[14]), .rdlo_in(a5_wr[46]),  .coef_in(coef[448]), .rdup_out(a6_wr[14]), .rdlo_out(a6_wr[46]));
			radix2 #(.width(width)) rd_st5_15  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[15]), .rdlo_in(a5_wr[47]),  .coef_in(coef[480]), .rdup_out(a6_wr[15]), .rdlo_out(a6_wr[47]));
			radix2 #(.width(width)) rd_st5_16  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[16]), .rdlo_in(a5_wr[48]),  .coef_in(coef[512]), .rdup_out(a6_wr[16]), .rdlo_out(a6_wr[48]));
			radix2 #(.width(width)) rd_st5_17  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[17]), .rdlo_in(a5_wr[49]),  .coef_in(coef[544]), .rdup_out(a6_wr[17]), .rdlo_out(a6_wr[49]));
			radix2 #(.width(width)) rd_st5_18  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[18]), .rdlo_in(a5_wr[50]),  .coef_in(coef[576]), .rdup_out(a6_wr[18]), .rdlo_out(a6_wr[50]));
			radix2 #(.width(width)) rd_st5_19  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[19]), .rdlo_in(a5_wr[51]),  .coef_in(coef[608]), .rdup_out(a6_wr[19]), .rdlo_out(a6_wr[51]));
			radix2 #(.width(width)) rd_st5_20  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[20]), .rdlo_in(a5_wr[52]),  .coef_in(coef[640]), .rdup_out(a6_wr[20]), .rdlo_out(a6_wr[52]));
			radix2 #(.width(width)) rd_st5_21  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[21]), .rdlo_in(a5_wr[53]),  .coef_in(coef[672]), .rdup_out(a6_wr[21]), .rdlo_out(a6_wr[53]));
			radix2 #(.width(width)) rd_st5_22  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[22]), .rdlo_in(a5_wr[54]),  .coef_in(coef[704]), .rdup_out(a6_wr[22]), .rdlo_out(a6_wr[54]));
			radix2 #(.width(width)) rd_st5_23  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[23]), .rdlo_in(a5_wr[55]),  .coef_in(coef[736]), .rdup_out(a6_wr[23]), .rdlo_out(a6_wr[55]));
			radix2 #(.width(width)) rd_st5_24  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[24]), .rdlo_in(a5_wr[56]),  .coef_in(coef[768]), .rdup_out(a6_wr[24]), .rdlo_out(a6_wr[56]));
			radix2 #(.width(width)) rd_st5_25  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[25]), .rdlo_in(a5_wr[57]),  .coef_in(coef[800]), .rdup_out(a6_wr[25]), .rdlo_out(a6_wr[57]));
			radix2 #(.width(width)) rd_st5_26  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[26]), .rdlo_in(a5_wr[58]),  .coef_in(coef[832]), .rdup_out(a6_wr[26]), .rdlo_out(a6_wr[58]));
			radix2 #(.width(width)) rd_st5_27  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[27]), .rdlo_in(a5_wr[59]),  .coef_in(coef[864]), .rdup_out(a6_wr[27]), .rdlo_out(a6_wr[59]));
			radix2 #(.width(width)) rd_st5_28  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[28]), .rdlo_in(a5_wr[60]),  .coef_in(coef[896]), .rdup_out(a6_wr[28]), .rdlo_out(a6_wr[60]));
			radix2 #(.width(width)) rd_st5_29  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[29]), .rdlo_in(a5_wr[61]),  .coef_in(coef[928]), .rdup_out(a6_wr[29]), .rdlo_out(a6_wr[61]));
			radix2 #(.width(width)) rd_st5_30  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[30]), .rdlo_in(a5_wr[62]),  .coef_in(coef[960]), .rdup_out(a6_wr[30]), .rdlo_out(a6_wr[62]));
			radix2 #(.width(width)) rd_st5_31  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[31]), .rdlo_in(a5_wr[63]),  .coef_in(coef[992]), .rdup_out(a6_wr[31]), .rdlo_out(a6_wr[63]));
			radix2 #(.width(width)) rd_st5_64  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[64]), .rdlo_in(a5_wr[96]),  .coef_in(coef[0]), .rdup_out(a6_wr[64]), .rdlo_out(a6_wr[96]));
			radix2 #(.width(width)) rd_st5_65  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[65]), .rdlo_in(a5_wr[97]),  .coef_in(coef[32]), .rdup_out(a6_wr[65]), .rdlo_out(a6_wr[97]));
			radix2 #(.width(width)) rd_st5_66  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[66]), .rdlo_in(a5_wr[98]),  .coef_in(coef[64]), .rdup_out(a6_wr[66]), .rdlo_out(a6_wr[98]));
			radix2 #(.width(width)) rd_st5_67  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[67]), .rdlo_in(a5_wr[99]),  .coef_in(coef[96]), .rdup_out(a6_wr[67]), .rdlo_out(a6_wr[99]));
			radix2 #(.width(width)) rd_st5_68  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[68]), .rdlo_in(a5_wr[100]),  .coef_in(coef[128]), .rdup_out(a6_wr[68]), .rdlo_out(a6_wr[100]));
			radix2 #(.width(width)) rd_st5_69  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[69]), .rdlo_in(a5_wr[101]),  .coef_in(coef[160]), .rdup_out(a6_wr[69]), .rdlo_out(a6_wr[101]));
			radix2 #(.width(width)) rd_st5_70  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[70]), .rdlo_in(a5_wr[102]),  .coef_in(coef[192]), .rdup_out(a6_wr[70]), .rdlo_out(a6_wr[102]));
			radix2 #(.width(width)) rd_st5_71  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[71]), .rdlo_in(a5_wr[103]),  .coef_in(coef[224]), .rdup_out(a6_wr[71]), .rdlo_out(a6_wr[103]));
			radix2 #(.width(width)) rd_st5_72  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[72]), .rdlo_in(a5_wr[104]),  .coef_in(coef[256]), .rdup_out(a6_wr[72]), .rdlo_out(a6_wr[104]));
			radix2 #(.width(width)) rd_st5_73  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[73]), .rdlo_in(a5_wr[105]),  .coef_in(coef[288]), .rdup_out(a6_wr[73]), .rdlo_out(a6_wr[105]));
			radix2 #(.width(width)) rd_st5_74  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[74]), .rdlo_in(a5_wr[106]),  .coef_in(coef[320]), .rdup_out(a6_wr[74]), .rdlo_out(a6_wr[106]));
			radix2 #(.width(width)) rd_st5_75  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[75]), .rdlo_in(a5_wr[107]),  .coef_in(coef[352]), .rdup_out(a6_wr[75]), .rdlo_out(a6_wr[107]));
			radix2 #(.width(width)) rd_st5_76  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[76]), .rdlo_in(a5_wr[108]),  .coef_in(coef[384]), .rdup_out(a6_wr[76]), .rdlo_out(a6_wr[108]));
			radix2 #(.width(width)) rd_st5_77  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[77]), .rdlo_in(a5_wr[109]),  .coef_in(coef[416]), .rdup_out(a6_wr[77]), .rdlo_out(a6_wr[109]));
			radix2 #(.width(width)) rd_st5_78  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[78]), .rdlo_in(a5_wr[110]),  .coef_in(coef[448]), .rdup_out(a6_wr[78]), .rdlo_out(a6_wr[110]));
			radix2 #(.width(width)) rd_st5_79  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[79]), .rdlo_in(a5_wr[111]),  .coef_in(coef[480]), .rdup_out(a6_wr[79]), .rdlo_out(a6_wr[111]));
			radix2 #(.width(width)) rd_st5_80  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[80]), .rdlo_in(a5_wr[112]),  .coef_in(coef[512]), .rdup_out(a6_wr[80]), .rdlo_out(a6_wr[112]));
			radix2 #(.width(width)) rd_st5_81  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[81]), .rdlo_in(a5_wr[113]),  .coef_in(coef[544]), .rdup_out(a6_wr[81]), .rdlo_out(a6_wr[113]));
			radix2 #(.width(width)) rd_st5_82  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[82]), .rdlo_in(a5_wr[114]),  .coef_in(coef[576]), .rdup_out(a6_wr[82]), .rdlo_out(a6_wr[114]));
			radix2 #(.width(width)) rd_st5_83  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[83]), .rdlo_in(a5_wr[115]),  .coef_in(coef[608]), .rdup_out(a6_wr[83]), .rdlo_out(a6_wr[115]));
			radix2 #(.width(width)) rd_st5_84  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[84]), .rdlo_in(a5_wr[116]),  .coef_in(coef[640]), .rdup_out(a6_wr[84]), .rdlo_out(a6_wr[116]));
			radix2 #(.width(width)) rd_st5_85  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[85]), .rdlo_in(a5_wr[117]),  .coef_in(coef[672]), .rdup_out(a6_wr[85]), .rdlo_out(a6_wr[117]));
			radix2 #(.width(width)) rd_st5_86  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[86]), .rdlo_in(a5_wr[118]),  .coef_in(coef[704]), .rdup_out(a6_wr[86]), .rdlo_out(a6_wr[118]));
			radix2 #(.width(width)) rd_st5_87  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[87]), .rdlo_in(a5_wr[119]),  .coef_in(coef[736]), .rdup_out(a6_wr[87]), .rdlo_out(a6_wr[119]));
			radix2 #(.width(width)) rd_st5_88  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[88]), .rdlo_in(a5_wr[120]),  .coef_in(coef[768]), .rdup_out(a6_wr[88]), .rdlo_out(a6_wr[120]));
			radix2 #(.width(width)) rd_st5_89  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[89]), .rdlo_in(a5_wr[121]),  .coef_in(coef[800]), .rdup_out(a6_wr[89]), .rdlo_out(a6_wr[121]));
			radix2 #(.width(width)) rd_st5_90  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[90]), .rdlo_in(a5_wr[122]),  .coef_in(coef[832]), .rdup_out(a6_wr[90]), .rdlo_out(a6_wr[122]));
			radix2 #(.width(width)) rd_st5_91  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[91]), .rdlo_in(a5_wr[123]),  .coef_in(coef[864]), .rdup_out(a6_wr[91]), .rdlo_out(a6_wr[123]));
			radix2 #(.width(width)) rd_st5_92  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[92]), .rdlo_in(a5_wr[124]),  .coef_in(coef[896]), .rdup_out(a6_wr[92]), .rdlo_out(a6_wr[124]));
			radix2 #(.width(width)) rd_st5_93  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[93]), .rdlo_in(a5_wr[125]),  .coef_in(coef[928]), .rdup_out(a6_wr[93]), .rdlo_out(a6_wr[125]));
			radix2 #(.width(width)) rd_st5_94  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[94]), .rdlo_in(a5_wr[126]),  .coef_in(coef[960]), .rdup_out(a6_wr[94]), .rdlo_out(a6_wr[126]));
			radix2 #(.width(width)) rd_st5_95  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[95]), .rdlo_in(a5_wr[127]),  .coef_in(coef[992]), .rdup_out(a6_wr[95]), .rdlo_out(a6_wr[127]));
			radix2 #(.width(width)) rd_st5_128  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[128]), .rdlo_in(a5_wr[160]),  .coef_in(coef[0]), .rdup_out(a6_wr[128]), .rdlo_out(a6_wr[160]));
			radix2 #(.width(width)) rd_st5_129  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[129]), .rdlo_in(a5_wr[161]),  .coef_in(coef[32]), .rdup_out(a6_wr[129]), .rdlo_out(a6_wr[161]));
			radix2 #(.width(width)) rd_st5_130  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[130]), .rdlo_in(a5_wr[162]),  .coef_in(coef[64]), .rdup_out(a6_wr[130]), .rdlo_out(a6_wr[162]));
			radix2 #(.width(width)) rd_st5_131  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[131]), .rdlo_in(a5_wr[163]),  .coef_in(coef[96]), .rdup_out(a6_wr[131]), .rdlo_out(a6_wr[163]));
			radix2 #(.width(width)) rd_st5_132  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[132]), .rdlo_in(a5_wr[164]),  .coef_in(coef[128]), .rdup_out(a6_wr[132]), .rdlo_out(a6_wr[164]));
			radix2 #(.width(width)) rd_st5_133  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[133]), .rdlo_in(a5_wr[165]),  .coef_in(coef[160]), .rdup_out(a6_wr[133]), .rdlo_out(a6_wr[165]));
			radix2 #(.width(width)) rd_st5_134  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[134]), .rdlo_in(a5_wr[166]),  .coef_in(coef[192]), .rdup_out(a6_wr[134]), .rdlo_out(a6_wr[166]));
			radix2 #(.width(width)) rd_st5_135  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[135]), .rdlo_in(a5_wr[167]),  .coef_in(coef[224]), .rdup_out(a6_wr[135]), .rdlo_out(a6_wr[167]));
			radix2 #(.width(width)) rd_st5_136  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[136]), .rdlo_in(a5_wr[168]),  .coef_in(coef[256]), .rdup_out(a6_wr[136]), .rdlo_out(a6_wr[168]));
			radix2 #(.width(width)) rd_st5_137  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[137]), .rdlo_in(a5_wr[169]),  .coef_in(coef[288]), .rdup_out(a6_wr[137]), .rdlo_out(a6_wr[169]));
			radix2 #(.width(width)) rd_st5_138  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[138]), .rdlo_in(a5_wr[170]),  .coef_in(coef[320]), .rdup_out(a6_wr[138]), .rdlo_out(a6_wr[170]));
			radix2 #(.width(width)) rd_st5_139  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[139]), .rdlo_in(a5_wr[171]),  .coef_in(coef[352]), .rdup_out(a6_wr[139]), .rdlo_out(a6_wr[171]));
			radix2 #(.width(width)) rd_st5_140  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[140]), .rdlo_in(a5_wr[172]),  .coef_in(coef[384]), .rdup_out(a6_wr[140]), .rdlo_out(a6_wr[172]));
			radix2 #(.width(width)) rd_st5_141  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[141]), .rdlo_in(a5_wr[173]),  .coef_in(coef[416]), .rdup_out(a6_wr[141]), .rdlo_out(a6_wr[173]));
			radix2 #(.width(width)) rd_st5_142  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[142]), .rdlo_in(a5_wr[174]),  .coef_in(coef[448]), .rdup_out(a6_wr[142]), .rdlo_out(a6_wr[174]));
			radix2 #(.width(width)) rd_st5_143  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[143]), .rdlo_in(a5_wr[175]),  .coef_in(coef[480]), .rdup_out(a6_wr[143]), .rdlo_out(a6_wr[175]));
			radix2 #(.width(width)) rd_st5_144  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[144]), .rdlo_in(a5_wr[176]),  .coef_in(coef[512]), .rdup_out(a6_wr[144]), .rdlo_out(a6_wr[176]));
			radix2 #(.width(width)) rd_st5_145  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[145]), .rdlo_in(a5_wr[177]),  .coef_in(coef[544]), .rdup_out(a6_wr[145]), .rdlo_out(a6_wr[177]));
			radix2 #(.width(width)) rd_st5_146  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[146]), .rdlo_in(a5_wr[178]),  .coef_in(coef[576]), .rdup_out(a6_wr[146]), .rdlo_out(a6_wr[178]));
			radix2 #(.width(width)) rd_st5_147  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[147]), .rdlo_in(a5_wr[179]),  .coef_in(coef[608]), .rdup_out(a6_wr[147]), .rdlo_out(a6_wr[179]));
			radix2 #(.width(width)) rd_st5_148  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[148]), .rdlo_in(a5_wr[180]),  .coef_in(coef[640]), .rdup_out(a6_wr[148]), .rdlo_out(a6_wr[180]));
			radix2 #(.width(width)) rd_st5_149  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[149]), .rdlo_in(a5_wr[181]),  .coef_in(coef[672]), .rdup_out(a6_wr[149]), .rdlo_out(a6_wr[181]));
			radix2 #(.width(width)) rd_st5_150  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[150]), .rdlo_in(a5_wr[182]),  .coef_in(coef[704]), .rdup_out(a6_wr[150]), .rdlo_out(a6_wr[182]));
			radix2 #(.width(width)) rd_st5_151  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[151]), .rdlo_in(a5_wr[183]),  .coef_in(coef[736]), .rdup_out(a6_wr[151]), .rdlo_out(a6_wr[183]));
			radix2 #(.width(width)) rd_st5_152  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[152]), .rdlo_in(a5_wr[184]),  .coef_in(coef[768]), .rdup_out(a6_wr[152]), .rdlo_out(a6_wr[184]));
			radix2 #(.width(width)) rd_st5_153  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[153]), .rdlo_in(a5_wr[185]),  .coef_in(coef[800]), .rdup_out(a6_wr[153]), .rdlo_out(a6_wr[185]));
			radix2 #(.width(width)) rd_st5_154  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[154]), .rdlo_in(a5_wr[186]),  .coef_in(coef[832]), .rdup_out(a6_wr[154]), .rdlo_out(a6_wr[186]));
			radix2 #(.width(width)) rd_st5_155  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[155]), .rdlo_in(a5_wr[187]),  .coef_in(coef[864]), .rdup_out(a6_wr[155]), .rdlo_out(a6_wr[187]));
			radix2 #(.width(width)) rd_st5_156  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[156]), .rdlo_in(a5_wr[188]),  .coef_in(coef[896]), .rdup_out(a6_wr[156]), .rdlo_out(a6_wr[188]));
			radix2 #(.width(width)) rd_st5_157  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[157]), .rdlo_in(a5_wr[189]),  .coef_in(coef[928]), .rdup_out(a6_wr[157]), .rdlo_out(a6_wr[189]));
			radix2 #(.width(width)) rd_st5_158  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[158]), .rdlo_in(a5_wr[190]),  .coef_in(coef[960]), .rdup_out(a6_wr[158]), .rdlo_out(a6_wr[190]));
			radix2 #(.width(width)) rd_st5_159  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[159]), .rdlo_in(a5_wr[191]),  .coef_in(coef[992]), .rdup_out(a6_wr[159]), .rdlo_out(a6_wr[191]));
			radix2 #(.width(width)) rd_st5_192  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[192]), .rdlo_in(a5_wr[224]),  .coef_in(coef[0]), .rdup_out(a6_wr[192]), .rdlo_out(a6_wr[224]));
			radix2 #(.width(width)) rd_st5_193  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[193]), .rdlo_in(a5_wr[225]),  .coef_in(coef[32]), .rdup_out(a6_wr[193]), .rdlo_out(a6_wr[225]));
			radix2 #(.width(width)) rd_st5_194  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[194]), .rdlo_in(a5_wr[226]),  .coef_in(coef[64]), .rdup_out(a6_wr[194]), .rdlo_out(a6_wr[226]));
			radix2 #(.width(width)) rd_st5_195  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[195]), .rdlo_in(a5_wr[227]),  .coef_in(coef[96]), .rdup_out(a6_wr[195]), .rdlo_out(a6_wr[227]));
			radix2 #(.width(width)) rd_st5_196  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[196]), .rdlo_in(a5_wr[228]),  .coef_in(coef[128]), .rdup_out(a6_wr[196]), .rdlo_out(a6_wr[228]));
			radix2 #(.width(width)) rd_st5_197  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[197]), .rdlo_in(a5_wr[229]),  .coef_in(coef[160]), .rdup_out(a6_wr[197]), .rdlo_out(a6_wr[229]));
			radix2 #(.width(width)) rd_st5_198  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[198]), .rdlo_in(a5_wr[230]),  .coef_in(coef[192]), .rdup_out(a6_wr[198]), .rdlo_out(a6_wr[230]));
			radix2 #(.width(width)) rd_st5_199  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[199]), .rdlo_in(a5_wr[231]),  .coef_in(coef[224]), .rdup_out(a6_wr[199]), .rdlo_out(a6_wr[231]));
			radix2 #(.width(width)) rd_st5_200  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[200]), .rdlo_in(a5_wr[232]),  .coef_in(coef[256]), .rdup_out(a6_wr[200]), .rdlo_out(a6_wr[232]));
			radix2 #(.width(width)) rd_st5_201  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[201]), .rdlo_in(a5_wr[233]),  .coef_in(coef[288]), .rdup_out(a6_wr[201]), .rdlo_out(a6_wr[233]));
			radix2 #(.width(width)) rd_st5_202  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[202]), .rdlo_in(a5_wr[234]),  .coef_in(coef[320]), .rdup_out(a6_wr[202]), .rdlo_out(a6_wr[234]));
			radix2 #(.width(width)) rd_st5_203  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[203]), .rdlo_in(a5_wr[235]),  .coef_in(coef[352]), .rdup_out(a6_wr[203]), .rdlo_out(a6_wr[235]));
			radix2 #(.width(width)) rd_st5_204  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[204]), .rdlo_in(a5_wr[236]),  .coef_in(coef[384]), .rdup_out(a6_wr[204]), .rdlo_out(a6_wr[236]));
			radix2 #(.width(width)) rd_st5_205  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[205]), .rdlo_in(a5_wr[237]),  .coef_in(coef[416]), .rdup_out(a6_wr[205]), .rdlo_out(a6_wr[237]));
			radix2 #(.width(width)) rd_st5_206  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[206]), .rdlo_in(a5_wr[238]),  .coef_in(coef[448]), .rdup_out(a6_wr[206]), .rdlo_out(a6_wr[238]));
			radix2 #(.width(width)) rd_st5_207  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[207]), .rdlo_in(a5_wr[239]),  .coef_in(coef[480]), .rdup_out(a6_wr[207]), .rdlo_out(a6_wr[239]));
			radix2 #(.width(width)) rd_st5_208  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[208]), .rdlo_in(a5_wr[240]),  .coef_in(coef[512]), .rdup_out(a6_wr[208]), .rdlo_out(a6_wr[240]));
			radix2 #(.width(width)) rd_st5_209  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[209]), .rdlo_in(a5_wr[241]),  .coef_in(coef[544]), .rdup_out(a6_wr[209]), .rdlo_out(a6_wr[241]));
			radix2 #(.width(width)) rd_st5_210  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[210]), .rdlo_in(a5_wr[242]),  .coef_in(coef[576]), .rdup_out(a6_wr[210]), .rdlo_out(a6_wr[242]));
			radix2 #(.width(width)) rd_st5_211  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[211]), .rdlo_in(a5_wr[243]),  .coef_in(coef[608]), .rdup_out(a6_wr[211]), .rdlo_out(a6_wr[243]));
			radix2 #(.width(width)) rd_st5_212  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[212]), .rdlo_in(a5_wr[244]),  .coef_in(coef[640]), .rdup_out(a6_wr[212]), .rdlo_out(a6_wr[244]));
			radix2 #(.width(width)) rd_st5_213  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[213]), .rdlo_in(a5_wr[245]),  .coef_in(coef[672]), .rdup_out(a6_wr[213]), .rdlo_out(a6_wr[245]));
			radix2 #(.width(width)) rd_st5_214  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[214]), .rdlo_in(a5_wr[246]),  .coef_in(coef[704]), .rdup_out(a6_wr[214]), .rdlo_out(a6_wr[246]));
			radix2 #(.width(width)) rd_st5_215  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[215]), .rdlo_in(a5_wr[247]),  .coef_in(coef[736]), .rdup_out(a6_wr[215]), .rdlo_out(a6_wr[247]));
			radix2 #(.width(width)) rd_st5_216  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[216]), .rdlo_in(a5_wr[248]),  .coef_in(coef[768]), .rdup_out(a6_wr[216]), .rdlo_out(a6_wr[248]));
			radix2 #(.width(width)) rd_st5_217  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[217]), .rdlo_in(a5_wr[249]),  .coef_in(coef[800]), .rdup_out(a6_wr[217]), .rdlo_out(a6_wr[249]));
			radix2 #(.width(width)) rd_st5_218  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[218]), .rdlo_in(a5_wr[250]),  .coef_in(coef[832]), .rdup_out(a6_wr[218]), .rdlo_out(a6_wr[250]));
			radix2 #(.width(width)) rd_st5_219  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[219]), .rdlo_in(a5_wr[251]),  .coef_in(coef[864]), .rdup_out(a6_wr[219]), .rdlo_out(a6_wr[251]));
			radix2 #(.width(width)) rd_st5_220  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[220]), .rdlo_in(a5_wr[252]),  .coef_in(coef[896]), .rdup_out(a6_wr[220]), .rdlo_out(a6_wr[252]));
			radix2 #(.width(width)) rd_st5_221  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[221]), .rdlo_in(a5_wr[253]),  .coef_in(coef[928]), .rdup_out(a6_wr[221]), .rdlo_out(a6_wr[253]));
			radix2 #(.width(width)) rd_st5_222  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[222]), .rdlo_in(a5_wr[254]),  .coef_in(coef[960]), .rdup_out(a6_wr[222]), .rdlo_out(a6_wr[254]));
			radix2 #(.width(width)) rd_st5_223  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[223]), .rdlo_in(a5_wr[255]),  .coef_in(coef[992]), .rdup_out(a6_wr[223]), .rdlo_out(a6_wr[255]));
			radix2 #(.width(width)) rd_st5_256  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[256]), .rdlo_in(a5_wr[288]),  .coef_in(coef[0]), .rdup_out(a6_wr[256]), .rdlo_out(a6_wr[288]));
			radix2 #(.width(width)) rd_st5_257  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[257]), .rdlo_in(a5_wr[289]),  .coef_in(coef[32]), .rdup_out(a6_wr[257]), .rdlo_out(a6_wr[289]));
			radix2 #(.width(width)) rd_st5_258  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[258]), .rdlo_in(a5_wr[290]),  .coef_in(coef[64]), .rdup_out(a6_wr[258]), .rdlo_out(a6_wr[290]));
			radix2 #(.width(width)) rd_st5_259  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[259]), .rdlo_in(a5_wr[291]),  .coef_in(coef[96]), .rdup_out(a6_wr[259]), .rdlo_out(a6_wr[291]));
			radix2 #(.width(width)) rd_st5_260  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[260]), .rdlo_in(a5_wr[292]),  .coef_in(coef[128]), .rdup_out(a6_wr[260]), .rdlo_out(a6_wr[292]));
			radix2 #(.width(width)) rd_st5_261  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[261]), .rdlo_in(a5_wr[293]),  .coef_in(coef[160]), .rdup_out(a6_wr[261]), .rdlo_out(a6_wr[293]));
			radix2 #(.width(width)) rd_st5_262  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[262]), .rdlo_in(a5_wr[294]),  .coef_in(coef[192]), .rdup_out(a6_wr[262]), .rdlo_out(a6_wr[294]));
			radix2 #(.width(width)) rd_st5_263  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[263]), .rdlo_in(a5_wr[295]),  .coef_in(coef[224]), .rdup_out(a6_wr[263]), .rdlo_out(a6_wr[295]));
			radix2 #(.width(width)) rd_st5_264  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[264]), .rdlo_in(a5_wr[296]),  .coef_in(coef[256]), .rdup_out(a6_wr[264]), .rdlo_out(a6_wr[296]));
			radix2 #(.width(width)) rd_st5_265  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[265]), .rdlo_in(a5_wr[297]),  .coef_in(coef[288]), .rdup_out(a6_wr[265]), .rdlo_out(a6_wr[297]));
			radix2 #(.width(width)) rd_st5_266  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[266]), .rdlo_in(a5_wr[298]),  .coef_in(coef[320]), .rdup_out(a6_wr[266]), .rdlo_out(a6_wr[298]));
			radix2 #(.width(width)) rd_st5_267  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[267]), .rdlo_in(a5_wr[299]),  .coef_in(coef[352]), .rdup_out(a6_wr[267]), .rdlo_out(a6_wr[299]));
			radix2 #(.width(width)) rd_st5_268  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[268]), .rdlo_in(a5_wr[300]),  .coef_in(coef[384]), .rdup_out(a6_wr[268]), .rdlo_out(a6_wr[300]));
			radix2 #(.width(width)) rd_st5_269  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[269]), .rdlo_in(a5_wr[301]),  .coef_in(coef[416]), .rdup_out(a6_wr[269]), .rdlo_out(a6_wr[301]));
			radix2 #(.width(width)) rd_st5_270  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[270]), .rdlo_in(a5_wr[302]),  .coef_in(coef[448]), .rdup_out(a6_wr[270]), .rdlo_out(a6_wr[302]));
			radix2 #(.width(width)) rd_st5_271  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[271]), .rdlo_in(a5_wr[303]),  .coef_in(coef[480]), .rdup_out(a6_wr[271]), .rdlo_out(a6_wr[303]));
			radix2 #(.width(width)) rd_st5_272  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[272]), .rdlo_in(a5_wr[304]),  .coef_in(coef[512]), .rdup_out(a6_wr[272]), .rdlo_out(a6_wr[304]));
			radix2 #(.width(width)) rd_st5_273  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[273]), .rdlo_in(a5_wr[305]),  .coef_in(coef[544]), .rdup_out(a6_wr[273]), .rdlo_out(a6_wr[305]));
			radix2 #(.width(width)) rd_st5_274  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[274]), .rdlo_in(a5_wr[306]),  .coef_in(coef[576]), .rdup_out(a6_wr[274]), .rdlo_out(a6_wr[306]));
			radix2 #(.width(width)) rd_st5_275  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[275]), .rdlo_in(a5_wr[307]),  .coef_in(coef[608]), .rdup_out(a6_wr[275]), .rdlo_out(a6_wr[307]));
			radix2 #(.width(width)) rd_st5_276  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[276]), .rdlo_in(a5_wr[308]),  .coef_in(coef[640]), .rdup_out(a6_wr[276]), .rdlo_out(a6_wr[308]));
			radix2 #(.width(width)) rd_st5_277  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[277]), .rdlo_in(a5_wr[309]),  .coef_in(coef[672]), .rdup_out(a6_wr[277]), .rdlo_out(a6_wr[309]));
			radix2 #(.width(width)) rd_st5_278  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[278]), .rdlo_in(a5_wr[310]),  .coef_in(coef[704]), .rdup_out(a6_wr[278]), .rdlo_out(a6_wr[310]));
			radix2 #(.width(width)) rd_st5_279  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[279]), .rdlo_in(a5_wr[311]),  .coef_in(coef[736]), .rdup_out(a6_wr[279]), .rdlo_out(a6_wr[311]));
			radix2 #(.width(width)) rd_st5_280  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[280]), .rdlo_in(a5_wr[312]),  .coef_in(coef[768]), .rdup_out(a6_wr[280]), .rdlo_out(a6_wr[312]));
			radix2 #(.width(width)) rd_st5_281  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[281]), .rdlo_in(a5_wr[313]),  .coef_in(coef[800]), .rdup_out(a6_wr[281]), .rdlo_out(a6_wr[313]));
			radix2 #(.width(width)) rd_st5_282  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[282]), .rdlo_in(a5_wr[314]),  .coef_in(coef[832]), .rdup_out(a6_wr[282]), .rdlo_out(a6_wr[314]));
			radix2 #(.width(width)) rd_st5_283  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[283]), .rdlo_in(a5_wr[315]),  .coef_in(coef[864]), .rdup_out(a6_wr[283]), .rdlo_out(a6_wr[315]));
			radix2 #(.width(width)) rd_st5_284  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[284]), .rdlo_in(a5_wr[316]),  .coef_in(coef[896]), .rdup_out(a6_wr[284]), .rdlo_out(a6_wr[316]));
			radix2 #(.width(width)) rd_st5_285  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[285]), .rdlo_in(a5_wr[317]),  .coef_in(coef[928]), .rdup_out(a6_wr[285]), .rdlo_out(a6_wr[317]));
			radix2 #(.width(width)) rd_st5_286  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[286]), .rdlo_in(a5_wr[318]),  .coef_in(coef[960]), .rdup_out(a6_wr[286]), .rdlo_out(a6_wr[318]));
			radix2 #(.width(width)) rd_st5_287  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[287]), .rdlo_in(a5_wr[319]),  .coef_in(coef[992]), .rdup_out(a6_wr[287]), .rdlo_out(a6_wr[319]));
			radix2 #(.width(width)) rd_st5_320  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[320]), .rdlo_in(a5_wr[352]),  .coef_in(coef[0]), .rdup_out(a6_wr[320]), .rdlo_out(a6_wr[352]));
			radix2 #(.width(width)) rd_st5_321  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[321]), .rdlo_in(a5_wr[353]),  .coef_in(coef[32]), .rdup_out(a6_wr[321]), .rdlo_out(a6_wr[353]));
			radix2 #(.width(width)) rd_st5_322  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[322]), .rdlo_in(a5_wr[354]),  .coef_in(coef[64]), .rdup_out(a6_wr[322]), .rdlo_out(a6_wr[354]));
			radix2 #(.width(width)) rd_st5_323  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[323]), .rdlo_in(a5_wr[355]),  .coef_in(coef[96]), .rdup_out(a6_wr[323]), .rdlo_out(a6_wr[355]));
			radix2 #(.width(width)) rd_st5_324  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[324]), .rdlo_in(a5_wr[356]),  .coef_in(coef[128]), .rdup_out(a6_wr[324]), .rdlo_out(a6_wr[356]));
			radix2 #(.width(width)) rd_st5_325  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[325]), .rdlo_in(a5_wr[357]),  .coef_in(coef[160]), .rdup_out(a6_wr[325]), .rdlo_out(a6_wr[357]));
			radix2 #(.width(width)) rd_st5_326  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[326]), .rdlo_in(a5_wr[358]),  .coef_in(coef[192]), .rdup_out(a6_wr[326]), .rdlo_out(a6_wr[358]));
			radix2 #(.width(width)) rd_st5_327  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[327]), .rdlo_in(a5_wr[359]),  .coef_in(coef[224]), .rdup_out(a6_wr[327]), .rdlo_out(a6_wr[359]));
			radix2 #(.width(width)) rd_st5_328  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[328]), .rdlo_in(a5_wr[360]),  .coef_in(coef[256]), .rdup_out(a6_wr[328]), .rdlo_out(a6_wr[360]));
			radix2 #(.width(width)) rd_st5_329  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[329]), .rdlo_in(a5_wr[361]),  .coef_in(coef[288]), .rdup_out(a6_wr[329]), .rdlo_out(a6_wr[361]));
			radix2 #(.width(width)) rd_st5_330  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[330]), .rdlo_in(a5_wr[362]),  .coef_in(coef[320]), .rdup_out(a6_wr[330]), .rdlo_out(a6_wr[362]));
			radix2 #(.width(width)) rd_st5_331  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[331]), .rdlo_in(a5_wr[363]),  .coef_in(coef[352]), .rdup_out(a6_wr[331]), .rdlo_out(a6_wr[363]));
			radix2 #(.width(width)) rd_st5_332  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[332]), .rdlo_in(a5_wr[364]),  .coef_in(coef[384]), .rdup_out(a6_wr[332]), .rdlo_out(a6_wr[364]));
			radix2 #(.width(width)) rd_st5_333  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[333]), .rdlo_in(a5_wr[365]),  .coef_in(coef[416]), .rdup_out(a6_wr[333]), .rdlo_out(a6_wr[365]));
			radix2 #(.width(width)) rd_st5_334  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[334]), .rdlo_in(a5_wr[366]),  .coef_in(coef[448]), .rdup_out(a6_wr[334]), .rdlo_out(a6_wr[366]));
			radix2 #(.width(width)) rd_st5_335  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[335]), .rdlo_in(a5_wr[367]),  .coef_in(coef[480]), .rdup_out(a6_wr[335]), .rdlo_out(a6_wr[367]));
			radix2 #(.width(width)) rd_st5_336  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[336]), .rdlo_in(a5_wr[368]),  .coef_in(coef[512]), .rdup_out(a6_wr[336]), .rdlo_out(a6_wr[368]));
			radix2 #(.width(width)) rd_st5_337  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[337]), .rdlo_in(a5_wr[369]),  .coef_in(coef[544]), .rdup_out(a6_wr[337]), .rdlo_out(a6_wr[369]));
			radix2 #(.width(width)) rd_st5_338  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[338]), .rdlo_in(a5_wr[370]),  .coef_in(coef[576]), .rdup_out(a6_wr[338]), .rdlo_out(a6_wr[370]));
			radix2 #(.width(width)) rd_st5_339  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[339]), .rdlo_in(a5_wr[371]),  .coef_in(coef[608]), .rdup_out(a6_wr[339]), .rdlo_out(a6_wr[371]));
			radix2 #(.width(width)) rd_st5_340  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[340]), .rdlo_in(a5_wr[372]),  .coef_in(coef[640]), .rdup_out(a6_wr[340]), .rdlo_out(a6_wr[372]));
			radix2 #(.width(width)) rd_st5_341  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[341]), .rdlo_in(a5_wr[373]),  .coef_in(coef[672]), .rdup_out(a6_wr[341]), .rdlo_out(a6_wr[373]));
			radix2 #(.width(width)) rd_st5_342  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[342]), .rdlo_in(a5_wr[374]),  .coef_in(coef[704]), .rdup_out(a6_wr[342]), .rdlo_out(a6_wr[374]));
			radix2 #(.width(width)) rd_st5_343  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[343]), .rdlo_in(a5_wr[375]),  .coef_in(coef[736]), .rdup_out(a6_wr[343]), .rdlo_out(a6_wr[375]));
			radix2 #(.width(width)) rd_st5_344  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[344]), .rdlo_in(a5_wr[376]),  .coef_in(coef[768]), .rdup_out(a6_wr[344]), .rdlo_out(a6_wr[376]));
			radix2 #(.width(width)) rd_st5_345  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[345]), .rdlo_in(a5_wr[377]),  .coef_in(coef[800]), .rdup_out(a6_wr[345]), .rdlo_out(a6_wr[377]));
			radix2 #(.width(width)) rd_st5_346  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[346]), .rdlo_in(a5_wr[378]),  .coef_in(coef[832]), .rdup_out(a6_wr[346]), .rdlo_out(a6_wr[378]));
			radix2 #(.width(width)) rd_st5_347  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[347]), .rdlo_in(a5_wr[379]),  .coef_in(coef[864]), .rdup_out(a6_wr[347]), .rdlo_out(a6_wr[379]));
			radix2 #(.width(width)) rd_st5_348  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[348]), .rdlo_in(a5_wr[380]),  .coef_in(coef[896]), .rdup_out(a6_wr[348]), .rdlo_out(a6_wr[380]));
			radix2 #(.width(width)) rd_st5_349  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[349]), .rdlo_in(a5_wr[381]),  .coef_in(coef[928]), .rdup_out(a6_wr[349]), .rdlo_out(a6_wr[381]));
			radix2 #(.width(width)) rd_st5_350  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[350]), .rdlo_in(a5_wr[382]),  .coef_in(coef[960]), .rdup_out(a6_wr[350]), .rdlo_out(a6_wr[382]));
			radix2 #(.width(width)) rd_st5_351  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[351]), .rdlo_in(a5_wr[383]),  .coef_in(coef[992]), .rdup_out(a6_wr[351]), .rdlo_out(a6_wr[383]));
			radix2 #(.width(width)) rd_st5_384  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[384]), .rdlo_in(a5_wr[416]),  .coef_in(coef[0]), .rdup_out(a6_wr[384]), .rdlo_out(a6_wr[416]));
			radix2 #(.width(width)) rd_st5_385  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[385]), .rdlo_in(a5_wr[417]),  .coef_in(coef[32]), .rdup_out(a6_wr[385]), .rdlo_out(a6_wr[417]));
			radix2 #(.width(width)) rd_st5_386  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[386]), .rdlo_in(a5_wr[418]),  .coef_in(coef[64]), .rdup_out(a6_wr[386]), .rdlo_out(a6_wr[418]));
			radix2 #(.width(width)) rd_st5_387  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[387]), .rdlo_in(a5_wr[419]),  .coef_in(coef[96]), .rdup_out(a6_wr[387]), .rdlo_out(a6_wr[419]));
			radix2 #(.width(width)) rd_st5_388  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[388]), .rdlo_in(a5_wr[420]),  .coef_in(coef[128]), .rdup_out(a6_wr[388]), .rdlo_out(a6_wr[420]));
			radix2 #(.width(width)) rd_st5_389  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[389]), .rdlo_in(a5_wr[421]),  .coef_in(coef[160]), .rdup_out(a6_wr[389]), .rdlo_out(a6_wr[421]));
			radix2 #(.width(width)) rd_st5_390  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[390]), .rdlo_in(a5_wr[422]),  .coef_in(coef[192]), .rdup_out(a6_wr[390]), .rdlo_out(a6_wr[422]));
			radix2 #(.width(width)) rd_st5_391  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[391]), .rdlo_in(a5_wr[423]),  .coef_in(coef[224]), .rdup_out(a6_wr[391]), .rdlo_out(a6_wr[423]));
			radix2 #(.width(width)) rd_st5_392  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[392]), .rdlo_in(a5_wr[424]),  .coef_in(coef[256]), .rdup_out(a6_wr[392]), .rdlo_out(a6_wr[424]));
			radix2 #(.width(width)) rd_st5_393  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[393]), .rdlo_in(a5_wr[425]),  .coef_in(coef[288]), .rdup_out(a6_wr[393]), .rdlo_out(a6_wr[425]));
			radix2 #(.width(width)) rd_st5_394  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[394]), .rdlo_in(a5_wr[426]),  .coef_in(coef[320]), .rdup_out(a6_wr[394]), .rdlo_out(a6_wr[426]));
			radix2 #(.width(width)) rd_st5_395  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[395]), .rdlo_in(a5_wr[427]),  .coef_in(coef[352]), .rdup_out(a6_wr[395]), .rdlo_out(a6_wr[427]));
			radix2 #(.width(width)) rd_st5_396  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[396]), .rdlo_in(a5_wr[428]),  .coef_in(coef[384]), .rdup_out(a6_wr[396]), .rdlo_out(a6_wr[428]));
			radix2 #(.width(width)) rd_st5_397  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[397]), .rdlo_in(a5_wr[429]),  .coef_in(coef[416]), .rdup_out(a6_wr[397]), .rdlo_out(a6_wr[429]));
			radix2 #(.width(width)) rd_st5_398  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[398]), .rdlo_in(a5_wr[430]),  .coef_in(coef[448]), .rdup_out(a6_wr[398]), .rdlo_out(a6_wr[430]));
			radix2 #(.width(width)) rd_st5_399  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[399]), .rdlo_in(a5_wr[431]),  .coef_in(coef[480]), .rdup_out(a6_wr[399]), .rdlo_out(a6_wr[431]));
			radix2 #(.width(width)) rd_st5_400  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[400]), .rdlo_in(a5_wr[432]),  .coef_in(coef[512]), .rdup_out(a6_wr[400]), .rdlo_out(a6_wr[432]));
			radix2 #(.width(width)) rd_st5_401  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[401]), .rdlo_in(a5_wr[433]),  .coef_in(coef[544]), .rdup_out(a6_wr[401]), .rdlo_out(a6_wr[433]));
			radix2 #(.width(width)) rd_st5_402  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[402]), .rdlo_in(a5_wr[434]),  .coef_in(coef[576]), .rdup_out(a6_wr[402]), .rdlo_out(a6_wr[434]));
			radix2 #(.width(width)) rd_st5_403  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[403]), .rdlo_in(a5_wr[435]),  .coef_in(coef[608]), .rdup_out(a6_wr[403]), .rdlo_out(a6_wr[435]));
			radix2 #(.width(width)) rd_st5_404  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[404]), .rdlo_in(a5_wr[436]),  .coef_in(coef[640]), .rdup_out(a6_wr[404]), .rdlo_out(a6_wr[436]));
			radix2 #(.width(width)) rd_st5_405  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[405]), .rdlo_in(a5_wr[437]),  .coef_in(coef[672]), .rdup_out(a6_wr[405]), .rdlo_out(a6_wr[437]));
			radix2 #(.width(width)) rd_st5_406  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[406]), .rdlo_in(a5_wr[438]),  .coef_in(coef[704]), .rdup_out(a6_wr[406]), .rdlo_out(a6_wr[438]));
			radix2 #(.width(width)) rd_st5_407  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[407]), .rdlo_in(a5_wr[439]),  .coef_in(coef[736]), .rdup_out(a6_wr[407]), .rdlo_out(a6_wr[439]));
			radix2 #(.width(width)) rd_st5_408  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[408]), .rdlo_in(a5_wr[440]),  .coef_in(coef[768]), .rdup_out(a6_wr[408]), .rdlo_out(a6_wr[440]));
			radix2 #(.width(width)) rd_st5_409  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[409]), .rdlo_in(a5_wr[441]),  .coef_in(coef[800]), .rdup_out(a6_wr[409]), .rdlo_out(a6_wr[441]));
			radix2 #(.width(width)) rd_st5_410  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[410]), .rdlo_in(a5_wr[442]),  .coef_in(coef[832]), .rdup_out(a6_wr[410]), .rdlo_out(a6_wr[442]));
			radix2 #(.width(width)) rd_st5_411  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[411]), .rdlo_in(a5_wr[443]),  .coef_in(coef[864]), .rdup_out(a6_wr[411]), .rdlo_out(a6_wr[443]));
			radix2 #(.width(width)) rd_st5_412  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[412]), .rdlo_in(a5_wr[444]),  .coef_in(coef[896]), .rdup_out(a6_wr[412]), .rdlo_out(a6_wr[444]));
			radix2 #(.width(width)) rd_st5_413  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[413]), .rdlo_in(a5_wr[445]),  .coef_in(coef[928]), .rdup_out(a6_wr[413]), .rdlo_out(a6_wr[445]));
			radix2 #(.width(width)) rd_st5_414  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[414]), .rdlo_in(a5_wr[446]),  .coef_in(coef[960]), .rdup_out(a6_wr[414]), .rdlo_out(a6_wr[446]));
			radix2 #(.width(width)) rd_st5_415  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[415]), .rdlo_in(a5_wr[447]),  .coef_in(coef[992]), .rdup_out(a6_wr[415]), .rdlo_out(a6_wr[447]));
			radix2 #(.width(width)) rd_st5_448  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[448]), .rdlo_in(a5_wr[480]),  .coef_in(coef[0]), .rdup_out(a6_wr[448]), .rdlo_out(a6_wr[480]));
			radix2 #(.width(width)) rd_st5_449  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[449]), .rdlo_in(a5_wr[481]),  .coef_in(coef[32]), .rdup_out(a6_wr[449]), .rdlo_out(a6_wr[481]));
			radix2 #(.width(width)) rd_st5_450  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[450]), .rdlo_in(a5_wr[482]),  .coef_in(coef[64]), .rdup_out(a6_wr[450]), .rdlo_out(a6_wr[482]));
			radix2 #(.width(width)) rd_st5_451  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[451]), .rdlo_in(a5_wr[483]),  .coef_in(coef[96]), .rdup_out(a6_wr[451]), .rdlo_out(a6_wr[483]));
			radix2 #(.width(width)) rd_st5_452  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[452]), .rdlo_in(a5_wr[484]),  .coef_in(coef[128]), .rdup_out(a6_wr[452]), .rdlo_out(a6_wr[484]));
			radix2 #(.width(width)) rd_st5_453  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[453]), .rdlo_in(a5_wr[485]),  .coef_in(coef[160]), .rdup_out(a6_wr[453]), .rdlo_out(a6_wr[485]));
			radix2 #(.width(width)) rd_st5_454  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[454]), .rdlo_in(a5_wr[486]),  .coef_in(coef[192]), .rdup_out(a6_wr[454]), .rdlo_out(a6_wr[486]));
			radix2 #(.width(width)) rd_st5_455  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[455]), .rdlo_in(a5_wr[487]),  .coef_in(coef[224]), .rdup_out(a6_wr[455]), .rdlo_out(a6_wr[487]));
			radix2 #(.width(width)) rd_st5_456  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[456]), .rdlo_in(a5_wr[488]),  .coef_in(coef[256]), .rdup_out(a6_wr[456]), .rdlo_out(a6_wr[488]));
			radix2 #(.width(width)) rd_st5_457  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[457]), .rdlo_in(a5_wr[489]),  .coef_in(coef[288]), .rdup_out(a6_wr[457]), .rdlo_out(a6_wr[489]));
			radix2 #(.width(width)) rd_st5_458  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[458]), .rdlo_in(a5_wr[490]),  .coef_in(coef[320]), .rdup_out(a6_wr[458]), .rdlo_out(a6_wr[490]));
			radix2 #(.width(width)) rd_st5_459  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[459]), .rdlo_in(a5_wr[491]),  .coef_in(coef[352]), .rdup_out(a6_wr[459]), .rdlo_out(a6_wr[491]));
			radix2 #(.width(width)) rd_st5_460  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[460]), .rdlo_in(a5_wr[492]),  .coef_in(coef[384]), .rdup_out(a6_wr[460]), .rdlo_out(a6_wr[492]));
			radix2 #(.width(width)) rd_st5_461  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[461]), .rdlo_in(a5_wr[493]),  .coef_in(coef[416]), .rdup_out(a6_wr[461]), .rdlo_out(a6_wr[493]));
			radix2 #(.width(width)) rd_st5_462  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[462]), .rdlo_in(a5_wr[494]),  .coef_in(coef[448]), .rdup_out(a6_wr[462]), .rdlo_out(a6_wr[494]));
			radix2 #(.width(width)) rd_st5_463  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[463]), .rdlo_in(a5_wr[495]),  .coef_in(coef[480]), .rdup_out(a6_wr[463]), .rdlo_out(a6_wr[495]));
			radix2 #(.width(width)) rd_st5_464  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[464]), .rdlo_in(a5_wr[496]),  .coef_in(coef[512]), .rdup_out(a6_wr[464]), .rdlo_out(a6_wr[496]));
			radix2 #(.width(width)) rd_st5_465  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[465]), .rdlo_in(a5_wr[497]),  .coef_in(coef[544]), .rdup_out(a6_wr[465]), .rdlo_out(a6_wr[497]));
			radix2 #(.width(width)) rd_st5_466  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[466]), .rdlo_in(a5_wr[498]),  .coef_in(coef[576]), .rdup_out(a6_wr[466]), .rdlo_out(a6_wr[498]));
			radix2 #(.width(width)) rd_st5_467  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[467]), .rdlo_in(a5_wr[499]),  .coef_in(coef[608]), .rdup_out(a6_wr[467]), .rdlo_out(a6_wr[499]));
			radix2 #(.width(width)) rd_st5_468  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[468]), .rdlo_in(a5_wr[500]),  .coef_in(coef[640]), .rdup_out(a6_wr[468]), .rdlo_out(a6_wr[500]));
			radix2 #(.width(width)) rd_st5_469  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[469]), .rdlo_in(a5_wr[501]),  .coef_in(coef[672]), .rdup_out(a6_wr[469]), .rdlo_out(a6_wr[501]));
			radix2 #(.width(width)) rd_st5_470  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[470]), .rdlo_in(a5_wr[502]),  .coef_in(coef[704]), .rdup_out(a6_wr[470]), .rdlo_out(a6_wr[502]));
			radix2 #(.width(width)) rd_st5_471  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[471]), .rdlo_in(a5_wr[503]),  .coef_in(coef[736]), .rdup_out(a6_wr[471]), .rdlo_out(a6_wr[503]));
			radix2 #(.width(width)) rd_st5_472  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[472]), .rdlo_in(a5_wr[504]),  .coef_in(coef[768]), .rdup_out(a6_wr[472]), .rdlo_out(a6_wr[504]));
			radix2 #(.width(width)) rd_st5_473  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[473]), .rdlo_in(a5_wr[505]),  .coef_in(coef[800]), .rdup_out(a6_wr[473]), .rdlo_out(a6_wr[505]));
			radix2 #(.width(width)) rd_st5_474  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[474]), .rdlo_in(a5_wr[506]),  .coef_in(coef[832]), .rdup_out(a6_wr[474]), .rdlo_out(a6_wr[506]));
			radix2 #(.width(width)) rd_st5_475  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[475]), .rdlo_in(a5_wr[507]),  .coef_in(coef[864]), .rdup_out(a6_wr[475]), .rdlo_out(a6_wr[507]));
			radix2 #(.width(width)) rd_st5_476  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[476]), .rdlo_in(a5_wr[508]),  .coef_in(coef[896]), .rdup_out(a6_wr[476]), .rdlo_out(a6_wr[508]));
			radix2 #(.width(width)) rd_st5_477  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[477]), .rdlo_in(a5_wr[509]),  .coef_in(coef[928]), .rdup_out(a6_wr[477]), .rdlo_out(a6_wr[509]));
			radix2 #(.width(width)) rd_st5_478  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[478]), .rdlo_in(a5_wr[510]),  .coef_in(coef[960]), .rdup_out(a6_wr[478]), .rdlo_out(a6_wr[510]));
			radix2 #(.width(width)) rd_st5_479  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[479]), .rdlo_in(a5_wr[511]),  .coef_in(coef[992]), .rdup_out(a6_wr[479]), .rdlo_out(a6_wr[511]));
			radix2 #(.width(width)) rd_st5_512  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[512]), .rdlo_in(a5_wr[544]),  .coef_in(coef[0]), .rdup_out(a6_wr[512]), .rdlo_out(a6_wr[544]));
			radix2 #(.width(width)) rd_st5_513  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[513]), .rdlo_in(a5_wr[545]),  .coef_in(coef[32]), .rdup_out(a6_wr[513]), .rdlo_out(a6_wr[545]));
			radix2 #(.width(width)) rd_st5_514  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[514]), .rdlo_in(a5_wr[546]),  .coef_in(coef[64]), .rdup_out(a6_wr[514]), .rdlo_out(a6_wr[546]));
			radix2 #(.width(width)) rd_st5_515  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[515]), .rdlo_in(a5_wr[547]),  .coef_in(coef[96]), .rdup_out(a6_wr[515]), .rdlo_out(a6_wr[547]));
			radix2 #(.width(width)) rd_st5_516  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[516]), .rdlo_in(a5_wr[548]),  .coef_in(coef[128]), .rdup_out(a6_wr[516]), .rdlo_out(a6_wr[548]));
			radix2 #(.width(width)) rd_st5_517  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[517]), .rdlo_in(a5_wr[549]),  .coef_in(coef[160]), .rdup_out(a6_wr[517]), .rdlo_out(a6_wr[549]));
			radix2 #(.width(width)) rd_st5_518  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[518]), .rdlo_in(a5_wr[550]),  .coef_in(coef[192]), .rdup_out(a6_wr[518]), .rdlo_out(a6_wr[550]));
			radix2 #(.width(width)) rd_st5_519  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[519]), .rdlo_in(a5_wr[551]),  .coef_in(coef[224]), .rdup_out(a6_wr[519]), .rdlo_out(a6_wr[551]));
			radix2 #(.width(width)) rd_st5_520  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[520]), .rdlo_in(a5_wr[552]),  .coef_in(coef[256]), .rdup_out(a6_wr[520]), .rdlo_out(a6_wr[552]));
			radix2 #(.width(width)) rd_st5_521  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[521]), .rdlo_in(a5_wr[553]),  .coef_in(coef[288]), .rdup_out(a6_wr[521]), .rdlo_out(a6_wr[553]));
			radix2 #(.width(width)) rd_st5_522  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[522]), .rdlo_in(a5_wr[554]),  .coef_in(coef[320]), .rdup_out(a6_wr[522]), .rdlo_out(a6_wr[554]));
			radix2 #(.width(width)) rd_st5_523  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[523]), .rdlo_in(a5_wr[555]),  .coef_in(coef[352]), .rdup_out(a6_wr[523]), .rdlo_out(a6_wr[555]));
			radix2 #(.width(width)) rd_st5_524  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[524]), .rdlo_in(a5_wr[556]),  .coef_in(coef[384]), .rdup_out(a6_wr[524]), .rdlo_out(a6_wr[556]));
			radix2 #(.width(width)) rd_st5_525  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[525]), .rdlo_in(a5_wr[557]),  .coef_in(coef[416]), .rdup_out(a6_wr[525]), .rdlo_out(a6_wr[557]));
			radix2 #(.width(width)) rd_st5_526  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[526]), .rdlo_in(a5_wr[558]),  .coef_in(coef[448]), .rdup_out(a6_wr[526]), .rdlo_out(a6_wr[558]));
			radix2 #(.width(width)) rd_st5_527  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[527]), .rdlo_in(a5_wr[559]),  .coef_in(coef[480]), .rdup_out(a6_wr[527]), .rdlo_out(a6_wr[559]));
			radix2 #(.width(width)) rd_st5_528  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[528]), .rdlo_in(a5_wr[560]),  .coef_in(coef[512]), .rdup_out(a6_wr[528]), .rdlo_out(a6_wr[560]));
			radix2 #(.width(width)) rd_st5_529  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[529]), .rdlo_in(a5_wr[561]),  .coef_in(coef[544]), .rdup_out(a6_wr[529]), .rdlo_out(a6_wr[561]));
			radix2 #(.width(width)) rd_st5_530  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[530]), .rdlo_in(a5_wr[562]),  .coef_in(coef[576]), .rdup_out(a6_wr[530]), .rdlo_out(a6_wr[562]));
			radix2 #(.width(width)) rd_st5_531  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[531]), .rdlo_in(a5_wr[563]),  .coef_in(coef[608]), .rdup_out(a6_wr[531]), .rdlo_out(a6_wr[563]));
			radix2 #(.width(width)) rd_st5_532  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[532]), .rdlo_in(a5_wr[564]),  .coef_in(coef[640]), .rdup_out(a6_wr[532]), .rdlo_out(a6_wr[564]));
			radix2 #(.width(width)) rd_st5_533  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[533]), .rdlo_in(a5_wr[565]),  .coef_in(coef[672]), .rdup_out(a6_wr[533]), .rdlo_out(a6_wr[565]));
			radix2 #(.width(width)) rd_st5_534  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[534]), .rdlo_in(a5_wr[566]),  .coef_in(coef[704]), .rdup_out(a6_wr[534]), .rdlo_out(a6_wr[566]));
			radix2 #(.width(width)) rd_st5_535  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[535]), .rdlo_in(a5_wr[567]),  .coef_in(coef[736]), .rdup_out(a6_wr[535]), .rdlo_out(a6_wr[567]));
			radix2 #(.width(width)) rd_st5_536  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[536]), .rdlo_in(a5_wr[568]),  .coef_in(coef[768]), .rdup_out(a6_wr[536]), .rdlo_out(a6_wr[568]));
			radix2 #(.width(width)) rd_st5_537  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[537]), .rdlo_in(a5_wr[569]),  .coef_in(coef[800]), .rdup_out(a6_wr[537]), .rdlo_out(a6_wr[569]));
			radix2 #(.width(width)) rd_st5_538  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[538]), .rdlo_in(a5_wr[570]),  .coef_in(coef[832]), .rdup_out(a6_wr[538]), .rdlo_out(a6_wr[570]));
			radix2 #(.width(width)) rd_st5_539  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[539]), .rdlo_in(a5_wr[571]),  .coef_in(coef[864]), .rdup_out(a6_wr[539]), .rdlo_out(a6_wr[571]));
			radix2 #(.width(width)) rd_st5_540  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[540]), .rdlo_in(a5_wr[572]),  .coef_in(coef[896]), .rdup_out(a6_wr[540]), .rdlo_out(a6_wr[572]));
			radix2 #(.width(width)) rd_st5_541  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[541]), .rdlo_in(a5_wr[573]),  .coef_in(coef[928]), .rdup_out(a6_wr[541]), .rdlo_out(a6_wr[573]));
			radix2 #(.width(width)) rd_st5_542  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[542]), .rdlo_in(a5_wr[574]),  .coef_in(coef[960]), .rdup_out(a6_wr[542]), .rdlo_out(a6_wr[574]));
			radix2 #(.width(width)) rd_st5_543  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[543]), .rdlo_in(a5_wr[575]),  .coef_in(coef[992]), .rdup_out(a6_wr[543]), .rdlo_out(a6_wr[575]));
			radix2 #(.width(width)) rd_st5_576  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[576]), .rdlo_in(a5_wr[608]),  .coef_in(coef[0]), .rdup_out(a6_wr[576]), .rdlo_out(a6_wr[608]));
			radix2 #(.width(width)) rd_st5_577  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[577]), .rdlo_in(a5_wr[609]),  .coef_in(coef[32]), .rdup_out(a6_wr[577]), .rdlo_out(a6_wr[609]));
			radix2 #(.width(width)) rd_st5_578  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[578]), .rdlo_in(a5_wr[610]),  .coef_in(coef[64]), .rdup_out(a6_wr[578]), .rdlo_out(a6_wr[610]));
			radix2 #(.width(width)) rd_st5_579  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[579]), .rdlo_in(a5_wr[611]),  .coef_in(coef[96]), .rdup_out(a6_wr[579]), .rdlo_out(a6_wr[611]));
			radix2 #(.width(width)) rd_st5_580  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[580]), .rdlo_in(a5_wr[612]),  .coef_in(coef[128]), .rdup_out(a6_wr[580]), .rdlo_out(a6_wr[612]));
			radix2 #(.width(width)) rd_st5_581  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[581]), .rdlo_in(a5_wr[613]),  .coef_in(coef[160]), .rdup_out(a6_wr[581]), .rdlo_out(a6_wr[613]));
			radix2 #(.width(width)) rd_st5_582  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[582]), .rdlo_in(a5_wr[614]),  .coef_in(coef[192]), .rdup_out(a6_wr[582]), .rdlo_out(a6_wr[614]));
			radix2 #(.width(width)) rd_st5_583  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[583]), .rdlo_in(a5_wr[615]),  .coef_in(coef[224]), .rdup_out(a6_wr[583]), .rdlo_out(a6_wr[615]));
			radix2 #(.width(width)) rd_st5_584  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[584]), .rdlo_in(a5_wr[616]),  .coef_in(coef[256]), .rdup_out(a6_wr[584]), .rdlo_out(a6_wr[616]));
			radix2 #(.width(width)) rd_st5_585  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[585]), .rdlo_in(a5_wr[617]),  .coef_in(coef[288]), .rdup_out(a6_wr[585]), .rdlo_out(a6_wr[617]));
			radix2 #(.width(width)) rd_st5_586  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[586]), .rdlo_in(a5_wr[618]),  .coef_in(coef[320]), .rdup_out(a6_wr[586]), .rdlo_out(a6_wr[618]));
			radix2 #(.width(width)) rd_st5_587  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[587]), .rdlo_in(a5_wr[619]),  .coef_in(coef[352]), .rdup_out(a6_wr[587]), .rdlo_out(a6_wr[619]));
			radix2 #(.width(width)) rd_st5_588  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[588]), .rdlo_in(a5_wr[620]),  .coef_in(coef[384]), .rdup_out(a6_wr[588]), .rdlo_out(a6_wr[620]));
			radix2 #(.width(width)) rd_st5_589  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[589]), .rdlo_in(a5_wr[621]),  .coef_in(coef[416]), .rdup_out(a6_wr[589]), .rdlo_out(a6_wr[621]));
			radix2 #(.width(width)) rd_st5_590  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[590]), .rdlo_in(a5_wr[622]),  .coef_in(coef[448]), .rdup_out(a6_wr[590]), .rdlo_out(a6_wr[622]));
			radix2 #(.width(width)) rd_st5_591  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[591]), .rdlo_in(a5_wr[623]),  .coef_in(coef[480]), .rdup_out(a6_wr[591]), .rdlo_out(a6_wr[623]));
			radix2 #(.width(width)) rd_st5_592  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[592]), .rdlo_in(a5_wr[624]),  .coef_in(coef[512]), .rdup_out(a6_wr[592]), .rdlo_out(a6_wr[624]));
			radix2 #(.width(width)) rd_st5_593  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[593]), .rdlo_in(a5_wr[625]),  .coef_in(coef[544]), .rdup_out(a6_wr[593]), .rdlo_out(a6_wr[625]));
			radix2 #(.width(width)) rd_st5_594  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[594]), .rdlo_in(a5_wr[626]),  .coef_in(coef[576]), .rdup_out(a6_wr[594]), .rdlo_out(a6_wr[626]));
			radix2 #(.width(width)) rd_st5_595  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[595]), .rdlo_in(a5_wr[627]),  .coef_in(coef[608]), .rdup_out(a6_wr[595]), .rdlo_out(a6_wr[627]));
			radix2 #(.width(width)) rd_st5_596  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[596]), .rdlo_in(a5_wr[628]),  .coef_in(coef[640]), .rdup_out(a6_wr[596]), .rdlo_out(a6_wr[628]));
			radix2 #(.width(width)) rd_st5_597  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[597]), .rdlo_in(a5_wr[629]),  .coef_in(coef[672]), .rdup_out(a6_wr[597]), .rdlo_out(a6_wr[629]));
			radix2 #(.width(width)) rd_st5_598  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[598]), .rdlo_in(a5_wr[630]),  .coef_in(coef[704]), .rdup_out(a6_wr[598]), .rdlo_out(a6_wr[630]));
			radix2 #(.width(width)) rd_st5_599  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[599]), .rdlo_in(a5_wr[631]),  .coef_in(coef[736]), .rdup_out(a6_wr[599]), .rdlo_out(a6_wr[631]));
			radix2 #(.width(width)) rd_st5_600  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[600]), .rdlo_in(a5_wr[632]),  .coef_in(coef[768]), .rdup_out(a6_wr[600]), .rdlo_out(a6_wr[632]));
			radix2 #(.width(width)) rd_st5_601  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[601]), .rdlo_in(a5_wr[633]),  .coef_in(coef[800]), .rdup_out(a6_wr[601]), .rdlo_out(a6_wr[633]));
			radix2 #(.width(width)) rd_st5_602  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[602]), .rdlo_in(a5_wr[634]),  .coef_in(coef[832]), .rdup_out(a6_wr[602]), .rdlo_out(a6_wr[634]));
			radix2 #(.width(width)) rd_st5_603  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[603]), .rdlo_in(a5_wr[635]),  .coef_in(coef[864]), .rdup_out(a6_wr[603]), .rdlo_out(a6_wr[635]));
			radix2 #(.width(width)) rd_st5_604  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[604]), .rdlo_in(a5_wr[636]),  .coef_in(coef[896]), .rdup_out(a6_wr[604]), .rdlo_out(a6_wr[636]));
			radix2 #(.width(width)) rd_st5_605  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[605]), .rdlo_in(a5_wr[637]),  .coef_in(coef[928]), .rdup_out(a6_wr[605]), .rdlo_out(a6_wr[637]));
			radix2 #(.width(width)) rd_st5_606  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[606]), .rdlo_in(a5_wr[638]),  .coef_in(coef[960]), .rdup_out(a6_wr[606]), .rdlo_out(a6_wr[638]));
			radix2 #(.width(width)) rd_st5_607  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[607]), .rdlo_in(a5_wr[639]),  .coef_in(coef[992]), .rdup_out(a6_wr[607]), .rdlo_out(a6_wr[639]));
			radix2 #(.width(width)) rd_st5_640  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[640]), .rdlo_in(a5_wr[672]),  .coef_in(coef[0]), .rdup_out(a6_wr[640]), .rdlo_out(a6_wr[672]));
			radix2 #(.width(width)) rd_st5_641  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[641]), .rdlo_in(a5_wr[673]),  .coef_in(coef[32]), .rdup_out(a6_wr[641]), .rdlo_out(a6_wr[673]));
			radix2 #(.width(width)) rd_st5_642  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[642]), .rdlo_in(a5_wr[674]),  .coef_in(coef[64]), .rdup_out(a6_wr[642]), .rdlo_out(a6_wr[674]));
			radix2 #(.width(width)) rd_st5_643  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[643]), .rdlo_in(a5_wr[675]),  .coef_in(coef[96]), .rdup_out(a6_wr[643]), .rdlo_out(a6_wr[675]));
			radix2 #(.width(width)) rd_st5_644  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[644]), .rdlo_in(a5_wr[676]),  .coef_in(coef[128]), .rdup_out(a6_wr[644]), .rdlo_out(a6_wr[676]));
			radix2 #(.width(width)) rd_st5_645  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[645]), .rdlo_in(a5_wr[677]),  .coef_in(coef[160]), .rdup_out(a6_wr[645]), .rdlo_out(a6_wr[677]));
			radix2 #(.width(width)) rd_st5_646  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[646]), .rdlo_in(a5_wr[678]),  .coef_in(coef[192]), .rdup_out(a6_wr[646]), .rdlo_out(a6_wr[678]));
			radix2 #(.width(width)) rd_st5_647  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[647]), .rdlo_in(a5_wr[679]),  .coef_in(coef[224]), .rdup_out(a6_wr[647]), .rdlo_out(a6_wr[679]));
			radix2 #(.width(width)) rd_st5_648  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[648]), .rdlo_in(a5_wr[680]),  .coef_in(coef[256]), .rdup_out(a6_wr[648]), .rdlo_out(a6_wr[680]));
			radix2 #(.width(width)) rd_st5_649  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[649]), .rdlo_in(a5_wr[681]),  .coef_in(coef[288]), .rdup_out(a6_wr[649]), .rdlo_out(a6_wr[681]));
			radix2 #(.width(width)) rd_st5_650  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[650]), .rdlo_in(a5_wr[682]),  .coef_in(coef[320]), .rdup_out(a6_wr[650]), .rdlo_out(a6_wr[682]));
			radix2 #(.width(width)) rd_st5_651  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[651]), .rdlo_in(a5_wr[683]),  .coef_in(coef[352]), .rdup_out(a6_wr[651]), .rdlo_out(a6_wr[683]));
			radix2 #(.width(width)) rd_st5_652  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[652]), .rdlo_in(a5_wr[684]),  .coef_in(coef[384]), .rdup_out(a6_wr[652]), .rdlo_out(a6_wr[684]));
			radix2 #(.width(width)) rd_st5_653  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[653]), .rdlo_in(a5_wr[685]),  .coef_in(coef[416]), .rdup_out(a6_wr[653]), .rdlo_out(a6_wr[685]));
			radix2 #(.width(width)) rd_st5_654  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[654]), .rdlo_in(a5_wr[686]),  .coef_in(coef[448]), .rdup_out(a6_wr[654]), .rdlo_out(a6_wr[686]));
			radix2 #(.width(width)) rd_st5_655  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[655]), .rdlo_in(a5_wr[687]),  .coef_in(coef[480]), .rdup_out(a6_wr[655]), .rdlo_out(a6_wr[687]));
			radix2 #(.width(width)) rd_st5_656  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[656]), .rdlo_in(a5_wr[688]),  .coef_in(coef[512]), .rdup_out(a6_wr[656]), .rdlo_out(a6_wr[688]));
			radix2 #(.width(width)) rd_st5_657  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[657]), .rdlo_in(a5_wr[689]),  .coef_in(coef[544]), .rdup_out(a6_wr[657]), .rdlo_out(a6_wr[689]));
			radix2 #(.width(width)) rd_st5_658  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[658]), .rdlo_in(a5_wr[690]),  .coef_in(coef[576]), .rdup_out(a6_wr[658]), .rdlo_out(a6_wr[690]));
			radix2 #(.width(width)) rd_st5_659  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[659]), .rdlo_in(a5_wr[691]),  .coef_in(coef[608]), .rdup_out(a6_wr[659]), .rdlo_out(a6_wr[691]));
			radix2 #(.width(width)) rd_st5_660  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[660]), .rdlo_in(a5_wr[692]),  .coef_in(coef[640]), .rdup_out(a6_wr[660]), .rdlo_out(a6_wr[692]));
			radix2 #(.width(width)) rd_st5_661  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[661]), .rdlo_in(a5_wr[693]),  .coef_in(coef[672]), .rdup_out(a6_wr[661]), .rdlo_out(a6_wr[693]));
			radix2 #(.width(width)) rd_st5_662  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[662]), .rdlo_in(a5_wr[694]),  .coef_in(coef[704]), .rdup_out(a6_wr[662]), .rdlo_out(a6_wr[694]));
			radix2 #(.width(width)) rd_st5_663  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[663]), .rdlo_in(a5_wr[695]),  .coef_in(coef[736]), .rdup_out(a6_wr[663]), .rdlo_out(a6_wr[695]));
			radix2 #(.width(width)) rd_st5_664  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[664]), .rdlo_in(a5_wr[696]),  .coef_in(coef[768]), .rdup_out(a6_wr[664]), .rdlo_out(a6_wr[696]));
			radix2 #(.width(width)) rd_st5_665  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[665]), .rdlo_in(a5_wr[697]),  .coef_in(coef[800]), .rdup_out(a6_wr[665]), .rdlo_out(a6_wr[697]));
			radix2 #(.width(width)) rd_st5_666  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[666]), .rdlo_in(a5_wr[698]),  .coef_in(coef[832]), .rdup_out(a6_wr[666]), .rdlo_out(a6_wr[698]));
			radix2 #(.width(width)) rd_st5_667  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[667]), .rdlo_in(a5_wr[699]),  .coef_in(coef[864]), .rdup_out(a6_wr[667]), .rdlo_out(a6_wr[699]));
			radix2 #(.width(width)) rd_st5_668  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[668]), .rdlo_in(a5_wr[700]),  .coef_in(coef[896]), .rdup_out(a6_wr[668]), .rdlo_out(a6_wr[700]));
			radix2 #(.width(width)) rd_st5_669  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[669]), .rdlo_in(a5_wr[701]),  .coef_in(coef[928]), .rdup_out(a6_wr[669]), .rdlo_out(a6_wr[701]));
			radix2 #(.width(width)) rd_st5_670  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[670]), .rdlo_in(a5_wr[702]),  .coef_in(coef[960]), .rdup_out(a6_wr[670]), .rdlo_out(a6_wr[702]));
			radix2 #(.width(width)) rd_st5_671  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[671]), .rdlo_in(a5_wr[703]),  .coef_in(coef[992]), .rdup_out(a6_wr[671]), .rdlo_out(a6_wr[703]));
			radix2 #(.width(width)) rd_st5_704  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[704]), .rdlo_in(a5_wr[736]),  .coef_in(coef[0]), .rdup_out(a6_wr[704]), .rdlo_out(a6_wr[736]));
			radix2 #(.width(width)) rd_st5_705  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[705]), .rdlo_in(a5_wr[737]),  .coef_in(coef[32]), .rdup_out(a6_wr[705]), .rdlo_out(a6_wr[737]));
			radix2 #(.width(width)) rd_st5_706  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[706]), .rdlo_in(a5_wr[738]),  .coef_in(coef[64]), .rdup_out(a6_wr[706]), .rdlo_out(a6_wr[738]));
			radix2 #(.width(width)) rd_st5_707  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[707]), .rdlo_in(a5_wr[739]),  .coef_in(coef[96]), .rdup_out(a6_wr[707]), .rdlo_out(a6_wr[739]));
			radix2 #(.width(width)) rd_st5_708  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[708]), .rdlo_in(a5_wr[740]),  .coef_in(coef[128]), .rdup_out(a6_wr[708]), .rdlo_out(a6_wr[740]));
			radix2 #(.width(width)) rd_st5_709  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[709]), .rdlo_in(a5_wr[741]),  .coef_in(coef[160]), .rdup_out(a6_wr[709]), .rdlo_out(a6_wr[741]));
			radix2 #(.width(width)) rd_st5_710  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[710]), .rdlo_in(a5_wr[742]),  .coef_in(coef[192]), .rdup_out(a6_wr[710]), .rdlo_out(a6_wr[742]));
			radix2 #(.width(width)) rd_st5_711  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[711]), .rdlo_in(a5_wr[743]),  .coef_in(coef[224]), .rdup_out(a6_wr[711]), .rdlo_out(a6_wr[743]));
			radix2 #(.width(width)) rd_st5_712  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[712]), .rdlo_in(a5_wr[744]),  .coef_in(coef[256]), .rdup_out(a6_wr[712]), .rdlo_out(a6_wr[744]));
			radix2 #(.width(width)) rd_st5_713  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[713]), .rdlo_in(a5_wr[745]),  .coef_in(coef[288]), .rdup_out(a6_wr[713]), .rdlo_out(a6_wr[745]));
			radix2 #(.width(width)) rd_st5_714  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[714]), .rdlo_in(a5_wr[746]),  .coef_in(coef[320]), .rdup_out(a6_wr[714]), .rdlo_out(a6_wr[746]));
			radix2 #(.width(width)) rd_st5_715  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[715]), .rdlo_in(a5_wr[747]),  .coef_in(coef[352]), .rdup_out(a6_wr[715]), .rdlo_out(a6_wr[747]));
			radix2 #(.width(width)) rd_st5_716  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[716]), .rdlo_in(a5_wr[748]),  .coef_in(coef[384]), .rdup_out(a6_wr[716]), .rdlo_out(a6_wr[748]));
			radix2 #(.width(width)) rd_st5_717  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[717]), .rdlo_in(a5_wr[749]),  .coef_in(coef[416]), .rdup_out(a6_wr[717]), .rdlo_out(a6_wr[749]));
			radix2 #(.width(width)) rd_st5_718  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[718]), .rdlo_in(a5_wr[750]),  .coef_in(coef[448]), .rdup_out(a6_wr[718]), .rdlo_out(a6_wr[750]));
			radix2 #(.width(width)) rd_st5_719  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[719]), .rdlo_in(a5_wr[751]),  .coef_in(coef[480]), .rdup_out(a6_wr[719]), .rdlo_out(a6_wr[751]));
			radix2 #(.width(width)) rd_st5_720  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[720]), .rdlo_in(a5_wr[752]),  .coef_in(coef[512]), .rdup_out(a6_wr[720]), .rdlo_out(a6_wr[752]));
			radix2 #(.width(width)) rd_st5_721  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[721]), .rdlo_in(a5_wr[753]),  .coef_in(coef[544]), .rdup_out(a6_wr[721]), .rdlo_out(a6_wr[753]));
			radix2 #(.width(width)) rd_st5_722  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[722]), .rdlo_in(a5_wr[754]),  .coef_in(coef[576]), .rdup_out(a6_wr[722]), .rdlo_out(a6_wr[754]));
			radix2 #(.width(width)) rd_st5_723  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[723]), .rdlo_in(a5_wr[755]),  .coef_in(coef[608]), .rdup_out(a6_wr[723]), .rdlo_out(a6_wr[755]));
			radix2 #(.width(width)) rd_st5_724  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[724]), .rdlo_in(a5_wr[756]),  .coef_in(coef[640]), .rdup_out(a6_wr[724]), .rdlo_out(a6_wr[756]));
			radix2 #(.width(width)) rd_st5_725  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[725]), .rdlo_in(a5_wr[757]),  .coef_in(coef[672]), .rdup_out(a6_wr[725]), .rdlo_out(a6_wr[757]));
			radix2 #(.width(width)) rd_st5_726  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[726]), .rdlo_in(a5_wr[758]),  .coef_in(coef[704]), .rdup_out(a6_wr[726]), .rdlo_out(a6_wr[758]));
			radix2 #(.width(width)) rd_st5_727  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[727]), .rdlo_in(a5_wr[759]),  .coef_in(coef[736]), .rdup_out(a6_wr[727]), .rdlo_out(a6_wr[759]));
			radix2 #(.width(width)) rd_st5_728  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[728]), .rdlo_in(a5_wr[760]),  .coef_in(coef[768]), .rdup_out(a6_wr[728]), .rdlo_out(a6_wr[760]));
			radix2 #(.width(width)) rd_st5_729  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[729]), .rdlo_in(a5_wr[761]),  .coef_in(coef[800]), .rdup_out(a6_wr[729]), .rdlo_out(a6_wr[761]));
			radix2 #(.width(width)) rd_st5_730  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[730]), .rdlo_in(a5_wr[762]),  .coef_in(coef[832]), .rdup_out(a6_wr[730]), .rdlo_out(a6_wr[762]));
			radix2 #(.width(width)) rd_st5_731  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[731]), .rdlo_in(a5_wr[763]),  .coef_in(coef[864]), .rdup_out(a6_wr[731]), .rdlo_out(a6_wr[763]));
			radix2 #(.width(width)) rd_st5_732  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[732]), .rdlo_in(a5_wr[764]),  .coef_in(coef[896]), .rdup_out(a6_wr[732]), .rdlo_out(a6_wr[764]));
			radix2 #(.width(width)) rd_st5_733  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[733]), .rdlo_in(a5_wr[765]),  .coef_in(coef[928]), .rdup_out(a6_wr[733]), .rdlo_out(a6_wr[765]));
			radix2 #(.width(width)) rd_st5_734  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[734]), .rdlo_in(a5_wr[766]),  .coef_in(coef[960]), .rdup_out(a6_wr[734]), .rdlo_out(a6_wr[766]));
			radix2 #(.width(width)) rd_st5_735  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[735]), .rdlo_in(a5_wr[767]),  .coef_in(coef[992]), .rdup_out(a6_wr[735]), .rdlo_out(a6_wr[767]));
			radix2 #(.width(width)) rd_st5_768  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[768]), .rdlo_in(a5_wr[800]),  .coef_in(coef[0]), .rdup_out(a6_wr[768]), .rdlo_out(a6_wr[800]));
			radix2 #(.width(width)) rd_st5_769  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[769]), .rdlo_in(a5_wr[801]),  .coef_in(coef[32]), .rdup_out(a6_wr[769]), .rdlo_out(a6_wr[801]));
			radix2 #(.width(width)) rd_st5_770  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[770]), .rdlo_in(a5_wr[802]),  .coef_in(coef[64]), .rdup_out(a6_wr[770]), .rdlo_out(a6_wr[802]));
			radix2 #(.width(width)) rd_st5_771  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[771]), .rdlo_in(a5_wr[803]),  .coef_in(coef[96]), .rdup_out(a6_wr[771]), .rdlo_out(a6_wr[803]));
			radix2 #(.width(width)) rd_st5_772  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[772]), .rdlo_in(a5_wr[804]),  .coef_in(coef[128]), .rdup_out(a6_wr[772]), .rdlo_out(a6_wr[804]));
			radix2 #(.width(width)) rd_st5_773  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[773]), .rdlo_in(a5_wr[805]),  .coef_in(coef[160]), .rdup_out(a6_wr[773]), .rdlo_out(a6_wr[805]));
			radix2 #(.width(width)) rd_st5_774  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[774]), .rdlo_in(a5_wr[806]),  .coef_in(coef[192]), .rdup_out(a6_wr[774]), .rdlo_out(a6_wr[806]));
			radix2 #(.width(width)) rd_st5_775  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[775]), .rdlo_in(a5_wr[807]),  .coef_in(coef[224]), .rdup_out(a6_wr[775]), .rdlo_out(a6_wr[807]));
			radix2 #(.width(width)) rd_st5_776  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[776]), .rdlo_in(a5_wr[808]),  .coef_in(coef[256]), .rdup_out(a6_wr[776]), .rdlo_out(a6_wr[808]));
			radix2 #(.width(width)) rd_st5_777  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[777]), .rdlo_in(a5_wr[809]),  .coef_in(coef[288]), .rdup_out(a6_wr[777]), .rdlo_out(a6_wr[809]));
			radix2 #(.width(width)) rd_st5_778  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[778]), .rdlo_in(a5_wr[810]),  .coef_in(coef[320]), .rdup_out(a6_wr[778]), .rdlo_out(a6_wr[810]));
			radix2 #(.width(width)) rd_st5_779  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[779]), .rdlo_in(a5_wr[811]),  .coef_in(coef[352]), .rdup_out(a6_wr[779]), .rdlo_out(a6_wr[811]));
			radix2 #(.width(width)) rd_st5_780  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[780]), .rdlo_in(a5_wr[812]),  .coef_in(coef[384]), .rdup_out(a6_wr[780]), .rdlo_out(a6_wr[812]));
			radix2 #(.width(width)) rd_st5_781  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[781]), .rdlo_in(a5_wr[813]),  .coef_in(coef[416]), .rdup_out(a6_wr[781]), .rdlo_out(a6_wr[813]));
			radix2 #(.width(width)) rd_st5_782  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[782]), .rdlo_in(a5_wr[814]),  .coef_in(coef[448]), .rdup_out(a6_wr[782]), .rdlo_out(a6_wr[814]));
			radix2 #(.width(width)) rd_st5_783  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[783]), .rdlo_in(a5_wr[815]),  .coef_in(coef[480]), .rdup_out(a6_wr[783]), .rdlo_out(a6_wr[815]));
			radix2 #(.width(width)) rd_st5_784  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[784]), .rdlo_in(a5_wr[816]),  .coef_in(coef[512]), .rdup_out(a6_wr[784]), .rdlo_out(a6_wr[816]));
			radix2 #(.width(width)) rd_st5_785  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[785]), .rdlo_in(a5_wr[817]),  .coef_in(coef[544]), .rdup_out(a6_wr[785]), .rdlo_out(a6_wr[817]));
			radix2 #(.width(width)) rd_st5_786  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[786]), .rdlo_in(a5_wr[818]),  .coef_in(coef[576]), .rdup_out(a6_wr[786]), .rdlo_out(a6_wr[818]));
			radix2 #(.width(width)) rd_st5_787  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[787]), .rdlo_in(a5_wr[819]),  .coef_in(coef[608]), .rdup_out(a6_wr[787]), .rdlo_out(a6_wr[819]));
			radix2 #(.width(width)) rd_st5_788  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[788]), .rdlo_in(a5_wr[820]),  .coef_in(coef[640]), .rdup_out(a6_wr[788]), .rdlo_out(a6_wr[820]));
			radix2 #(.width(width)) rd_st5_789  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[789]), .rdlo_in(a5_wr[821]),  .coef_in(coef[672]), .rdup_out(a6_wr[789]), .rdlo_out(a6_wr[821]));
			radix2 #(.width(width)) rd_st5_790  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[790]), .rdlo_in(a5_wr[822]),  .coef_in(coef[704]), .rdup_out(a6_wr[790]), .rdlo_out(a6_wr[822]));
			radix2 #(.width(width)) rd_st5_791  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[791]), .rdlo_in(a5_wr[823]),  .coef_in(coef[736]), .rdup_out(a6_wr[791]), .rdlo_out(a6_wr[823]));
			radix2 #(.width(width)) rd_st5_792  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[792]), .rdlo_in(a5_wr[824]),  .coef_in(coef[768]), .rdup_out(a6_wr[792]), .rdlo_out(a6_wr[824]));
			radix2 #(.width(width)) rd_st5_793  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[793]), .rdlo_in(a5_wr[825]),  .coef_in(coef[800]), .rdup_out(a6_wr[793]), .rdlo_out(a6_wr[825]));
			radix2 #(.width(width)) rd_st5_794  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[794]), .rdlo_in(a5_wr[826]),  .coef_in(coef[832]), .rdup_out(a6_wr[794]), .rdlo_out(a6_wr[826]));
			radix2 #(.width(width)) rd_st5_795  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[795]), .rdlo_in(a5_wr[827]),  .coef_in(coef[864]), .rdup_out(a6_wr[795]), .rdlo_out(a6_wr[827]));
			radix2 #(.width(width)) rd_st5_796  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[796]), .rdlo_in(a5_wr[828]),  .coef_in(coef[896]), .rdup_out(a6_wr[796]), .rdlo_out(a6_wr[828]));
			radix2 #(.width(width)) rd_st5_797  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[797]), .rdlo_in(a5_wr[829]),  .coef_in(coef[928]), .rdup_out(a6_wr[797]), .rdlo_out(a6_wr[829]));
			radix2 #(.width(width)) rd_st5_798  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[798]), .rdlo_in(a5_wr[830]),  .coef_in(coef[960]), .rdup_out(a6_wr[798]), .rdlo_out(a6_wr[830]));
			radix2 #(.width(width)) rd_st5_799  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[799]), .rdlo_in(a5_wr[831]),  .coef_in(coef[992]), .rdup_out(a6_wr[799]), .rdlo_out(a6_wr[831]));
			radix2 #(.width(width)) rd_st5_832  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[832]), .rdlo_in(a5_wr[864]),  .coef_in(coef[0]), .rdup_out(a6_wr[832]), .rdlo_out(a6_wr[864]));
			radix2 #(.width(width)) rd_st5_833  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[833]), .rdlo_in(a5_wr[865]),  .coef_in(coef[32]), .rdup_out(a6_wr[833]), .rdlo_out(a6_wr[865]));
			radix2 #(.width(width)) rd_st5_834  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[834]), .rdlo_in(a5_wr[866]),  .coef_in(coef[64]), .rdup_out(a6_wr[834]), .rdlo_out(a6_wr[866]));
			radix2 #(.width(width)) rd_st5_835  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[835]), .rdlo_in(a5_wr[867]),  .coef_in(coef[96]), .rdup_out(a6_wr[835]), .rdlo_out(a6_wr[867]));
			radix2 #(.width(width)) rd_st5_836  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[836]), .rdlo_in(a5_wr[868]),  .coef_in(coef[128]), .rdup_out(a6_wr[836]), .rdlo_out(a6_wr[868]));
			radix2 #(.width(width)) rd_st5_837  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[837]), .rdlo_in(a5_wr[869]),  .coef_in(coef[160]), .rdup_out(a6_wr[837]), .rdlo_out(a6_wr[869]));
			radix2 #(.width(width)) rd_st5_838  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[838]), .rdlo_in(a5_wr[870]),  .coef_in(coef[192]), .rdup_out(a6_wr[838]), .rdlo_out(a6_wr[870]));
			radix2 #(.width(width)) rd_st5_839  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[839]), .rdlo_in(a5_wr[871]),  .coef_in(coef[224]), .rdup_out(a6_wr[839]), .rdlo_out(a6_wr[871]));
			radix2 #(.width(width)) rd_st5_840  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[840]), .rdlo_in(a5_wr[872]),  .coef_in(coef[256]), .rdup_out(a6_wr[840]), .rdlo_out(a6_wr[872]));
			radix2 #(.width(width)) rd_st5_841  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[841]), .rdlo_in(a5_wr[873]),  .coef_in(coef[288]), .rdup_out(a6_wr[841]), .rdlo_out(a6_wr[873]));
			radix2 #(.width(width)) rd_st5_842  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[842]), .rdlo_in(a5_wr[874]),  .coef_in(coef[320]), .rdup_out(a6_wr[842]), .rdlo_out(a6_wr[874]));
			radix2 #(.width(width)) rd_st5_843  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[843]), .rdlo_in(a5_wr[875]),  .coef_in(coef[352]), .rdup_out(a6_wr[843]), .rdlo_out(a6_wr[875]));
			radix2 #(.width(width)) rd_st5_844  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[844]), .rdlo_in(a5_wr[876]),  .coef_in(coef[384]), .rdup_out(a6_wr[844]), .rdlo_out(a6_wr[876]));
			radix2 #(.width(width)) rd_st5_845  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[845]), .rdlo_in(a5_wr[877]),  .coef_in(coef[416]), .rdup_out(a6_wr[845]), .rdlo_out(a6_wr[877]));
			radix2 #(.width(width)) rd_st5_846  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[846]), .rdlo_in(a5_wr[878]),  .coef_in(coef[448]), .rdup_out(a6_wr[846]), .rdlo_out(a6_wr[878]));
			radix2 #(.width(width)) rd_st5_847  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[847]), .rdlo_in(a5_wr[879]),  .coef_in(coef[480]), .rdup_out(a6_wr[847]), .rdlo_out(a6_wr[879]));
			radix2 #(.width(width)) rd_st5_848  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[848]), .rdlo_in(a5_wr[880]),  .coef_in(coef[512]), .rdup_out(a6_wr[848]), .rdlo_out(a6_wr[880]));
			radix2 #(.width(width)) rd_st5_849  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[849]), .rdlo_in(a5_wr[881]),  .coef_in(coef[544]), .rdup_out(a6_wr[849]), .rdlo_out(a6_wr[881]));
			radix2 #(.width(width)) rd_st5_850  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[850]), .rdlo_in(a5_wr[882]),  .coef_in(coef[576]), .rdup_out(a6_wr[850]), .rdlo_out(a6_wr[882]));
			radix2 #(.width(width)) rd_st5_851  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[851]), .rdlo_in(a5_wr[883]),  .coef_in(coef[608]), .rdup_out(a6_wr[851]), .rdlo_out(a6_wr[883]));
			radix2 #(.width(width)) rd_st5_852  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[852]), .rdlo_in(a5_wr[884]),  .coef_in(coef[640]), .rdup_out(a6_wr[852]), .rdlo_out(a6_wr[884]));
			radix2 #(.width(width)) rd_st5_853  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[853]), .rdlo_in(a5_wr[885]),  .coef_in(coef[672]), .rdup_out(a6_wr[853]), .rdlo_out(a6_wr[885]));
			radix2 #(.width(width)) rd_st5_854  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[854]), .rdlo_in(a5_wr[886]),  .coef_in(coef[704]), .rdup_out(a6_wr[854]), .rdlo_out(a6_wr[886]));
			radix2 #(.width(width)) rd_st5_855  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[855]), .rdlo_in(a5_wr[887]),  .coef_in(coef[736]), .rdup_out(a6_wr[855]), .rdlo_out(a6_wr[887]));
			radix2 #(.width(width)) rd_st5_856  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[856]), .rdlo_in(a5_wr[888]),  .coef_in(coef[768]), .rdup_out(a6_wr[856]), .rdlo_out(a6_wr[888]));
			radix2 #(.width(width)) rd_st5_857  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[857]), .rdlo_in(a5_wr[889]),  .coef_in(coef[800]), .rdup_out(a6_wr[857]), .rdlo_out(a6_wr[889]));
			radix2 #(.width(width)) rd_st5_858  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[858]), .rdlo_in(a5_wr[890]),  .coef_in(coef[832]), .rdup_out(a6_wr[858]), .rdlo_out(a6_wr[890]));
			radix2 #(.width(width)) rd_st5_859  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[859]), .rdlo_in(a5_wr[891]),  .coef_in(coef[864]), .rdup_out(a6_wr[859]), .rdlo_out(a6_wr[891]));
			radix2 #(.width(width)) rd_st5_860  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[860]), .rdlo_in(a5_wr[892]),  .coef_in(coef[896]), .rdup_out(a6_wr[860]), .rdlo_out(a6_wr[892]));
			radix2 #(.width(width)) rd_st5_861  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[861]), .rdlo_in(a5_wr[893]),  .coef_in(coef[928]), .rdup_out(a6_wr[861]), .rdlo_out(a6_wr[893]));
			radix2 #(.width(width)) rd_st5_862  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[862]), .rdlo_in(a5_wr[894]),  .coef_in(coef[960]), .rdup_out(a6_wr[862]), .rdlo_out(a6_wr[894]));
			radix2 #(.width(width)) rd_st5_863  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[863]), .rdlo_in(a5_wr[895]),  .coef_in(coef[992]), .rdup_out(a6_wr[863]), .rdlo_out(a6_wr[895]));
			radix2 #(.width(width)) rd_st5_896  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[896]), .rdlo_in(a5_wr[928]),  .coef_in(coef[0]), .rdup_out(a6_wr[896]), .rdlo_out(a6_wr[928]));
			radix2 #(.width(width)) rd_st5_897  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[897]), .rdlo_in(a5_wr[929]),  .coef_in(coef[32]), .rdup_out(a6_wr[897]), .rdlo_out(a6_wr[929]));
			radix2 #(.width(width)) rd_st5_898  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[898]), .rdlo_in(a5_wr[930]),  .coef_in(coef[64]), .rdup_out(a6_wr[898]), .rdlo_out(a6_wr[930]));
			radix2 #(.width(width)) rd_st5_899  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[899]), .rdlo_in(a5_wr[931]),  .coef_in(coef[96]), .rdup_out(a6_wr[899]), .rdlo_out(a6_wr[931]));
			radix2 #(.width(width)) rd_st5_900  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[900]), .rdlo_in(a5_wr[932]),  .coef_in(coef[128]), .rdup_out(a6_wr[900]), .rdlo_out(a6_wr[932]));
			radix2 #(.width(width)) rd_st5_901  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[901]), .rdlo_in(a5_wr[933]),  .coef_in(coef[160]), .rdup_out(a6_wr[901]), .rdlo_out(a6_wr[933]));
			radix2 #(.width(width)) rd_st5_902  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[902]), .rdlo_in(a5_wr[934]),  .coef_in(coef[192]), .rdup_out(a6_wr[902]), .rdlo_out(a6_wr[934]));
			radix2 #(.width(width)) rd_st5_903  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[903]), .rdlo_in(a5_wr[935]),  .coef_in(coef[224]), .rdup_out(a6_wr[903]), .rdlo_out(a6_wr[935]));
			radix2 #(.width(width)) rd_st5_904  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[904]), .rdlo_in(a5_wr[936]),  .coef_in(coef[256]), .rdup_out(a6_wr[904]), .rdlo_out(a6_wr[936]));
			radix2 #(.width(width)) rd_st5_905  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[905]), .rdlo_in(a5_wr[937]),  .coef_in(coef[288]), .rdup_out(a6_wr[905]), .rdlo_out(a6_wr[937]));
			radix2 #(.width(width)) rd_st5_906  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[906]), .rdlo_in(a5_wr[938]),  .coef_in(coef[320]), .rdup_out(a6_wr[906]), .rdlo_out(a6_wr[938]));
			radix2 #(.width(width)) rd_st5_907  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[907]), .rdlo_in(a5_wr[939]),  .coef_in(coef[352]), .rdup_out(a6_wr[907]), .rdlo_out(a6_wr[939]));
			radix2 #(.width(width)) rd_st5_908  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[908]), .rdlo_in(a5_wr[940]),  .coef_in(coef[384]), .rdup_out(a6_wr[908]), .rdlo_out(a6_wr[940]));
			radix2 #(.width(width)) rd_st5_909  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[909]), .rdlo_in(a5_wr[941]),  .coef_in(coef[416]), .rdup_out(a6_wr[909]), .rdlo_out(a6_wr[941]));
			radix2 #(.width(width)) rd_st5_910  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[910]), .rdlo_in(a5_wr[942]),  .coef_in(coef[448]), .rdup_out(a6_wr[910]), .rdlo_out(a6_wr[942]));
			radix2 #(.width(width)) rd_st5_911  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[911]), .rdlo_in(a5_wr[943]),  .coef_in(coef[480]), .rdup_out(a6_wr[911]), .rdlo_out(a6_wr[943]));
			radix2 #(.width(width)) rd_st5_912  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[912]), .rdlo_in(a5_wr[944]),  .coef_in(coef[512]), .rdup_out(a6_wr[912]), .rdlo_out(a6_wr[944]));
			radix2 #(.width(width)) rd_st5_913  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[913]), .rdlo_in(a5_wr[945]),  .coef_in(coef[544]), .rdup_out(a6_wr[913]), .rdlo_out(a6_wr[945]));
			radix2 #(.width(width)) rd_st5_914  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[914]), .rdlo_in(a5_wr[946]),  .coef_in(coef[576]), .rdup_out(a6_wr[914]), .rdlo_out(a6_wr[946]));
			radix2 #(.width(width)) rd_st5_915  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[915]), .rdlo_in(a5_wr[947]),  .coef_in(coef[608]), .rdup_out(a6_wr[915]), .rdlo_out(a6_wr[947]));
			radix2 #(.width(width)) rd_st5_916  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[916]), .rdlo_in(a5_wr[948]),  .coef_in(coef[640]), .rdup_out(a6_wr[916]), .rdlo_out(a6_wr[948]));
			radix2 #(.width(width)) rd_st5_917  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[917]), .rdlo_in(a5_wr[949]),  .coef_in(coef[672]), .rdup_out(a6_wr[917]), .rdlo_out(a6_wr[949]));
			radix2 #(.width(width)) rd_st5_918  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[918]), .rdlo_in(a5_wr[950]),  .coef_in(coef[704]), .rdup_out(a6_wr[918]), .rdlo_out(a6_wr[950]));
			radix2 #(.width(width)) rd_st5_919  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[919]), .rdlo_in(a5_wr[951]),  .coef_in(coef[736]), .rdup_out(a6_wr[919]), .rdlo_out(a6_wr[951]));
			radix2 #(.width(width)) rd_st5_920  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[920]), .rdlo_in(a5_wr[952]),  .coef_in(coef[768]), .rdup_out(a6_wr[920]), .rdlo_out(a6_wr[952]));
			radix2 #(.width(width)) rd_st5_921  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[921]), .rdlo_in(a5_wr[953]),  .coef_in(coef[800]), .rdup_out(a6_wr[921]), .rdlo_out(a6_wr[953]));
			radix2 #(.width(width)) rd_st5_922  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[922]), .rdlo_in(a5_wr[954]),  .coef_in(coef[832]), .rdup_out(a6_wr[922]), .rdlo_out(a6_wr[954]));
			radix2 #(.width(width)) rd_st5_923  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[923]), .rdlo_in(a5_wr[955]),  .coef_in(coef[864]), .rdup_out(a6_wr[923]), .rdlo_out(a6_wr[955]));
			radix2 #(.width(width)) rd_st5_924  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[924]), .rdlo_in(a5_wr[956]),  .coef_in(coef[896]), .rdup_out(a6_wr[924]), .rdlo_out(a6_wr[956]));
			radix2 #(.width(width)) rd_st5_925  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[925]), .rdlo_in(a5_wr[957]),  .coef_in(coef[928]), .rdup_out(a6_wr[925]), .rdlo_out(a6_wr[957]));
			radix2 #(.width(width)) rd_st5_926  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[926]), .rdlo_in(a5_wr[958]),  .coef_in(coef[960]), .rdup_out(a6_wr[926]), .rdlo_out(a6_wr[958]));
			radix2 #(.width(width)) rd_st5_927  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[927]), .rdlo_in(a5_wr[959]),  .coef_in(coef[992]), .rdup_out(a6_wr[927]), .rdlo_out(a6_wr[959]));
			radix2 #(.width(width)) rd_st5_960  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[960]), .rdlo_in(a5_wr[992]),  .coef_in(coef[0]), .rdup_out(a6_wr[960]), .rdlo_out(a6_wr[992]));
			radix2 #(.width(width)) rd_st5_961  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[961]), .rdlo_in(a5_wr[993]),  .coef_in(coef[32]), .rdup_out(a6_wr[961]), .rdlo_out(a6_wr[993]));
			radix2 #(.width(width)) rd_st5_962  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[962]), .rdlo_in(a5_wr[994]),  .coef_in(coef[64]), .rdup_out(a6_wr[962]), .rdlo_out(a6_wr[994]));
			radix2 #(.width(width)) rd_st5_963  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[963]), .rdlo_in(a5_wr[995]),  .coef_in(coef[96]), .rdup_out(a6_wr[963]), .rdlo_out(a6_wr[995]));
			radix2 #(.width(width)) rd_st5_964  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[964]), .rdlo_in(a5_wr[996]),  .coef_in(coef[128]), .rdup_out(a6_wr[964]), .rdlo_out(a6_wr[996]));
			radix2 #(.width(width)) rd_st5_965  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[965]), .rdlo_in(a5_wr[997]),  .coef_in(coef[160]), .rdup_out(a6_wr[965]), .rdlo_out(a6_wr[997]));
			radix2 #(.width(width)) rd_st5_966  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[966]), .rdlo_in(a5_wr[998]),  .coef_in(coef[192]), .rdup_out(a6_wr[966]), .rdlo_out(a6_wr[998]));
			radix2 #(.width(width)) rd_st5_967  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[967]), .rdlo_in(a5_wr[999]),  .coef_in(coef[224]), .rdup_out(a6_wr[967]), .rdlo_out(a6_wr[999]));
			radix2 #(.width(width)) rd_st5_968  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[968]), .rdlo_in(a5_wr[1000]),  .coef_in(coef[256]), .rdup_out(a6_wr[968]), .rdlo_out(a6_wr[1000]));
			radix2 #(.width(width)) rd_st5_969  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[969]), .rdlo_in(a5_wr[1001]),  .coef_in(coef[288]), .rdup_out(a6_wr[969]), .rdlo_out(a6_wr[1001]));
			radix2 #(.width(width)) rd_st5_970  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[970]), .rdlo_in(a5_wr[1002]),  .coef_in(coef[320]), .rdup_out(a6_wr[970]), .rdlo_out(a6_wr[1002]));
			radix2 #(.width(width)) rd_st5_971  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[971]), .rdlo_in(a5_wr[1003]),  .coef_in(coef[352]), .rdup_out(a6_wr[971]), .rdlo_out(a6_wr[1003]));
			radix2 #(.width(width)) rd_st5_972  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[972]), .rdlo_in(a5_wr[1004]),  .coef_in(coef[384]), .rdup_out(a6_wr[972]), .rdlo_out(a6_wr[1004]));
			radix2 #(.width(width)) rd_st5_973  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[973]), .rdlo_in(a5_wr[1005]),  .coef_in(coef[416]), .rdup_out(a6_wr[973]), .rdlo_out(a6_wr[1005]));
			radix2 #(.width(width)) rd_st5_974  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[974]), .rdlo_in(a5_wr[1006]),  .coef_in(coef[448]), .rdup_out(a6_wr[974]), .rdlo_out(a6_wr[1006]));
			radix2 #(.width(width)) rd_st5_975  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[975]), .rdlo_in(a5_wr[1007]),  .coef_in(coef[480]), .rdup_out(a6_wr[975]), .rdlo_out(a6_wr[1007]));
			radix2 #(.width(width)) rd_st5_976  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[976]), .rdlo_in(a5_wr[1008]),  .coef_in(coef[512]), .rdup_out(a6_wr[976]), .rdlo_out(a6_wr[1008]));
			radix2 #(.width(width)) rd_st5_977  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[977]), .rdlo_in(a5_wr[1009]),  .coef_in(coef[544]), .rdup_out(a6_wr[977]), .rdlo_out(a6_wr[1009]));
			radix2 #(.width(width)) rd_st5_978  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[978]), .rdlo_in(a5_wr[1010]),  .coef_in(coef[576]), .rdup_out(a6_wr[978]), .rdlo_out(a6_wr[1010]));
			radix2 #(.width(width)) rd_st5_979  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[979]), .rdlo_in(a5_wr[1011]),  .coef_in(coef[608]), .rdup_out(a6_wr[979]), .rdlo_out(a6_wr[1011]));
			radix2 #(.width(width)) rd_st5_980  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[980]), .rdlo_in(a5_wr[1012]),  .coef_in(coef[640]), .rdup_out(a6_wr[980]), .rdlo_out(a6_wr[1012]));
			radix2 #(.width(width)) rd_st5_981  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[981]), .rdlo_in(a5_wr[1013]),  .coef_in(coef[672]), .rdup_out(a6_wr[981]), .rdlo_out(a6_wr[1013]));
			radix2 #(.width(width)) rd_st5_982  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[982]), .rdlo_in(a5_wr[1014]),  .coef_in(coef[704]), .rdup_out(a6_wr[982]), .rdlo_out(a6_wr[1014]));
			radix2 #(.width(width)) rd_st5_983  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[983]), .rdlo_in(a5_wr[1015]),  .coef_in(coef[736]), .rdup_out(a6_wr[983]), .rdlo_out(a6_wr[1015]));
			radix2 #(.width(width)) rd_st5_984  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[984]), .rdlo_in(a5_wr[1016]),  .coef_in(coef[768]), .rdup_out(a6_wr[984]), .rdlo_out(a6_wr[1016]));
			radix2 #(.width(width)) rd_st5_985  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[985]), .rdlo_in(a5_wr[1017]),  .coef_in(coef[800]), .rdup_out(a6_wr[985]), .rdlo_out(a6_wr[1017]));
			radix2 #(.width(width)) rd_st5_986  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[986]), .rdlo_in(a5_wr[1018]),  .coef_in(coef[832]), .rdup_out(a6_wr[986]), .rdlo_out(a6_wr[1018]));
			radix2 #(.width(width)) rd_st5_987  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[987]), .rdlo_in(a5_wr[1019]),  .coef_in(coef[864]), .rdup_out(a6_wr[987]), .rdlo_out(a6_wr[1019]));
			radix2 #(.width(width)) rd_st5_988  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[988]), .rdlo_in(a5_wr[1020]),  .coef_in(coef[896]), .rdup_out(a6_wr[988]), .rdlo_out(a6_wr[1020]));
			radix2 #(.width(width)) rd_st5_989  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[989]), .rdlo_in(a5_wr[1021]),  .coef_in(coef[928]), .rdup_out(a6_wr[989]), .rdlo_out(a6_wr[1021]));
			radix2 #(.width(width)) rd_st5_990  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[990]), .rdlo_in(a5_wr[1022]),  .coef_in(coef[960]), .rdup_out(a6_wr[990]), .rdlo_out(a6_wr[1022]));
			radix2 #(.width(width)) rd_st5_991  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[991]), .rdlo_in(a5_wr[1023]),  .coef_in(coef[992]), .rdup_out(a6_wr[991]), .rdlo_out(a6_wr[1023]));
			radix2 #(.width(width)) rd_st5_1024  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1024]), .rdlo_in(a5_wr[1056]),  .coef_in(coef[0]), .rdup_out(a6_wr[1024]), .rdlo_out(a6_wr[1056]));
			radix2 #(.width(width)) rd_st5_1025  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1025]), .rdlo_in(a5_wr[1057]),  .coef_in(coef[32]), .rdup_out(a6_wr[1025]), .rdlo_out(a6_wr[1057]));
			radix2 #(.width(width)) rd_st5_1026  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1026]), .rdlo_in(a5_wr[1058]),  .coef_in(coef[64]), .rdup_out(a6_wr[1026]), .rdlo_out(a6_wr[1058]));
			radix2 #(.width(width)) rd_st5_1027  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1027]), .rdlo_in(a5_wr[1059]),  .coef_in(coef[96]), .rdup_out(a6_wr[1027]), .rdlo_out(a6_wr[1059]));
			radix2 #(.width(width)) rd_st5_1028  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1028]), .rdlo_in(a5_wr[1060]),  .coef_in(coef[128]), .rdup_out(a6_wr[1028]), .rdlo_out(a6_wr[1060]));
			radix2 #(.width(width)) rd_st5_1029  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1029]), .rdlo_in(a5_wr[1061]),  .coef_in(coef[160]), .rdup_out(a6_wr[1029]), .rdlo_out(a6_wr[1061]));
			radix2 #(.width(width)) rd_st5_1030  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1030]), .rdlo_in(a5_wr[1062]),  .coef_in(coef[192]), .rdup_out(a6_wr[1030]), .rdlo_out(a6_wr[1062]));
			radix2 #(.width(width)) rd_st5_1031  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1031]), .rdlo_in(a5_wr[1063]),  .coef_in(coef[224]), .rdup_out(a6_wr[1031]), .rdlo_out(a6_wr[1063]));
			radix2 #(.width(width)) rd_st5_1032  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1032]), .rdlo_in(a5_wr[1064]),  .coef_in(coef[256]), .rdup_out(a6_wr[1032]), .rdlo_out(a6_wr[1064]));
			radix2 #(.width(width)) rd_st5_1033  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1033]), .rdlo_in(a5_wr[1065]),  .coef_in(coef[288]), .rdup_out(a6_wr[1033]), .rdlo_out(a6_wr[1065]));
			radix2 #(.width(width)) rd_st5_1034  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1034]), .rdlo_in(a5_wr[1066]),  .coef_in(coef[320]), .rdup_out(a6_wr[1034]), .rdlo_out(a6_wr[1066]));
			radix2 #(.width(width)) rd_st5_1035  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1035]), .rdlo_in(a5_wr[1067]),  .coef_in(coef[352]), .rdup_out(a6_wr[1035]), .rdlo_out(a6_wr[1067]));
			radix2 #(.width(width)) rd_st5_1036  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1036]), .rdlo_in(a5_wr[1068]),  .coef_in(coef[384]), .rdup_out(a6_wr[1036]), .rdlo_out(a6_wr[1068]));
			radix2 #(.width(width)) rd_st5_1037  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1037]), .rdlo_in(a5_wr[1069]),  .coef_in(coef[416]), .rdup_out(a6_wr[1037]), .rdlo_out(a6_wr[1069]));
			radix2 #(.width(width)) rd_st5_1038  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1038]), .rdlo_in(a5_wr[1070]),  .coef_in(coef[448]), .rdup_out(a6_wr[1038]), .rdlo_out(a6_wr[1070]));
			radix2 #(.width(width)) rd_st5_1039  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1039]), .rdlo_in(a5_wr[1071]),  .coef_in(coef[480]), .rdup_out(a6_wr[1039]), .rdlo_out(a6_wr[1071]));
			radix2 #(.width(width)) rd_st5_1040  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1040]), .rdlo_in(a5_wr[1072]),  .coef_in(coef[512]), .rdup_out(a6_wr[1040]), .rdlo_out(a6_wr[1072]));
			radix2 #(.width(width)) rd_st5_1041  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1041]), .rdlo_in(a5_wr[1073]),  .coef_in(coef[544]), .rdup_out(a6_wr[1041]), .rdlo_out(a6_wr[1073]));
			radix2 #(.width(width)) rd_st5_1042  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1042]), .rdlo_in(a5_wr[1074]),  .coef_in(coef[576]), .rdup_out(a6_wr[1042]), .rdlo_out(a6_wr[1074]));
			radix2 #(.width(width)) rd_st5_1043  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1043]), .rdlo_in(a5_wr[1075]),  .coef_in(coef[608]), .rdup_out(a6_wr[1043]), .rdlo_out(a6_wr[1075]));
			radix2 #(.width(width)) rd_st5_1044  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1044]), .rdlo_in(a5_wr[1076]),  .coef_in(coef[640]), .rdup_out(a6_wr[1044]), .rdlo_out(a6_wr[1076]));
			radix2 #(.width(width)) rd_st5_1045  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1045]), .rdlo_in(a5_wr[1077]),  .coef_in(coef[672]), .rdup_out(a6_wr[1045]), .rdlo_out(a6_wr[1077]));
			radix2 #(.width(width)) rd_st5_1046  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1046]), .rdlo_in(a5_wr[1078]),  .coef_in(coef[704]), .rdup_out(a6_wr[1046]), .rdlo_out(a6_wr[1078]));
			radix2 #(.width(width)) rd_st5_1047  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1047]), .rdlo_in(a5_wr[1079]),  .coef_in(coef[736]), .rdup_out(a6_wr[1047]), .rdlo_out(a6_wr[1079]));
			radix2 #(.width(width)) rd_st5_1048  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1048]), .rdlo_in(a5_wr[1080]),  .coef_in(coef[768]), .rdup_out(a6_wr[1048]), .rdlo_out(a6_wr[1080]));
			radix2 #(.width(width)) rd_st5_1049  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1049]), .rdlo_in(a5_wr[1081]),  .coef_in(coef[800]), .rdup_out(a6_wr[1049]), .rdlo_out(a6_wr[1081]));
			radix2 #(.width(width)) rd_st5_1050  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1050]), .rdlo_in(a5_wr[1082]),  .coef_in(coef[832]), .rdup_out(a6_wr[1050]), .rdlo_out(a6_wr[1082]));
			radix2 #(.width(width)) rd_st5_1051  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1051]), .rdlo_in(a5_wr[1083]),  .coef_in(coef[864]), .rdup_out(a6_wr[1051]), .rdlo_out(a6_wr[1083]));
			radix2 #(.width(width)) rd_st5_1052  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1052]), .rdlo_in(a5_wr[1084]),  .coef_in(coef[896]), .rdup_out(a6_wr[1052]), .rdlo_out(a6_wr[1084]));
			radix2 #(.width(width)) rd_st5_1053  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1053]), .rdlo_in(a5_wr[1085]),  .coef_in(coef[928]), .rdup_out(a6_wr[1053]), .rdlo_out(a6_wr[1085]));
			radix2 #(.width(width)) rd_st5_1054  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1054]), .rdlo_in(a5_wr[1086]),  .coef_in(coef[960]), .rdup_out(a6_wr[1054]), .rdlo_out(a6_wr[1086]));
			radix2 #(.width(width)) rd_st5_1055  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1055]), .rdlo_in(a5_wr[1087]),  .coef_in(coef[992]), .rdup_out(a6_wr[1055]), .rdlo_out(a6_wr[1087]));
			radix2 #(.width(width)) rd_st5_1088  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1088]), .rdlo_in(a5_wr[1120]),  .coef_in(coef[0]), .rdup_out(a6_wr[1088]), .rdlo_out(a6_wr[1120]));
			radix2 #(.width(width)) rd_st5_1089  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1089]), .rdlo_in(a5_wr[1121]),  .coef_in(coef[32]), .rdup_out(a6_wr[1089]), .rdlo_out(a6_wr[1121]));
			radix2 #(.width(width)) rd_st5_1090  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1090]), .rdlo_in(a5_wr[1122]),  .coef_in(coef[64]), .rdup_out(a6_wr[1090]), .rdlo_out(a6_wr[1122]));
			radix2 #(.width(width)) rd_st5_1091  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1091]), .rdlo_in(a5_wr[1123]),  .coef_in(coef[96]), .rdup_out(a6_wr[1091]), .rdlo_out(a6_wr[1123]));
			radix2 #(.width(width)) rd_st5_1092  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1092]), .rdlo_in(a5_wr[1124]),  .coef_in(coef[128]), .rdup_out(a6_wr[1092]), .rdlo_out(a6_wr[1124]));
			radix2 #(.width(width)) rd_st5_1093  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1093]), .rdlo_in(a5_wr[1125]),  .coef_in(coef[160]), .rdup_out(a6_wr[1093]), .rdlo_out(a6_wr[1125]));
			radix2 #(.width(width)) rd_st5_1094  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1094]), .rdlo_in(a5_wr[1126]),  .coef_in(coef[192]), .rdup_out(a6_wr[1094]), .rdlo_out(a6_wr[1126]));
			radix2 #(.width(width)) rd_st5_1095  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1095]), .rdlo_in(a5_wr[1127]),  .coef_in(coef[224]), .rdup_out(a6_wr[1095]), .rdlo_out(a6_wr[1127]));
			radix2 #(.width(width)) rd_st5_1096  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1096]), .rdlo_in(a5_wr[1128]),  .coef_in(coef[256]), .rdup_out(a6_wr[1096]), .rdlo_out(a6_wr[1128]));
			radix2 #(.width(width)) rd_st5_1097  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1097]), .rdlo_in(a5_wr[1129]),  .coef_in(coef[288]), .rdup_out(a6_wr[1097]), .rdlo_out(a6_wr[1129]));
			radix2 #(.width(width)) rd_st5_1098  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1098]), .rdlo_in(a5_wr[1130]),  .coef_in(coef[320]), .rdup_out(a6_wr[1098]), .rdlo_out(a6_wr[1130]));
			radix2 #(.width(width)) rd_st5_1099  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1099]), .rdlo_in(a5_wr[1131]),  .coef_in(coef[352]), .rdup_out(a6_wr[1099]), .rdlo_out(a6_wr[1131]));
			radix2 #(.width(width)) rd_st5_1100  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1100]), .rdlo_in(a5_wr[1132]),  .coef_in(coef[384]), .rdup_out(a6_wr[1100]), .rdlo_out(a6_wr[1132]));
			radix2 #(.width(width)) rd_st5_1101  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1101]), .rdlo_in(a5_wr[1133]),  .coef_in(coef[416]), .rdup_out(a6_wr[1101]), .rdlo_out(a6_wr[1133]));
			radix2 #(.width(width)) rd_st5_1102  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1102]), .rdlo_in(a5_wr[1134]),  .coef_in(coef[448]), .rdup_out(a6_wr[1102]), .rdlo_out(a6_wr[1134]));
			radix2 #(.width(width)) rd_st5_1103  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1103]), .rdlo_in(a5_wr[1135]),  .coef_in(coef[480]), .rdup_out(a6_wr[1103]), .rdlo_out(a6_wr[1135]));
			radix2 #(.width(width)) rd_st5_1104  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1104]), .rdlo_in(a5_wr[1136]),  .coef_in(coef[512]), .rdup_out(a6_wr[1104]), .rdlo_out(a6_wr[1136]));
			radix2 #(.width(width)) rd_st5_1105  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1105]), .rdlo_in(a5_wr[1137]),  .coef_in(coef[544]), .rdup_out(a6_wr[1105]), .rdlo_out(a6_wr[1137]));
			radix2 #(.width(width)) rd_st5_1106  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1106]), .rdlo_in(a5_wr[1138]),  .coef_in(coef[576]), .rdup_out(a6_wr[1106]), .rdlo_out(a6_wr[1138]));
			radix2 #(.width(width)) rd_st5_1107  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1107]), .rdlo_in(a5_wr[1139]),  .coef_in(coef[608]), .rdup_out(a6_wr[1107]), .rdlo_out(a6_wr[1139]));
			radix2 #(.width(width)) rd_st5_1108  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1108]), .rdlo_in(a5_wr[1140]),  .coef_in(coef[640]), .rdup_out(a6_wr[1108]), .rdlo_out(a6_wr[1140]));
			radix2 #(.width(width)) rd_st5_1109  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1109]), .rdlo_in(a5_wr[1141]),  .coef_in(coef[672]), .rdup_out(a6_wr[1109]), .rdlo_out(a6_wr[1141]));
			radix2 #(.width(width)) rd_st5_1110  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1110]), .rdlo_in(a5_wr[1142]),  .coef_in(coef[704]), .rdup_out(a6_wr[1110]), .rdlo_out(a6_wr[1142]));
			radix2 #(.width(width)) rd_st5_1111  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1111]), .rdlo_in(a5_wr[1143]),  .coef_in(coef[736]), .rdup_out(a6_wr[1111]), .rdlo_out(a6_wr[1143]));
			radix2 #(.width(width)) rd_st5_1112  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1112]), .rdlo_in(a5_wr[1144]),  .coef_in(coef[768]), .rdup_out(a6_wr[1112]), .rdlo_out(a6_wr[1144]));
			radix2 #(.width(width)) rd_st5_1113  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1113]), .rdlo_in(a5_wr[1145]),  .coef_in(coef[800]), .rdup_out(a6_wr[1113]), .rdlo_out(a6_wr[1145]));
			radix2 #(.width(width)) rd_st5_1114  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1114]), .rdlo_in(a5_wr[1146]),  .coef_in(coef[832]), .rdup_out(a6_wr[1114]), .rdlo_out(a6_wr[1146]));
			radix2 #(.width(width)) rd_st5_1115  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1115]), .rdlo_in(a5_wr[1147]),  .coef_in(coef[864]), .rdup_out(a6_wr[1115]), .rdlo_out(a6_wr[1147]));
			radix2 #(.width(width)) rd_st5_1116  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1116]), .rdlo_in(a5_wr[1148]),  .coef_in(coef[896]), .rdup_out(a6_wr[1116]), .rdlo_out(a6_wr[1148]));
			radix2 #(.width(width)) rd_st5_1117  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1117]), .rdlo_in(a5_wr[1149]),  .coef_in(coef[928]), .rdup_out(a6_wr[1117]), .rdlo_out(a6_wr[1149]));
			radix2 #(.width(width)) rd_st5_1118  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1118]), .rdlo_in(a5_wr[1150]),  .coef_in(coef[960]), .rdup_out(a6_wr[1118]), .rdlo_out(a6_wr[1150]));
			radix2 #(.width(width)) rd_st5_1119  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1119]), .rdlo_in(a5_wr[1151]),  .coef_in(coef[992]), .rdup_out(a6_wr[1119]), .rdlo_out(a6_wr[1151]));
			radix2 #(.width(width)) rd_st5_1152  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1152]), .rdlo_in(a5_wr[1184]),  .coef_in(coef[0]), .rdup_out(a6_wr[1152]), .rdlo_out(a6_wr[1184]));
			radix2 #(.width(width)) rd_st5_1153  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1153]), .rdlo_in(a5_wr[1185]),  .coef_in(coef[32]), .rdup_out(a6_wr[1153]), .rdlo_out(a6_wr[1185]));
			radix2 #(.width(width)) rd_st5_1154  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1154]), .rdlo_in(a5_wr[1186]),  .coef_in(coef[64]), .rdup_out(a6_wr[1154]), .rdlo_out(a6_wr[1186]));
			radix2 #(.width(width)) rd_st5_1155  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1155]), .rdlo_in(a5_wr[1187]),  .coef_in(coef[96]), .rdup_out(a6_wr[1155]), .rdlo_out(a6_wr[1187]));
			radix2 #(.width(width)) rd_st5_1156  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1156]), .rdlo_in(a5_wr[1188]),  .coef_in(coef[128]), .rdup_out(a6_wr[1156]), .rdlo_out(a6_wr[1188]));
			radix2 #(.width(width)) rd_st5_1157  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1157]), .rdlo_in(a5_wr[1189]),  .coef_in(coef[160]), .rdup_out(a6_wr[1157]), .rdlo_out(a6_wr[1189]));
			radix2 #(.width(width)) rd_st5_1158  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1158]), .rdlo_in(a5_wr[1190]),  .coef_in(coef[192]), .rdup_out(a6_wr[1158]), .rdlo_out(a6_wr[1190]));
			radix2 #(.width(width)) rd_st5_1159  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1159]), .rdlo_in(a5_wr[1191]),  .coef_in(coef[224]), .rdup_out(a6_wr[1159]), .rdlo_out(a6_wr[1191]));
			radix2 #(.width(width)) rd_st5_1160  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1160]), .rdlo_in(a5_wr[1192]),  .coef_in(coef[256]), .rdup_out(a6_wr[1160]), .rdlo_out(a6_wr[1192]));
			radix2 #(.width(width)) rd_st5_1161  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1161]), .rdlo_in(a5_wr[1193]),  .coef_in(coef[288]), .rdup_out(a6_wr[1161]), .rdlo_out(a6_wr[1193]));
			radix2 #(.width(width)) rd_st5_1162  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1162]), .rdlo_in(a5_wr[1194]),  .coef_in(coef[320]), .rdup_out(a6_wr[1162]), .rdlo_out(a6_wr[1194]));
			radix2 #(.width(width)) rd_st5_1163  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1163]), .rdlo_in(a5_wr[1195]),  .coef_in(coef[352]), .rdup_out(a6_wr[1163]), .rdlo_out(a6_wr[1195]));
			radix2 #(.width(width)) rd_st5_1164  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1164]), .rdlo_in(a5_wr[1196]),  .coef_in(coef[384]), .rdup_out(a6_wr[1164]), .rdlo_out(a6_wr[1196]));
			radix2 #(.width(width)) rd_st5_1165  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1165]), .rdlo_in(a5_wr[1197]),  .coef_in(coef[416]), .rdup_out(a6_wr[1165]), .rdlo_out(a6_wr[1197]));
			radix2 #(.width(width)) rd_st5_1166  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1166]), .rdlo_in(a5_wr[1198]),  .coef_in(coef[448]), .rdup_out(a6_wr[1166]), .rdlo_out(a6_wr[1198]));
			radix2 #(.width(width)) rd_st5_1167  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1167]), .rdlo_in(a5_wr[1199]),  .coef_in(coef[480]), .rdup_out(a6_wr[1167]), .rdlo_out(a6_wr[1199]));
			radix2 #(.width(width)) rd_st5_1168  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1168]), .rdlo_in(a5_wr[1200]),  .coef_in(coef[512]), .rdup_out(a6_wr[1168]), .rdlo_out(a6_wr[1200]));
			radix2 #(.width(width)) rd_st5_1169  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1169]), .rdlo_in(a5_wr[1201]),  .coef_in(coef[544]), .rdup_out(a6_wr[1169]), .rdlo_out(a6_wr[1201]));
			radix2 #(.width(width)) rd_st5_1170  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1170]), .rdlo_in(a5_wr[1202]),  .coef_in(coef[576]), .rdup_out(a6_wr[1170]), .rdlo_out(a6_wr[1202]));
			radix2 #(.width(width)) rd_st5_1171  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1171]), .rdlo_in(a5_wr[1203]),  .coef_in(coef[608]), .rdup_out(a6_wr[1171]), .rdlo_out(a6_wr[1203]));
			radix2 #(.width(width)) rd_st5_1172  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1172]), .rdlo_in(a5_wr[1204]),  .coef_in(coef[640]), .rdup_out(a6_wr[1172]), .rdlo_out(a6_wr[1204]));
			radix2 #(.width(width)) rd_st5_1173  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1173]), .rdlo_in(a5_wr[1205]),  .coef_in(coef[672]), .rdup_out(a6_wr[1173]), .rdlo_out(a6_wr[1205]));
			radix2 #(.width(width)) rd_st5_1174  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1174]), .rdlo_in(a5_wr[1206]),  .coef_in(coef[704]), .rdup_out(a6_wr[1174]), .rdlo_out(a6_wr[1206]));
			radix2 #(.width(width)) rd_st5_1175  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1175]), .rdlo_in(a5_wr[1207]),  .coef_in(coef[736]), .rdup_out(a6_wr[1175]), .rdlo_out(a6_wr[1207]));
			radix2 #(.width(width)) rd_st5_1176  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1176]), .rdlo_in(a5_wr[1208]),  .coef_in(coef[768]), .rdup_out(a6_wr[1176]), .rdlo_out(a6_wr[1208]));
			radix2 #(.width(width)) rd_st5_1177  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1177]), .rdlo_in(a5_wr[1209]),  .coef_in(coef[800]), .rdup_out(a6_wr[1177]), .rdlo_out(a6_wr[1209]));
			radix2 #(.width(width)) rd_st5_1178  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1178]), .rdlo_in(a5_wr[1210]),  .coef_in(coef[832]), .rdup_out(a6_wr[1178]), .rdlo_out(a6_wr[1210]));
			radix2 #(.width(width)) rd_st5_1179  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1179]), .rdlo_in(a5_wr[1211]),  .coef_in(coef[864]), .rdup_out(a6_wr[1179]), .rdlo_out(a6_wr[1211]));
			radix2 #(.width(width)) rd_st5_1180  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1180]), .rdlo_in(a5_wr[1212]),  .coef_in(coef[896]), .rdup_out(a6_wr[1180]), .rdlo_out(a6_wr[1212]));
			radix2 #(.width(width)) rd_st5_1181  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1181]), .rdlo_in(a5_wr[1213]),  .coef_in(coef[928]), .rdup_out(a6_wr[1181]), .rdlo_out(a6_wr[1213]));
			radix2 #(.width(width)) rd_st5_1182  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1182]), .rdlo_in(a5_wr[1214]),  .coef_in(coef[960]), .rdup_out(a6_wr[1182]), .rdlo_out(a6_wr[1214]));
			radix2 #(.width(width)) rd_st5_1183  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1183]), .rdlo_in(a5_wr[1215]),  .coef_in(coef[992]), .rdup_out(a6_wr[1183]), .rdlo_out(a6_wr[1215]));
			radix2 #(.width(width)) rd_st5_1216  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1216]), .rdlo_in(a5_wr[1248]),  .coef_in(coef[0]), .rdup_out(a6_wr[1216]), .rdlo_out(a6_wr[1248]));
			radix2 #(.width(width)) rd_st5_1217  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1217]), .rdlo_in(a5_wr[1249]),  .coef_in(coef[32]), .rdup_out(a6_wr[1217]), .rdlo_out(a6_wr[1249]));
			radix2 #(.width(width)) rd_st5_1218  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1218]), .rdlo_in(a5_wr[1250]),  .coef_in(coef[64]), .rdup_out(a6_wr[1218]), .rdlo_out(a6_wr[1250]));
			radix2 #(.width(width)) rd_st5_1219  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1219]), .rdlo_in(a5_wr[1251]),  .coef_in(coef[96]), .rdup_out(a6_wr[1219]), .rdlo_out(a6_wr[1251]));
			radix2 #(.width(width)) rd_st5_1220  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1220]), .rdlo_in(a5_wr[1252]),  .coef_in(coef[128]), .rdup_out(a6_wr[1220]), .rdlo_out(a6_wr[1252]));
			radix2 #(.width(width)) rd_st5_1221  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1221]), .rdlo_in(a5_wr[1253]),  .coef_in(coef[160]), .rdup_out(a6_wr[1221]), .rdlo_out(a6_wr[1253]));
			radix2 #(.width(width)) rd_st5_1222  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1222]), .rdlo_in(a5_wr[1254]),  .coef_in(coef[192]), .rdup_out(a6_wr[1222]), .rdlo_out(a6_wr[1254]));
			radix2 #(.width(width)) rd_st5_1223  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1223]), .rdlo_in(a5_wr[1255]),  .coef_in(coef[224]), .rdup_out(a6_wr[1223]), .rdlo_out(a6_wr[1255]));
			radix2 #(.width(width)) rd_st5_1224  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1224]), .rdlo_in(a5_wr[1256]),  .coef_in(coef[256]), .rdup_out(a6_wr[1224]), .rdlo_out(a6_wr[1256]));
			radix2 #(.width(width)) rd_st5_1225  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1225]), .rdlo_in(a5_wr[1257]),  .coef_in(coef[288]), .rdup_out(a6_wr[1225]), .rdlo_out(a6_wr[1257]));
			radix2 #(.width(width)) rd_st5_1226  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1226]), .rdlo_in(a5_wr[1258]),  .coef_in(coef[320]), .rdup_out(a6_wr[1226]), .rdlo_out(a6_wr[1258]));
			radix2 #(.width(width)) rd_st5_1227  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1227]), .rdlo_in(a5_wr[1259]),  .coef_in(coef[352]), .rdup_out(a6_wr[1227]), .rdlo_out(a6_wr[1259]));
			radix2 #(.width(width)) rd_st5_1228  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1228]), .rdlo_in(a5_wr[1260]),  .coef_in(coef[384]), .rdup_out(a6_wr[1228]), .rdlo_out(a6_wr[1260]));
			radix2 #(.width(width)) rd_st5_1229  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1229]), .rdlo_in(a5_wr[1261]),  .coef_in(coef[416]), .rdup_out(a6_wr[1229]), .rdlo_out(a6_wr[1261]));
			radix2 #(.width(width)) rd_st5_1230  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1230]), .rdlo_in(a5_wr[1262]),  .coef_in(coef[448]), .rdup_out(a6_wr[1230]), .rdlo_out(a6_wr[1262]));
			radix2 #(.width(width)) rd_st5_1231  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1231]), .rdlo_in(a5_wr[1263]),  .coef_in(coef[480]), .rdup_out(a6_wr[1231]), .rdlo_out(a6_wr[1263]));
			radix2 #(.width(width)) rd_st5_1232  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1232]), .rdlo_in(a5_wr[1264]),  .coef_in(coef[512]), .rdup_out(a6_wr[1232]), .rdlo_out(a6_wr[1264]));
			radix2 #(.width(width)) rd_st5_1233  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1233]), .rdlo_in(a5_wr[1265]),  .coef_in(coef[544]), .rdup_out(a6_wr[1233]), .rdlo_out(a6_wr[1265]));
			radix2 #(.width(width)) rd_st5_1234  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1234]), .rdlo_in(a5_wr[1266]),  .coef_in(coef[576]), .rdup_out(a6_wr[1234]), .rdlo_out(a6_wr[1266]));
			radix2 #(.width(width)) rd_st5_1235  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1235]), .rdlo_in(a5_wr[1267]),  .coef_in(coef[608]), .rdup_out(a6_wr[1235]), .rdlo_out(a6_wr[1267]));
			radix2 #(.width(width)) rd_st5_1236  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1236]), .rdlo_in(a5_wr[1268]),  .coef_in(coef[640]), .rdup_out(a6_wr[1236]), .rdlo_out(a6_wr[1268]));
			radix2 #(.width(width)) rd_st5_1237  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1237]), .rdlo_in(a5_wr[1269]),  .coef_in(coef[672]), .rdup_out(a6_wr[1237]), .rdlo_out(a6_wr[1269]));
			radix2 #(.width(width)) rd_st5_1238  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1238]), .rdlo_in(a5_wr[1270]),  .coef_in(coef[704]), .rdup_out(a6_wr[1238]), .rdlo_out(a6_wr[1270]));
			radix2 #(.width(width)) rd_st5_1239  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1239]), .rdlo_in(a5_wr[1271]),  .coef_in(coef[736]), .rdup_out(a6_wr[1239]), .rdlo_out(a6_wr[1271]));
			radix2 #(.width(width)) rd_st5_1240  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1240]), .rdlo_in(a5_wr[1272]),  .coef_in(coef[768]), .rdup_out(a6_wr[1240]), .rdlo_out(a6_wr[1272]));
			radix2 #(.width(width)) rd_st5_1241  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1241]), .rdlo_in(a5_wr[1273]),  .coef_in(coef[800]), .rdup_out(a6_wr[1241]), .rdlo_out(a6_wr[1273]));
			radix2 #(.width(width)) rd_st5_1242  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1242]), .rdlo_in(a5_wr[1274]),  .coef_in(coef[832]), .rdup_out(a6_wr[1242]), .rdlo_out(a6_wr[1274]));
			radix2 #(.width(width)) rd_st5_1243  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1243]), .rdlo_in(a5_wr[1275]),  .coef_in(coef[864]), .rdup_out(a6_wr[1243]), .rdlo_out(a6_wr[1275]));
			radix2 #(.width(width)) rd_st5_1244  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1244]), .rdlo_in(a5_wr[1276]),  .coef_in(coef[896]), .rdup_out(a6_wr[1244]), .rdlo_out(a6_wr[1276]));
			radix2 #(.width(width)) rd_st5_1245  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1245]), .rdlo_in(a5_wr[1277]),  .coef_in(coef[928]), .rdup_out(a6_wr[1245]), .rdlo_out(a6_wr[1277]));
			radix2 #(.width(width)) rd_st5_1246  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1246]), .rdlo_in(a5_wr[1278]),  .coef_in(coef[960]), .rdup_out(a6_wr[1246]), .rdlo_out(a6_wr[1278]));
			radix2 #(.width(width)) rd_st5_1247  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1247]), .rdlo_in(a5_wr[1279]),  .coef_in(coef[992]), .rdup_out(a6_wr[1247]), .rdlo_out(a6_wr[1279]));
			radix2 #(.width(width)) rd_st5_1280  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1280]), .rdlo_in(a5_wr[1312]),  .coef_in(coef[0]), .rdup_out(a6_wr[1280]), .rdlo_out(a6_wr[1312]));
			radix2 #(.width(width)) rd_st5_1281  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1281]), .rdlo_in(a5_wr[1313]),  .coef_in(coef[32]), .rdup_out(a6_wr[1281]), .rdlo_out(a6_wr[1313]));
			radix2 #(.width(width)) rd_st5_1282  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1282]), .rdlo_in(a5_wr[1314]),  .coef_in(coef[64]), .rdup_out(a6_wr[1282]), .rdlo_out(a6_wr[1314]));
			radix2 #(.width(width)) rd_st5_1283  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1283]), .rdlo_in(a5_wr[1315]),  .coef_in(coef[96]), .rdup_out(a6_wr[1283]), .rdlo_out(a6_wr[1315]));
			radix2 #(.width(width)) rd_st5_1284  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1284]), .rdlo_in(a5_wr[1316]),  .coef_in(coef[128]), .rdup_out(a6_wr[1284]), .rdlo_out(a6_wr[1316]));
			radix2 #(.width(width)) rd_st5_1285  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1285]), .rdlo_in(a5_wr[1317]),  .coef_in(coef[160]), .rdup_out(a6_wr[1285]), .rdlo_out(a6_wr[1317]));
			radix2 #(.width(width)) rd_st5_1286  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1286]), .rdlo_in(a5_wr[1318]),  .coef_in(coef[192]), .rdup_out(a6_wr[1286]), .rdlo_out(a6_wr[1318]));
			radix2 #(.width(width)) rd_st5_1287  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1287]), .rdlo_in(a5_wr[1319]),  .coef_in(coef[224]), .rdup_out(a6_wr[1287]), .rdlo_out(a6_wr[1319]));
			radix2 #(.width(width)) rd_st5_1288  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1288]), .rdlo_in(a5_wr[1320]),  .coef_in(coef[256]), .rdup_out(a6_wr[1288]), .rdlo_out(a6_wr[1320]));
			radix2 #(.width(width)) rd_st5_1289  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1289]), .rdlo_in(a5_wr[1321]),  .coef_in(coef[288]), .rdup_out(a6_wr[1289]), .rdlo_out(a6_wr[1321]));
			radix2 #(.width(width)) rd_st5_1290  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1290]), .rdlo_in(a5_wr[1322]),  .coef_in(coef[320]), .rdup_out(a6_wr[1290]), .rdlo_out(a6_wr[1322]));
			radix2 #(.width(width)) rd_st5_1291  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1291]), .rdlo_in(a5_wr[1323]),  .coef_in(coef[352]), .rdup_out(a6_wr[1291]), .rdlo_out(a6_wr[1323]));
			radix2 #(.width(width)) rd_st5_1292  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1292]), .rdlo_in(a5_wr[1324]),  .coef_in(coef[384]), .rdup_out(a6_wr[1292]), .rdlo_out(a6_wr[1324]));
			radix2 #(.width(width)) rd_st5_1293  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1293]), .rdlo_in(a5_wr[1325]),  .coef_in(coef[416]), .rdup_out(a6_wr[1293]), .rdlo_out(a6_wr[1325]));
			radix2 #(.width(width)) rd_st5_1294  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1294]), .rdlo_in(a5_wr[1326]),  .coef_in(coef[448]), .rdup_out(a6_wr[1294]), .rdlo_out(a6_wr[1326]));
			radix2 #(.width(width)) rd_st5_1295  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1295]), .rdlo_in(a5_wr[1327]),  .coef_in(coef[480]), .rdup_out(a6_wr[1295]), .rdlo_out(a6_wr[1327]));
			radix2 #(.width(width)) rd_st5_1296  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1296]), .rdlo_in(a5_wr[1328]),  .coef_in(coef[512]), .rdup_out(a6_wr[1296]), .rdlo_out(a6_wr[1328]));
			radix2 #(.width(width)) rd_st5_1297  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1297]), .rdlo_in(a5_wr[1329]),  .coef_in(coef[544]), .rdup_out(a6_wr[1297]), .rdlo_out(a6_wr[1329]));
			radix2 #(.width(width)) rd_st5_1298  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1298]), .rdlo_in(a5_wr[1330]),  .coef_in(coef[576]), .rdup_out(a6_wr[1298]), .rdlo_out(a6_wr[1330]));
			radix2 #(.width(width)) rd_st5_1299  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1299]), .rdlo_in(a5_wr[1331]),  .coef_in(coef[608]), .rdup_out(a6_wr[1299]), .rdlo_out(a6_wr[1331]));
			radix2 #(.width(width)) rd_st5_1300  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1300]), .rdlo_in(a5_wr[1332]),  .coef_in(coef[640]), .rdup_out(a6_wr[1300]), .rdlo_out(a6_wr[1332]));
			radix2 #(.width(width)) rd_st5_1301  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1301]), .rdlo_in(a5_wr[1333]),  .coef_in(coef[672]), .rdup_out(a6_wr[1301]), .rdlo_out(a6_wr[1333]));
			radix2 #(.width(width)) rd_st5_1302  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1302]), .rdlo_in(a5_wr[1334]),  .coef_in(coef[704]), .rdup_out(a6_wr[1302]), .rdlo_out(a6_wr[1334]));
			radix2 #(.width(width)) rd_st5_1303  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1303]), .rdlo_in(a5_wr[1335]),  .coef_in(coef[736]), .rdup_out(a6_wr[1303]), .rdlo_out(a6_wr[1335]));
			radix2 #(.width(width)) rd_st5_1304  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1304]), .rdlo_in(a5_wr[1336]),  .coef_in(coef[768]), .rdup_out(a6_wr[1304]), .rdlo_out(a6_wr[1336]));
			radix2 #(.width(width)) rd_st5_1305  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1305]), .rdlo_in(a5_wr[1337]),  .coef_in(coef[800]), .rdup_out(a6_wr[1305]), .rdlo_out(a6_wr[1337]));
			radix2 #(.width(width)) rd_st5_1306  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1306]), .rdlo_in(a5_wr[1338]),  .coef_in(coef[832]), .rdup_out(a6_wr[1306]), .rdlo_out(a6_wr[1338]));
			radix2 #(.width(width)) rd_st5_1307  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1307]), .rdlo_in(a5_wr[1339]),  .coef_in(coef[864]), .rdup_out(a6_wr[1307]), .rdlo_out(a6_wr[1339]));
			radix2 #(.width(width)) rd_st5_1308  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1308]), .rdlo_in(a5_wr[1340]),  .coef_in(coef[896]), .rdup_out(a6_wr[1308]), .rdlo_out(a6_wr[1340]));
			radix2 #(.width(width)) rd_st5_1309  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1309]), .rdlo_in(a5_wr[1341]),  .coef_in(coef[928]), .rdup_out(a6_wr[1309]), .rdlo_out(a6_wr[1341]));
			radix2 #(.width(width)) rd_st5_1310  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1310]), .rdlo_in(a5_wr[1342]),  .coef_in(coef[960]), .rdup_out(a6_wr[1310]), .rdlo_out(a6_wr[1342]));
			radix2 #(.width(width)) rd_st5_1311  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1311]), .rdlo_in(a5_wr[1343]),  .coef_in(coef[992]), .rdup_out(a6_wr[1311]), .rdlo_out(a6_wr[1343]));
			radix2 #(.width(width)) rd_st5_1344  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1344]), .rdlo_in(a5_wr[1376]),  .coef_in(coef[0]), .rdup_out(a6_wr[1344]), .rdlo_out(a6_wr[1376]));
			radix2 #(.width(width)) rd_st5_1345  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1345]), .rdlo_in(a5_wr[1377]),  .coef_in(coef[32]), .rdup_out(a6_wr[1345]), .rdlo_out(a6_wr[1377]));
			radix2 #(.width(width)) rd_st5_1346  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1346]), .rdlo_in(a5_wr[1378]),  .coef_in(coef[64]), .rdup_out(a6_wr[1346]), .rdlo_out(a6_wr[1378]));
			radix2 #(.width(width)) rd_st5_1347  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1347]), .rdlo_in(a5_wr[1379]),  .coef_in(coef[96]), .rdup_out(a6_wr[1347]), .rdlo_out(a6_wr[1379]));
			radix2 #(.width(width)) rd_st5_1348  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1348]), .rdlo_in(a5_wr[1380]),  .coef_in(coef[128]), .rdup_out(a6_wr[1348]), .rdlo_out(a6_wr[1380]));
			radix2 #(.width(width)) rd_st5_1349  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1349]), .rdlo_in(a5_wr[1381]),  .coef_in(coef[160]), .rdup_out(a6_wr[1349]), .rdlo_out(a6_wr[1381]));
			radix2 #(.width(width)) rd_st5_1350  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1350]), .rdlo_in(a5_wr[1382]),  .coef_in(coef[192]), .rdup_out(a6_wr[1350]), .rdlo_out(a6_wr[1382]));
			radix2 #(.width(width)) rd_st5_1351  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1351]), .rdlo_in(a5_wr[1383]),  .coef_in(coef[224]), .rdup_out(a6_wr[1351]), .rdlo_out(a6_wr[1383]));
			radix2 #(.width(width)) rd_st5_1352  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1352]), .rdlo_in(a5_wr[1384]),  .coef_in(coef[256]), .rdup_out(a6_wr[1352]), .rdlo_out(a6_wr[1384]));
			radix2 #(.width(width)) rd_st5_1353  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1353]), .rdlo_in(a5_wr[1385]),  .coef_in(coef[288]), .rdup_out(a6_wr[1353]), .rdlo_out(a6_wr[1385]));
			radix2 #(.width(width)) rd_st5_1354  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1354]), .rdlo_in(a5_wr[1386]),  .coef_in(coef[320]), .rdup_out(a6_wr[1354]), .rdlo_out(a6_wr[1386]));
			radix2 #(.width(width)) rd_st5_1355  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1355]), .rdlo_in(a5_wr[1387]),  .coef_in(coef[352]), .rdup_out(a6_wr[1355]), .rdlo_out(a6_wr[1387]));
			radix2 #(.width(width)) rd_st5_1356  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1356]), .rdlo_in(a5_wr[1388]),  .coef_in(coef[384]), .rdup_out(a6_wr[1356]), .rdlo_out(a6_wr[1388]));
			radix2 #(.width(width)) rd_st5_1357  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1357]), .rdlo_in(a5_wr[1389]),  .coef_in(coef[416]), .rdup_out(a6_wr[1357]), .rdlo_out(a6_wr[1389]));
			radix2 #(.width(width)) rd_st5_1358  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1358]), .rdlo_in(a5_wr[1390]),  .coef_in(coef[448]), .rdup_out(a6_wr[1358]), .rdlo_out(a6_wr[1390]));
			radix2 #(.width(width)) rd_st5_1359  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1359]), .rdlo_in(a5_wr[1391]),  .coef_in(coef[480]), .rdup_out(a6_wr[1359]), .rdlo_out(a6_wr[1391]));
			radix2 #(.width(width)) rd_st5_1360  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1360]), .rdlo_in(a5_wr[1392]),  .coef_in(coef[512]), .rdup_out(a6_wr[1360]), .rdlo_out(a6_wr[1392]));
			radix2 #(.width(width)) rd_st5_1361  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1361]), .rdlo_in(a5_wr[1393]),  .coef_in(coef[544]), .rdup_out(a6_wr[1361]), .rdlo_out(a6_wr[1393]));
			radix2 #(.width(width)) rd_st5_1362  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1362]), .rdlo_in(a5_wr[1394]),  .coef_in(coef[576]), .rdup_out(a6_wr[1362]), .rdlo_out(a6_wr[1394]));
			radix2 #(.width(width)) rd_st5_1363  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1363]), .rdlo_in(a5_wr[1395]),  .coef_in(coef[608]), .rdup_out(a6_wr[1363]), .rdlo_out(a6_wr[1395]));
			radix2 #(.width(width)) rd_st5_1364  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1364]), .rdlo_in(a5_wr[1396]),  .coef_in(coef[640]), .rdup_out(a6_wr[1364]), .rdlo_out(a6_wr[1396]));
			radix2 #(.width(width)) rd_st5_1365  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1365]), .rdlo_in(a5_wr[1397]),  .coef_in(coef[672]), .rdup_out(a6_wr[1365]), .rdlo_out(a6_wr[1397]));
			radix2 #(.width(width)) rd_st5_1366  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1366]), .rdlo_in(a5_wr[1398]),  .coef_in(coef[704]), .rdup_out(a6_wr[1366]), .rdlo_out(a6_wr[1398]));
			radix2 #(.width(width)) rd_st5_1367  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1367]), .rdlo_in(a5_wr[1399]),  .coef_in(coef[736]), .rdup_out(a6_wr[1367]), .rdlo_out(a6_wr[1399]));
			radix2 #(.width(width)) rd_st5_1368  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1368]), .rdlo_in(a5_wr[1400]),  .coef_in(coef[768]), .rdup_out(a6_wr[1368]), .rdlo_out(a6_wr[1400]));
			radix2 #(.width(width)) rd_st5_1369  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1369]), .rdlo_in(a5_wr[1401]),  .coef_in(coef[800]), .rdup_out(a6_wr[1369]), .rdlo_out(a6_wr[1401]));
			radix2 #(.width(width)) rd_st5_1370  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1370]), .rdlo_in(a5_wr[1402]),  .coef_in(coef[832]), .rdup_out(a6_wr[1370]), .rdlo_out(a6_wr[1402]));
			radix2 #(.width(width)) rd_st5_1371  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1371]), .rdlo_in(a5_wr[1403]),  .coef_in(coef[864]), .rdup_out(a6_wr[1371]), .rdlo_out(a6_wr[1403]));
			radix2 #(.width(width)) rd_st5_1372  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1372]), .rdlo_in(a5_wr[1404]),  .coef_in(coef[896]), .rdup_out(a6_wr[1372]), .rdlo_out(a6_wr[1404]));
			radix2 #(.width(width)) rd_st5_1373  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1373]), .rdlo_in(a5_wr[1405]),  .coef_in(coef[928]), .rdup_out(a6_wr[1373]), .rdlo_out(a6_wr[1405]));
			radix2 #(.width(width)) rd_st5_1374  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1374]), .rdlo_in(a5_wr[1406]),  .coef_in(coef[960]), .rdup_out(a6_wr[1374]), .rdlo_out(a6_wr[1406]));
			radix2 #(.width(width)) rd_st5_1375  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1375]), .rdlo_in(a5_wr[1407]),  .coef_in(coef[992]), .rdup_out(a6_wr[1375]), .rdlo_out(a6_wr[1407]));
			radix2 #(.width(width)) rd_st5_1408  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1408]), .rdlo_in(a5_wr[1440]),  .coef_in(coef[0]), .rdup_out(a6_wr[1408]), .rdlo_out(a6_wr[1440]));
			radix2 #(.width(width)) rd_st5_1409  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1409]), .rdlo_in(a5_wr[1441]),  .coef_in(coef[32]), .rdup_out(a6_wr[1409]), .rdlo_out(a6_wr[1441]));
			radix2 #(.width(width)) rd_st5_1410  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1410]), .rdlo_in(a5_wr[1442]),  .coef_in(coef[64]), .rdup_out(a6_wr[1410]), .rdlo_out(a6_wr[1442]));
			radix2 #(.width(width)) rd_st5_1411  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1411]), .rdlo_in(a5_wr[1443]),  .coef_in(coef[96]), .rdup_out(a6_wr[1411]), .rdlo_out(a6_wr[1443]));
			radix2 #(.width(width)) rd_st5_1412  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1412]), .rdlo_in(a5_wr[1444]),  .coef_in(coef[128]), .rdup_out(a6_wr[1412]), .rdlo_out(a6_wr[1444]));
			radix2 #(.width(width)) rd_st5_1413  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1413]), .rdlo_in(a5_wr[1445]),  .coef_in(coef[160]), .rdup_out(a6_wr[1413]), .rdlo_out(a6_wr[1445]));
			radix2 #(.width(width)) rd_st5_1414  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1414]), .rdlo_in(a5_wr[1446]),  .coef_in(coef[192]), .rdup_out(a6_wr[1414]), .rdlo_out(a6_wr[1446]));
			radix2 #(.width(width)) rd_st5_1415  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1415]), .rdlo_in(a5_wr[1447]),  .coef_in(coef[224]), .rdup_out(a6_wr[1415]), .rdlo_out(a6_wr[1447]));
			radix2 #(.width(width)) rd_st5_1416  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1416]), .rdlo_in(a5_wr[1448]),  .coef_in(coef[256]), .rdup_out(a6_wr[1416]), .rdlo_out(a6_wr[1448]));
			radix2 #(.width(width)) rd_st5_1417  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1417]), .rdlo_in(a5_wr[1449]),  .coef_in(coef[288]), .rdup_out(a6_wr[1417]), .rdlo_out(a6_wr[1449]));
			radix2 #(.width(width)) rd_st5_1418  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1418]), .rdlo_in(a5_wr[1450]),  .coef_in(coef[320]), .rdup_out(a6_wr[1418]), .rdlo_out(a6_wr[1450]));
			radix2 #(.width(width)) rd_st5_1419  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1419]), .rdlo_in(a5_wr[1451]),  .coef_in(coef[352]), .rdup_out(a6_wr[1419]), .rdlo_out(a6_wr[1451]));
			radix2 #(.width(width)) rd_st5_1420  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1420]), .rdlo_in(a5_wr[1452]),  .coef_in(coef[384]), .rdup_out(a6_wr[1420]), .rdlo_out(a6_wr[1452]));
			radix2 #(.width(width)) rd_st5_1421  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1421]), .rdlo_in(a5_wr[1453]),  .coef_in(coef[416]), .rdup_out(a6_wr[1421]), .rdlo_out(a6_wr[1453]));
			radix2 #(.width(width)) rd_st5_1422  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1422]), .rdlo_in(a5_wr[1454]),  .coef_in(coef[448]), .rdup_out(a6_wr[1422]), .rdlo_out(a6_wr[1454]));
			radix2 #(.width(width)) rd_st5_1423  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1423]), .rdlo_in(a5_wr[1455]),  .coef_in(coef[480]), .rdup_out(a6_wr[1423]), .rdlo_out(a6_wr[1455]));
			radix2 #(.width(width)) rd_st5_1424  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1424]), .rdlo_in(a5_wr[1456]),  .coef_in(coef[512]), .rdup_out(a6_wr[1424]), .rdlo_out(a6_wr[1456]));
			radix2 #(.width(width)) rd_st5_1425  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1425]), .rdlo_in(a5_wr[1457]),  .coef_in(coef[544]), .rdup_out(a6_wr[1425]), .rdlo_out(a6_wr[1457]));
			radix2 #(.width(width)) rd_st5_1426  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1426]), .rdlo_in(a5_wr[1458]),  .coef_in(coef[576]), .rdup_out(a6_wr[1426]), .rdlo_out(a6_wr[1458]));
			radix2 #(.width(width)) rd_st5_1427  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1427]), .rdlo_in(a5_wr[1459]),  .coef_in(coef[608]), .rdup_out(a6_wr[1427]), .rdlo_out(a6_wr[1459]));
			radix2 #(.width(width)) rd_st5_1428  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1428]), .rdlo_in(a5_wr[1460]),  .coef_in(coef[640]), .rdup_out(a6_wr[1428]), .rdlo_out(a6_wr[1460]));
			radix2 #(.width(width)) rd_st5_1429  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1429]), .rdlo_in(a5_wr[1461]),  .coef_in(coef[672]), .rdup_out(a6_wr[1429]), .rdlo_out(a6_wr[1461]));
			radix2 #(.width(width)) rd_st5_1430  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1430]), .rdlo_in(a5_wr[1462]),  .coef_in(coef[704]), .rdup_out(a6_wr[1430]), .rdlo_out(a6_wr[1462]));
			radix2 #(.width(width)) rd_st5_1431  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1431]), .rdlo_in(a5_wr[1463]),  .coef_in(coef[736]), .rdup_out(a6_wr[1431]), .rdlo_out(a6_wr[1463]));
			radix2 #(.width(width)) rd_st5_1432  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1432]), .rdlo_in(a5_wr[1464]),  .coef_in(coef[768]), .rdup_out(a6_wr[1432]), .rdlo_out(a6_wr[1464]));
			radix2 #(.width(width)) rd_st5_1433  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1433]), .rdlo_in(a5_wr[1465]),  .coef_in(coef[800]), .rdup_out(a6_wr[1433]), .rdlo_out(a6_wr[1465]));
			radix2 #(.width(width)) rd_st5_1434  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1434]), .rdlo_in(a5_wr[1466]),  .coef_in(coef[832]), .rdup_out(a6_wr[1434]), .rdlo_out(a6_wr[1466]));
			radix2 #(.width(width)) rd_st5_1435  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1435]), .rdlo_in(a5_wr[1467]),  .coef_in(coef[864]), .rdup_out(a6_wr[1435]), .rdlo_out(a6_wr[1467]));
			radix2 #(.width(width)) rd_st5_1436  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1436]), .rdlo_in(a5_wr[1468]),  .coef_in(coef[896]), .rdup_out(a6_wr[1436]), .rdlo_out(a6_wr[1468]));
			radix2 #(.width(width)) rd_st5_1437  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1437]), .rdlo_in(a5_wr[1469]),  .coef_in(coef[928]), .rdup_out(a6_wr[1437]), .rdlo_out(a6_wr[1469]));
			radix2 #(.width(width)) rd_st5_1438  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1438]), .rdlo_in(a5_wr[1470]),  .coef_in(coef[960]), .rdup_out(a6_wr[1438]), .rdlo_out(a6_wr[1470]));
			radix2 #(.width(width)) rd_st5_1439  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1439]), .rdlo_in(a5_wr[1471]),  .coef_in(coef[992]), .rdup_out(a6_wr[1439]), .rdlo_out(a6_wr[1471]));
			radix2 #(.width(width)) rd_st5_1472  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1472]), .rdlo_in(a5_wr[1504]),  .coef_in(coef[0]), .rdup_out(a6_wr[1472]), .rdlo_out(a6_wr[1504]));
			radix2 #(.width(width)) rd_st5_1473  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1473]), .rdlo_in(a5_wr[1505]),  .coef_in(coef[32]), .rdup_out(a6_wr[1473]), .rdlo_out(a6_wr[1505]));
			radix2 #(.width(width)) rd_st5_1474  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1474]), .rdlo_in(a5_wr[1506]),  .coef_in(coef[64]), .rdup_out(a6_wr[1474]), .rdlo_out(a6_wr[1506]));
			radix2 #(.width(width)) rd_st5_1475  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1475]), .rdlo_in(a5_wr[1507]),  .coef_in(coef[96]), .rdup_out(a6_wr[1475]), .rdlo_out(a6_wr[1507]));
			radix2 #(.width(width)) rd_st5_1476  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1476]), .rdlo_in(a5_wr[1508]),  .coef_in(coef[128]), .rdup_out(a6_wr[1476]), .rdlo_out(a6_wr[1508]));
			radix2 #(.width(width)) rd_st5_1477  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1477]), .rdlo_in(a5_wr[1509]),  .coef_in(coef[160]), .rdup_out(a6_wr[1477]), .rdlo_out(a6_wr[1509]));
			radix2 #(.width(width)) rd_st5_1478  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1478]), .rdlo_in(a5_wr[1510]),  .coef_in(coef[192]), .rdup_out(a6_wr[1478]), .rdlo_out(a6_wr[1510]));
			radix2 #(.width(width)) rd_st5_1479  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1479]), .rdlo_in(a5_wr[1511]),  .coef_in(coef[224]), .rdup_out(a6_wr[1479]), .rdlo_out(a6_wr[1511]));
			radix2 #(.width(width)) rd_st5_1480  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1480]), .rdlo_in(a5_wr[1512]),  .coef_in(coef[256]), .rdup_out(a6_wr[1480]), .rdlo_out(a6_wr[1512]));
			radix2 #(.width(width)) rd_st5_1481  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1481]), .rdlo_in(a5_wr[1513]),  .coef_in(coef[288]), .rdup_out(a6_wr[1481]), .rdlo_out(a6_wr[1513]));
			radix2 #(.width(width)) rd_st5_1482  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1482]), .rdlo_in(a5_wr[1514]),  .coef_in(coef[320]), .rdup_out(a6_wr[1482]), .rdlo_out(a6_wr[1514]));
			radix2 #(.width(width)) rd_st5_1483  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1483]), .rdlo_in(a5_wr[1515]),  .coef_in(coef[352]), .rdup_out(a6_wr[1483]), .rdlo_out(a6_wr[1515]));
			radix2 #(.width(width)) rd_st5_1484  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1484]), .rdlo_in(a5_wr[1516]),  .coef_in(coef[384]), .rdup_out(a6_wr[1484]), .rdlo_out(a6_wr[1516]));
			radix2 #(.width(width)) rd_st5_1485  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1485]), .rdlo_in(a5_wr[1517]),  .coef_in(coef[416]), .rdup_out(a6_wr[1485]), .rdlo_out(a6_wr[1517]));
			radix2 #(.width(width)) rd_st5_1486  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1486]), .rdlo_in(a5_wr[1518]),  .coef_in(coef[448]), .rdup_out(a6_wr[1486]), .rdlo_out(a6_wr[1518]));
			radix2 #(.width(width)) rd_st5_1487  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1487]), .rdlo_in(a5_wr[1519]),  .coef_in(coef[480]), .rdup_out(a6_wr[1487]), .rdlo_out(a6_wr[1519]));
			radix2 #(.width(width)) rd_st5_1488  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1488]), .rdlo_in(a5_wr[1520]),  .coef_in(coef[512]), .rdup_out(a6_wr[1488]), .rdlo_out(a6_wr[1520]));
			radix2 #(.width(width)) rd_st5_1489  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1489]), .rdlo_in(a5_wr[1521]),  .coef_in(coef[544]), .rdup_out(a6_wr[1489]), .rdlo_out(a6_wr[1521]));
			radix2 #(.width(width)) rd_st5_1490  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1490]), .rdlo_in(a5_wr[1522]),  .coef_in(coef[576]), .rdup_out(a6_wr[1490]), .rdlo_out(a6_wr[1522]));
			radix2 #(.width(width)) rd_st5_1491  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1491]), .rdlo_in(a5_wr[1523]),  .coef_in(coef[608]), .rdup_out(a6_wr[1491]), .rdlo_out(a6_wr[1523]));
			radix2 #(.width(width)) rd_st5_1492  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1492]), .rdlo_in(a5_wr[1524]),  .coef_in(coef[640]), .rdup_out(a6_wr[1492]), .rdlo_out(a6_wr[1524]));
			radix2 #(.width(width)) rd_st5_1493  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1493]), .rdlo_in(a5_wr[1525]),  .coef_in(coef[672]), .rdup_out(a6_wr[1493]), .rdlo_out(a6_wr[1525]));
			radix2 #(.width(width)) rd_st5_1494  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1494]), .rdlo_in(a5_wr[1526]),  .coef_in(coef[704]), .rdup_out(a6_wr[1494]), .rdlo_out(a6_wr[1526]));
			radix2 #(.width(width)) rd_st5_1495  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1495]), .rdlo_in(a5_wr[1527]),  .coef_in(coef[736]), .rdup_out(a6_wr[1495]), .rdlo_out(a6_wr[1527]));
			radix2 #(.width(width)) rd_st5_1496  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1496]), .rdlo_in(a5_wr[1528]),  .coef_in(coef[768]), .rdup_out(a6_wr[1496]), .rdlo_out(a6_wr[1528]));
			radix2 #(.width(width)) rd_st5_1497  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1497]), .rdlo_in(a5_wr[1529]),  .coef_in(coef[800]), .rdup_out(a6_wr[1497]), .rdlo_out(a6_wr[1529]));
			radix2 #(.width(width)) rd_st5_1498  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1498]), .rdlo_in(a5_wr[1530]),  .coef_in(coef[832]), .rdup_out(a6_wr[1498]), .rdlo_out(a6_wr[1530]));
			radix2 #(.width(width)) rd_st5_1499  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1499]), .rdlo_in(a5_wr[1531]),  .coef_in(coef[864]), .rdup_out(a6_wr[1499]), .rdlo_out(a6_wr[1531]));
			radix2 #(.width(width)) rd_st5_1500  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1500]), .rdlo_in(a5_wr[1532]),  .coef_in(coef[896]), .rdup_out(a6_wr[1500]), .rdlo_out(a6_wr[1532]));
			radix2 #(.width(width)) rd_st5_1501  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1501]), .rdlo_in(a5_wr[1533]),  .coef_in(coef[928]), .rdup_out(a6_wr[1501]), .rdlo_out(a6_wr[1533]));
			radix2 #(.width(width)) rd_st5_1502  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1502]), .rdlo_in(a5_wr[1534]),  .coef_in(coef[960]), .rdup_out(a6_wr[1502]), .rdlo_out(a6_wr[1534]));
			radix2 #(.width(width)) rd_st5_1503  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1503]), .rdlo_in(a5_wr[1535]),  .coef_in(coef[992]), .rdup_out(a6_wr[1503]), .rdlo_out(a6_wr[1535]));
			radix2 #(.width(width)) rd_st5_1536  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1536]), .rdlo_in(a5_wr[1568]),  .coef_in(coef[0]), .rdup_out(a6_wr[1536]), .rdlo_out(a6_wr[1568]));
			radix2 #(.width(width)) rd_st5_1537  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1537]), .rdlo_in(a5_wr[1569]),  .coef_in(coef[32]), .rdup_out(a6_wr[1537]), .rdlo_out(a6_wr[1569]));
			radix2 #(.width(width)) rd_st5_1538  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1538]), .rdlo_in(a5_wr[1570]),  .coef_in(coef[64]), .rdup_out(a6_wr[1538]), .rdlo_out(a6_wr[1570]));
			radix2 #(.width(width)) rd_st5_1539  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1539]), .rdlo_in(a5_wr[1571]),  .coef_in(coef[96]), .rdup_out(a6_wr[1539]), .rdlo_out(a6_wr[1571]));
			radix2 #(.width(width)) rd_st5_1540  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1540]), .rdlo_in(a5_wr[1572]),  .coef_in(coef[128]), .rdup_out(a6_wr[1540]), .rdlo_out(a6_wr[1572]));
			radix2 #(.width(width)) rd_st5_1541  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1541]), .rdlo_in(a5_wr[1573]),  .coef_in(coef[160]), .rdup_out(a6_wr[1541]), .rdlo_out(a6_wr[1573]));
			radix2 #(.width(width)) rd_st5_1542  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1542]), .rdlo_in(a5_wr[1574]),  .coef_in(coef[192]), .rdup_out(a6_wr[1542]), .rdlo_out(a6_wr[1574]));
			radix2 #(.width(width)) rd_st5_1543  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1543]), .rdlo_in(a5_wr[1575]),  .coef_in(coef[224]), .rdup_out(a6_wr[1543]), .rdlo_out(a6_wr[1575]));
			radix2 #(.width(width)) rd_st5_1544  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1544]), .rdlo_in(a5_wr[1576]),  .coef_in(coef[256]), .rdup_out(a6_wr[1544]), .rdlo_out(a6_wr[1576]));
			radix2 #(.width(width)) rd_st5_1545  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1545]), .rdlo_in(a5_wr[1577]),  .coef_in(coef[288]), .rdup_out(a6_wr[1545]), .rdlo_out(a6_wr[1577]));
			radix2 #(.width(width)) rd_st5_1546  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1546]), .rdlo_in(a5_wr[1578]),  .coef_in(coef[320]), .rdup_out(a6_wr[1546]), .rdlo_out(a6_wr[1578]));
			radix2 #(.width(width)) rd_st5_1547  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1547]), .rdlo_in(a5_wr[1579]),  .coef_in(coef[352]), .rdup_out(a6_wr[1547]), .rdlo_out(a6_wr[1579]));
			radix2 #(.width(width)) rd_st5_1548  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1548]), .rdlo_in(a5_wr[1580]),  .coef_in(coef[384]), .rdup_out(a6_wr[1548]), .rdlo_out(a6_wr[1580]));
			radix2 #(.width(width)) rd_st5_1549  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1549]), .rdlo_in(a5_wr[1581]),  .coef_in(coef[416]), .rdup_out(a6_wr[1549]), .rdlo_out(a6_wr[1581]));
			radix2 #(.width(width)) rd_st5_1550  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1550]), .rdlo_in(a5_wr[1582]),  .coef_in(coef[448]), .rdup_out(a6_wr[1550]), .rdlo_out(a6_wr[1582]));
			radix2 #(.width(width)) rd_st5_1551  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1551]), .rdlo_in(a5_wr[1583]),  .coef_in(coef[480]), .rdup_out(a6_wr[1551]), .rdlo_out(a6_wr[1583]));
			radix2 #(.width(width)) rd_st5_1552  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1552]), .rdlo_in(a5_wr[1584]),  .coef_in(coef[512]), .rdup_out(a6_wr[1552]), .rdlo_out(a6_wr[1584]));
			radix2 #(.width(width)) rd_st5_1553  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1553]), .rdlo_in(a5_wr[1585]),  .coef_in(coef[544]), .rdup_out(a6_wr[1553]), .rdlo_out(a6_wr[1585]));
			radix2 #(.width(width)) rd_st5_1554  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1554]), .rdlo_in(a5_wr[1586]),  .coef_in(coef[576]), .rdup_out(a6_wr[1554]), .rdlo_out(a6_wr[1586]));
			radix2 #(.width(width)) rd_st5_1555  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1555]), .rdlo_in(a5_wr[1587]),  .coef_in(coef[608]), .rdup_out(a6_wr[1555]), .rdlo_out(a6_wr[1587]));
			radix2 #(.width(width)) rd_st5_1556  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1556]), .rdlo_in(a5_wr[1588]),  .coef_in(coef[640]), .rdup_out(a6_wr[1556]), .rdlo_out(a6_wr[1588]));
			radix2 #(.width(width)) rd_st5_1557  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1557]), .rdlo_in(a5_wr[1589]),  .coef_in(coef[672]), .rdup_out(a6_wr[1557]), .rdlo_out(a6_wr[1589]));
			radix2 #(.width(width)) rd_st5_1558  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1558]), .rdlo_in(a5_wr[1590]),  .coef_in(coef[704]), .rdup_out(a6_wr[1558]), .rdlo_out(a6_wr[1590]));
			radix2 #(.width(width)) rd_st5_1559  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1559]), .rdlo_in(a5_wr[1591]),  .coef_in(coef[736]), .rdup_out(a6_wr[1559]), .rdlo_out(a6_wr[1591]));
			radix2 #(.width(width)) rd_st5_1560  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1560]), .rdlo_in(a5_wr[1592]),  .coef_in(coef[768]), .rdup_out(a6_wr[1560]), .rdlo_out(a6_wr[1592]));
			radix2 #(.width(width)) rd_st5_1561  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1561]), .rdlo_in(a5_wr[1593]),  .coef_in(coef[800]), .rdup_out(a6_wr[1561]), .rdlo_out(a6_wr[1593]));
			radix2 #(.width(width)) rd_st5_1562  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1562]), .rdlo_in(a5_wr[1594]),  .coef_in(coef[832]), .rdup_out(a6_wr[1562]), .rdlo_out(a6_wr[1594]));
			radix2 #(.width(width)) rd_st5_1563  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1563]), .rdlo_in(a5_wr[1595]),  .coef_in(coef[864]), .rdup_out(a6_wr[1563]), .rdlo_out(a6_wr[1595]));
			radix2 #(.width(width)) rd_st5_1564  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1564]), .rdlo_in(a5_wr[1596]),  .coef_in(coef[896]), .rdup_out(a6_wr[1564]), .rdlo_out(a6_wr[1596]));
			radix2 #(.width(width)) rd_st5_1565  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1565]), .rdlo_in(a5_wr[1597]),  .coef_in(coef[928]), .rdup_out(a6_wr[1565]), .rdlo_out(a6_wr[1597]));
			radix2 #(.width(width)) rd_st5_1566  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1566]), .rdlo_in(a5_wr[1598]),  .coef_in(coef[960]), .rdup_out(a6_wr[1566]), .rdlo_out(a6_wr[1598]));
			radix2 #(.width(width)) rd_st5_1567  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1567]), .rdlo_in(a5_wr[1599]),  .coef_in(coef[992]), .rdup_out(a6_wr[1567]), .rdlo_out(a6_wr[1599]));
			radix2 #(.width(width)) rd_st5_1600  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1600]), .rdlo_in(a5_wr[1632]),  .coef_in(coef[0]), .rdup_out(a6_wr[1600]), .rdlo_out(a6_wr[1632]));
			radix2 #(.width(width)) rd_st5_1601  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1601]), .rdlo_in(a5_wr[1633]),  .coef_in(coef[32]), .rdup_out(a6_wr[1601]), .rdlo_out(a6_wr[1633]));
			radix2 #(.width(width)) rd_st5_1602  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1602]), .rdlo_in(a5_wr[1634]),  .coef_in(coef[64]), .rdup_out(a6_wr[1602]), .rdlo_out(a6_wr[1634]));
			radix2 #(.width(width)) rd_st5_1603  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1603]), .rdlo_in(a5_wr[1635]),  .coef_in(coef[96]), .rdup_out(a6_wr[1603]), .rdlo_out(a6_wr[1635]));
			radix2 #(.width(width)) rd_st5_1604  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1604]), .rdlo_in(a5_wr[1636]),  .coef_in(coef[128]), .rdup_out(a6_wr[1604]), .rdlo_out(a6_wr[1636]));
			radix2 #(.width(width)) rd_st5_1605  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1605]), .rdlo_in(a5_wr[1637]),  .coef_in(coef[160]), .rdup_out(a6_wr[1605]), .rdlo_out(a6_wr[1637]));
			radix2 #(.width(width)) rd_st5_1606  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1606]), .rdlo_in(a5_wr[1638]),  .coef_in(coef[192]), .rdup_out(a6_wr[1606]), .rdlo_out(a6_wr[1638]));
			radix2 #(.width(width)) rd_st5_1607  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1607]), .rdlo_in(a5_wr[1639]),  .coef_in(coef[224]), .rdup_out(a6_wr[1607]), .rdlo_out(a6_wr[1639]));
			radix2 #(.width(width)) rd_st5_1608  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1608]), .rdlo_in(a5_wr[1640]),  .coef_in(coef[256]), .rdup_out(a6_wr[1608]), .rdlo_out(a6_wr[1640]));
			radix2 #(.width(width)) rd_st5_1609  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1609]), .rdlo_in(a5_wr[1641]),  .coef_in(coef[288]), .rdup_out(a6_wr[1609]), .rdlo_out(a6_wr[1641]));
			radix2 #(.width(width)) rd_st5_1610  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1610]), .rdlo_in(a5_wr[1642]),  .coef_in(coef[320]), .rdup_out(a6_wr[1610]), .rdlo_out(a6_wr[1642]));
			radix2 #(.width(width)) rd_st5_1611  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1611]), .rdlo_in(a5_wr[1643]),  .coef_in(coef[352]), .rdup_out(a6_wr[1611]), .rdlo_out(a6_wr[1643]));
			radix2 #(.width(width)) rd_st5_1612  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1612]), .rdlo_in(a5_wr[1644]),  .coef_in(coef[384]), .rdup_out(a6_wr[1612]), .rdlo_out(a6_wr[1644]));
			radix2 #(.width(width)) rd_st5_1613  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1613]), .rdlo_in(a5_wr[1645]),  .coef_in(coef[416]), .rdup_out(a6_wr[1613]), .rdlo_out(a6_wr[1645]));
			radix2 #(.width(width)) rd_st5_1614  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1614]), .rdlo_in(a5_wr[1646]),  .coef_in(coef[448]), .rdup_out(a6_wr[1614]), .rdlo_out(a6_wr[1646]));
			radix2 #(.width(width)) rd_st5_1615  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1615]), .rdlo_in(a5_wr[1647]),  .coef_in(coef[480]), .rdup_out(a6_wr[1615]), .rdlo_out(a6_wr[1647]));
			radix2 #(.width(width)) rd_st5_1616  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1616]), .rdlo_in(a5_wr[1648]),  .coef_in(coef[512]), .rdup_out(a6_wr[1616]), .rdlo_out(a6_wr[1648]));
			radix2 #(.width(width)) rd_st5_1617  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1617]), .rdlo_in(a5_wr[1649]),  .coef_in(coef[544]), .rdup_out(a6_wr[1617]), .rdlo_out(a6_wr[1649]));
			radix2 #(.width(width)) rd_st5_1618  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1618]), .rdlo_in(a5_wr[1650]),  .coef_in(coef[576]), .rdup_out(a6_wr[1618]), .rdlo_out(a6_wr[1650]));
			radix2 #(.width(width)) rd_st5_1619  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1619]), .rdlo_in(a5_wr[1651]),  .coef_in(coef[608]), .rdup_out(a6_wr[1619]), .rdlo_out(a6_wr[1651]));
			radix2 #(.width(width)) rd_st5_1620  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1620]), .rdlo_in(a5_wr[1652]),  .coef_in(coef[640]), .rdup_out(a6_wr[1620]), .rdlo_out(a6_wr[1652]));
			radix2 #(.width(width)) rd_st5_1621  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1621]), .rdlo_in(a5_wr[1653]),  .coef_in(coef[672]), .rdup_out(a6_wr[1621]), .rdlo_out(a6_wr[1653]));
			radix2 #(.width(width)) rd_st5_1622  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1622]), .rdlo_in(a5_wr[1654]),  .coef_in(coef[704]), .rdup_out(a6_wr[1622]), .rdlo_out(a6_wr[1654]));
			radix2 #(.width(width)) rd_st5_1623  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1623]), .rdlo_in(a5_wr[1655]),  .coef_in(coef[736]), .rdup_out(a6_wr[1623]), .rdlo_out(a6_wr[1655]));
			radix2 #(.width(width)) rd_st5_1624  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1624]), .rdlo_in(a5_wr[1656]),  .coef_in(coef[768]), .rdup_out(a6_wr[1624]), .rdlo_out(a6_wr[1656]));
			radix2 #(.width(width)) rd_st5_1625  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1625]), .rdlo_in(a5_wr[1657]),  .coef_in(coef[800]), .rdup_out(a6_wr[1625]), .rdlo_out(a6_wr[1657]));
			radix2 #(.width(width)) rd_st5_1626  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1626]), .rdlo_in(a5_wr[1658]),  .coef_in(coef[832]), .rdup_out(a6_wr[1626]), .rdlo_out(a6_wr[1658]));
			radix2 #(.width(width)) rd_st5_1627  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1627]), .rdlo_in(a5_wr[1659]),  .coef_in(coef[864]), .rdup_out(a6_wr[1627]), .rdlo_out(a6_wr[1659]));
			radix2 #(.width(width)) rd_st5_1628  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1628]), .rdlo_in(a5_wr[1660]),  .coef_in(coef[896]), .rdup_out(a6_wr[1628]), .rdlo_out(a6_wr[1660]));
			radix2 #(.width(width)) rd_st5_1629  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1629]), .rdlo_in(a5_wr[1661]),  .coef_in(coef[928]), .rdup_out(a6_wr[1629]), .rdlo_out(a6_wr[1661]));
			radix2 #(.width(width)) rd_st5_1630  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1630]), .rdlo_in(a5_wr[1662]),  .coef_in(coef[960]), .rdup_out(a6_wr[1630]), .rdlo_out(a6_wr[1662]));
			radix2 #(.width(width)) rd_st5_1631  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1631]), .rdlo_in(a5_wr[1663]),  .coef_in(coef[992]), .rdup_out(a6_wr[1631]), .rdlo_out(a6_wr[1663]));
			radix2 #(.width(width)) rd_st5_1664  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1664]), .rdlo_in(a5_wr[1696]),  .coef_in(coef[0]), .rdup_out(a6_wr[1664]), .rdlo_out(a6_wr[1696]));
			radix2 #(.width(width)) rd_st5_1665  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1665]), .rdlo_in(a5_wr[1697]),  .coef_in(coef[32]), .rdup_out(a6_wr[1665]), .rdlo_out(a6_wr[1697]));
			radix2 #(.width(width)) rd_st5_1666  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1666]), .rdlo_in(a5_wr[1698]),  .coef_in(coef[64]), .rdup_out(a6_wr[1666]), .rdlo_out(a6_wr[1698]));
			radix2 #(.width(width)) rd_st5_1667  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1667]), .rdlo_in(a5_wr[1699]),  .coef_in(coef[96]), .rdup_out(a6_wr[1667]), .rdlo_out(a6_wr[1699]));
			radix2 #(.width(width)) rd_st5_1668  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1668]), .rdlo_in(a5_wr[1700]),  .coef_in(coef[128]), .rdup_out(a6_wr[1668]), .rdlo_out(a6_wr[1700]));
			radix2 #(.width(width)) rd_st5_1669  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1669]), .rdlo_in(a5_wr[1701]),  .coef_in(coef[160]), .rdup_out(a6_wr[1669]), .rdlo_out(a6_wr[1701]));
			radix2 #(.width(width)) rd_st5_1670  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1670]), .rdlo_in(a5_wr[1702]),  .coef_in(coef[192]), .rdup_out(a6_wr[1670]), .rdlo_out(a6_wr[1702]));
			radix2 #(.width(width)) rd_st5_1671  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1671]), .rdlo_in(a5_wr[1703]),  .coef_in(coef[224]), .rdup_out(a6_wr[1671]), .rdlo_out(a6_wr[1703]));
			radix2 #(.width(width)) rd_st5_1672  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1672]), .rdlo_in(a5_wr[1704]),  .coef_in(coef[256]), .rdup_out(a6_wr[1672]), .rdlo_out(a6_wr[1704]));
			radix2 #(.width(width)) rd_st5_1673  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1673]), .rdlo_in(a5_wr[1705]),  .coef_in(coef[288]), .rdup_out(a6_wr[1673]), .rdlo_out(a6_wr[1705]));
			radix2 #(.width(width)) rd_st5_1674  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1674]), .rdlo_in(a5_wr[1706]),  .coef_in(coef[320]), .rdup_out(a6_wr[1674]), .rdlo_out(a6_wr[1706]));
			radix2 #(.width(width)) rd_st5_1675  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1675]), .rdlo_in(a5_wr[1707]),  .coef_in(coef[352]), .rdup_out(a6_wr[1675]), .rdlo_out(a6_wr[1707]));
			radix2 #(.width(width)) rd_st5_1676  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1676]), .rdlo_in(a5_wr[1708]),  .coef_in(coef[384]), .rdup_out(a6_wr[1676]), .rdlo_out(a6_wr[1708]));
			radix2 #(.width(width)) rd_st5_1677  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1677]), .rdlo_in(a5_wr[1709]),  .coef_in(coef[416]), .rdup_out(a6_wr[1677]), .rdlo_out(a6_wr[1709]));
			radix2 #(.width(width)) rd_st5_1678  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1678]), .rdlo_in(a5_wr[1710]),  .coef_in(coef[448]), .rdup_out(a6_wr[1678]), .rdlo_out(a6_wr[1710]));
			radix2 #(.width(width)) rd_st5_1679  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1679]), .rdlo_in(a5_wr[1711]),  .coef_in(coef[480]), .rdup_out(a6_wr[1679]), .rdlo_out(a6_wr[1711]));
			radix2 #(.width(width)) rd_st5_1680  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1680]), .rdlo_in(a5_wr[1712]),  .coef_in(coef[512]), .rdup_out(a6_wr[1680]), .rdlo_out(a6_wr[1712]));
			radix2 #(.width(width)) rd_st5_1681  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1681]), .rdlo_in(a5_wr[1713]),  .coef_in(coef[544]), .rdup_out(a6_wr[1681]), .rdlo_out(a6_wr[1713]));
			radix2 #(.width(width)) rd_st5_1682  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1682]), .rdlo_in(a5_wr[1714]),  .coef_in(coef[576]), .rdup_out(a6_wr[1682]), .rdlo_out(a6_wr[1714]));
			radix2 #(.width(width)) rd_st5_1683  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1683]), .rdlo_in(a5_wr[1715]),  .coef_in(coef[608]), .rdup_out(a6_wr[1683]), .rdlo_out(a6_wr[1715]));
			radix2 #(.width(width)) rd_st5_1684  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1684]), .rdlo_in(a5_wr[1716]),  .coef_in(coef[640]), .rdup_out(a6_wr[1684]), .rdlo_out(a6_wr[1716]));
			radix2 #(.width(width)) rd_st5_1685  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1685]), .rdlo_in(a5_wr[1717]),  .coef_in(coef[672]), .rdup_out(a6_wr[1685]), .rdlo_out(a6_wr[1717]));
			radix2 #(.width(width)) rd_st5_1686  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1686]), .rdlo_in(a5_wr[1718]),  .coef_in(coef[704]), .rdup_out(a6_wr[1686]), .rdlo_out(a6_wr[1718]));
			radix2 #(.width(width)) rd_st5_1687  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1687]), .rdlo_in(a5_wr[1719]),  .coef_in(coef[736]), .rdup_out(a6_wr[1687]), .rdlo_out(a6_wr[1719]));
			radix2 #(.width(width)) rd_st5_1688  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1688]), .rdlo_in(a5_wr[1720]),  .coef_in(coef[768]), .rdup_out(a6_wr[1688]), .rdlo_out(a6_wr[1720]));
			radix2 #(.width(width)) rd_st5_1689  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1689]), .rdlo_in(a5_wr[1721]),  .coef_in(coef[800]), .rdup_out(a6_wr[1689]), .rdlo_out(a6_wr[1721]));
			radix2 #(.width(width)) rd_st5_1690  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1690]), .rdlo_in(a5_wr[1722]),  .coef_in(coef[832]), .rdup_out(a6_wr[1690]), .rdlo_out(a6_wr[1722]));
			radix2 #(.width(width)) rd_st5_1691  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1691]), .rdlo_in(a5_wr[1723]),  .coef_in(coef[864]), .rdup_out(a6_wr[1691]), .rdlo_out(a6_wr[1723]));
			radix2 #(.width(width)) rd_st5_1692  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1692]), .rdlo_in(a5_wr[1724]),  .coef_in(coef[896]), .rdup_out(a6_wr[1692]), .rdlo_out(a6_wr[1724]));
			radix2 #(.width(width)) rd_st5_1693  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1693]), .rdlo_in(a5_wr[1725]),  .coef_in(coef[928]), .rdup_out(a6_wr[1693]), .rdlo_out(a6_wr[1725]));
			radix2 #(.width(width)) rd_st5_1694  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1694]), .rdlo_in(a5_wr[1726]),  .coef_in(coef[960]), .rdup_out(a6_wr[1694]), .rdlo_out(a6_wr[1726]));
			radix2 #(.width(width)) rd_st5_1695  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1695]), .rdlo_in(a5_wr[1727]),  .coef_in(coef[992]), .rdup_out(a6_wr[1695]), .rdlo_out(a6_wr[1727]));
			radix2 #(.width(width)) rd_st5_1728  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1728]), .rdlo_in(a5_wr[1760]),  .coef_in(coef[0]), .rdup_out(a6_wr[1728]), .rdlo_out(a6_wr[1760]));
			radix2 #(.width(width)) rd_st5_1729  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1729]), .rdlo_in(a5_wr[1761]),  .coef_in(coef[32]), .rdup_out(a6_wr[1729]), .rdlo_out(a6_wr[1761]));
			radix2 #(.width(width)) rd_st5_1730  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1730]), .rdlo_in(a5_wr[1762]),  .coef_in(coef[64]), .rdup_out(a6_wr[1730]), .rdlo_out(a6_wr[1762]));
			radix2 #(.width(width)) rd_st5_1731  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1731]), .rdlo_in(a5_wr[1763]),  .coef_in(coef[96]), .rdup_out(a6_wr[1731]), .rdlo_out(a6_wr[1763]));
			radix2 #(.width(width)) rd_st5_1732  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1732]), .rdlo_in(a5_wr[1764]),  .coef_in(coef[128]), .rdup_out(a6_wr[1732]), .rdlo_out(a6_wr[1764]));
			radix2 #(.width(width)) rd_st5_1733  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1733]), .rdlo_in(a5_wr[1765]),  .coef_in(coef[160]), .rdup_out(a6_wr[1733]), .rdlo_out(a6_wr[1765]));
			radix2 #(.width(width)) rd_st5_1734  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1734]), .rdlo_in(a5_wr[1766]),  .coef_in(coef[192]), .rdup_out(a6_wr[1734]), .rdlo_out(a6_wr[1766]));
			radix2 #(.width(width)) rd_st5_1735  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1735]), .rdlo_in(a5_wr[1767]),  .coef_in(coef[224]), .rdup_out(a6_wr[1735]), .rdlo_out(a6_wr[1767]));
			radix2 #(.width(width)) rd_st5_1736  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1736]), .rdlo_in(a5_wr[1768]),  .coef_in(coef[256]), .rdup_out(a6_wr[1736]), .rdlo_out(a6_wr[1768]));
			radix2 #(.width(width)) rd_st5_1737  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1737]), .rdlo_in(a5_wr[1769]),  .coef_in(coef[288]), .rdup_out(a6_wr[1737]), .rdlo_out(a6_wr[1769]));
			radix2 #(.width(width)) rd_st5_1738  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1738]), .rdlo_in(a5_wr[1770]),  .coef_in(coef[320]), .rdup_out(a6_wr[1738]), .rdlo_out(a6_wr[1770]));
			radix2 #(.width(width)) rd_st5_1739  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1739]), .rdlo_in(a5_wr[1771]),  .coef_in(coef[352]), .rdup_out(a6_wr[1739]), .rdlo_out(a6_wr[1771]));
			radix2 #(.width(width)) rd_st5_1740  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1740]), .rdlo_in(a5_wr[1772]),  .coef_in(coef[384]), .rdup_out(a6_wr[1740]), .rdlo_out(a6_wr[1772]));
			radix2 #(.width(width)) rd_st5_1741  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1741]), .rdlo_in(a5_wr[1773]),  .coef_in(coef[416]), .rdup_out(a6_wr[1741]), .rdlo_out(a6_wr[1773]));
			radix2 #(.width(width)) rd_st5_1742  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1742]), .rdlo_in(a5_wr[1774]),  .coef_in(coef[448]), .rdup_out(a6_wr[1742]), .rdlo_out(a6_wr[1774]));
			radix2 #(.width(width)) rd_st5_1743  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1743]), .rdlo_in(a5_wr[1775]),  .coef_in(coef[480]), .rdup_out(a6_wr[1743]), .rdlo_out(a6_wr[1775]));
			radix2 #(.width(width)) rd_st5_1744  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1744]), .rdlo_in(a5_wr[1776]),  .coef_in(coef[512]), .rdup_out(a6_wr[1744]), .rdlo_out(a6_wr[1776]));
			radix2 #(.width(width)) rd_st5_1745  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1745]), .rdlo_in(a5_wr[1777]),  .coef_in(coef[544]), .rdup_out(a6_wr[1745]), .rdlo_out(a6_wr[1777]));
			radix2 #(.width(width)) rd_st5_1746  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1746]), .rdlo_in(a5_wr[1778]),  .coef_in(coef[576]), .rdup_out(a6_wr[1746]), .rdlo_out(a6_wr[1778]));
			radix2 #(.width(width)) rd_st5_1747  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1747]), .rdlo_in(a5_wr[1779]),  .coef_in(coef[608]), .rdup_out(a6_wr[1747]), .rdlo_out(a6_wr[1779]));
			radix2 #(.width(width)) rd_st5_1748  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1748]), .rdlo_in(a5_wr[1780]),  .coef_in(coef[640]), .rdup_out(a6_wr[1748]), .rdlo_out(a6_wr[1780]));
			radix2 #(.width(width)) rd_st5_1749  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1749]), .rdlo_in(a5_wr[1781]),  .coef_in(coef[672]), .rdup_out(a6_wr[1749]), .rdlo_out(a6_wr[1781]));
			radix2 #(.width(width)) rd_st5_1750  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1750]), .rdlo_in(a5_wr[1782]),  .coef_in(coef[704]), .rdup_out(a6_wr[1750]), .rdlo_out(a6_wr[1782]));
			radix2 #(.width(width)) rd_st5_1751  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1751]), .rdlo_in(a5_wr[1783]),  .coef_in(coef[736]), .rdup_out(a6_wr[1751]), .rdlo_out(a6_wr[1783]));
			radix2 #(.width(width)) rd_st5_1752  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1752]), .rdlo_in(a5_wr[1784]),  .coef_in(coef[768]), .rdup_out(a6_wr[1752]), .rdlo_out(a6_wr[1784]));
			radix2 #(.width(width)) rd_st5_1753  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1753]), .rdlo_in(a5_wr[1785]),  .coef_in(coef[800]), .rdup_out(a6_wr[1753]), .rdlo_out(a6_wr[1785]));
			radix2 #(.width(width)) rd_st5_1754  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1754]), .rdlo_in(a5_wr[1786]),  .coef_in(coef[832]), .rdup_out(a6_wr[1754]), .rdlo_out(a6_wr[1786]));
			radix2 #(.width(width)) rd_st5_1755  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1755]), .rdlo_in(a5_wr[1787]),  .coef_in(coef[864]), .rdup_out(a6_wr[1755]), .rdlo_out(a6_wr[1787]));
			radix2 #(.width(width)) rd_st5_1756  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1756]), .rdlo_in(a5_wr[1788]),  .coef_in(coef[896]), .rdup_out(a6_wr[1756]), .rdlo_out(a6_wr[1788]));
			radix2 #(.width(width)) rd_st5_1757  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1757]), .rdlo_in(a5_wr[1789]),  .coef_in(coef[928]), .rdup_out(a6_wr[1757]), .rdlo_out(a6_wr[1789]));
			radix2 #(.width(width)) rd_st5_1758  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1758]), .rdlo_in(a5_wr[1790]),  .coef_in(coef[960]), .rdup_out(a6_wr[1758]), .rdlo_out(a6_wr[1790]));
			radix2 #(.width(width)) rd_st5_1759  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1759]), .rdlo_in(a5_wr[1791]),  .coef_in(coef[992]), .rdup_out(a6_wr[1759]), .rdlo_out(a6_wr[1791]));
			radix2 #(.width(width)) rd_st5_1792  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1792]), .rdlo_in(a5_wr[1824]),  .coef_in(coef[0]), .rdup_out(a6_wr[1792]), .rdlo_out(a6_wr[1824]));
			radix2 #(.width(width)) rd_st5_1793  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1793]), .rdlo_in(a5_wr[1825]),  .coef_in(coef[32]), .rdup_out(a6_wr[1793]), .rdlo_out(a6_wr[1825]));
			radix2 #(.width(width)) rd_st5_1794  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1794]), .rdlo_in(a5_wr[1826]),  .coef_in(coef[64]), .rdup_out(a6_wr[1794]), .rdlo_out(a6_wr[1826]));
			radix2 #(.width(width)) rd_st5_1795  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1795]), .rdlo_in(a5_wr[1827]),  .coef_in(coef[96]), .rdup_out(a6_wr[1795]), .rdlo_out(a6_wr[1827]));
			radix2 #(.width(width)) rd_st5_1796  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1796]), .rdlo_in(a5_wr[1828]),  .coef_in(coef[128]), .rdup_out(a6_wr[1796]), .rdlo_out(a6_wr[1828]));
			radix2 #(.width(width)) rd_st5_1797  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1797]), .rdlo_in(a5_wr[1829]),  .coef_in(coef[160]), .rdup_out(a6_wr[1797]), .rdlo_out(a6_wr[1829]));
			radix2 #(.width(width)) rd_st5_1798  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1798]), .rdlo_in(a5_wr[1830]),  .coef_in(coef[192]), .rdup_out(a6_wr[1798]), .rdlo_out(a6_wr[1830]));
			radix2 #(.width(width)) rd_st5_1799  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1799]), .rdlo_in(a5_wr[1831]),  .coef_in(coef[224]), .rdup_out(a6_wr[1799]), .rdlo_out(a6_wr[1831]));
			radix2 #(.width(width)) rd_st5_1800  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1800]), .rdlo_in(a5_wr[1832]),  .coef_in(coef[256]), .rdup_out(a6_wr[1800]), .rdlo_out(a6_wr[1832]));
			radix2 #(.width(width)) rd_st5_1801  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1801]), .rdlo_in(a5_wr[1833]),  .coef_in(coef[288]), .rdup_out(a6_wr[1801]), .rdlo_out(a6_wr[1833]));
			radix2 #(.width(width)) rd_st5_1802  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1802]), .rdlo_in(a5_wr[1834]),  .coef_in(coef[320]), .rdup_out(a6_wr[1802]), .rdlo_out(a6_wr[1834]));
			radix2 #(.width(width)) rd_st5_1803  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1803]), .rdlo_in(a5_wr[1835]),  .coef_in(coef[352]), .rdup_out(a6_wr[1803]), .rdlo_out(a6_wr[1835]));
			radix2 #(.width(width)) rd_st5_1804  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1804]), .rdlo_in(a5_wr[1836]),  .coef_in(coef[384]), .rdup_out(a6_wr[1804]), .rdlo_out(a6_wr[1836]));
			radix2 #(.width(width)) rd_st5_1805  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1805]), .rdlo_in(a5_wr[1837]),  .coef_in(coef[416]), .rdup_out(a6_wr[1805]), .rdlo_out(a6_wr[1837]));
			radix2 #(.width(width)) rd_st5_1806  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1806]), .rdlo_in(a5_wr[1838]),  .coef_in(coef[448]), .rdup_out(a6_wr[1806]), .rdlo_out(a6_wr[1838]));
			radix2 #(.width(width)) rd_st5_1807  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1807]), .rdlo_in(a5_wr[1839]),  .coef_in(coef[480]), .rdup_out(a6_wr[1807]), .rdlo_out(a6_wr[1839]));
			radix2 #(.width(width)) rd_st5_1808  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1808]), .rdlo_in(a5_wr[1840]),  .coef_in(coef[512]), .rdup_out(a6_wr[1808]), .rdlo_out(a6_wr[1840]));
			radix2 #(.width(width)) rd_st5_1809  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1809]), .rdlo_in(a5_wr[1841]),  .coef_in(coef[544]), .rdup_out(a6_wr[1809]), .rdlo_out(a6_wr[1841]));
			radix2 #(.width(width)) rd_st5_1810  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1810]), .rdlo_in(a5_wr[1842]),  .coef_in(coef[576]), .rdup_out(a6_wr[1810]), .rdlo_out(a6_wr[1842]));
			radix2 #(.width(width)) rd_st5_1811  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1811]), .rdlo_in(a5_wr[1843]),  .coef_in(coef[608]), .rdup_out(a6_wr[1811]), .rdlo_out(a6_wr[1843]));
			radix2 #(.width(width)) rd_st5_1812  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1812]), .rdlo_in(a5_wr[1844]),  .coef_in(coef[640]), .rdup_out(a6_wr[1812]), .rdlo_out(a6_wr[1844]));
			radix2 #(.width(width)) rd_st5_1813  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1813]), .rdlo_in(a5_wr[1845]),  .coef_in(coef[672]), .rdup_out(a6_wr[1813]), .rdlo_out(a6_wr[1845]));
			radix2 #(.width(width)) rd_st5_1814  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1814]), .rdlo_in(a5_wr[1846]),  .coef_in(coef[704]), .rdup_out(a6_wr[1814]), .rdlo_out(a6_wr[1846]));
			radix2 #(.width(width)) rd_st5_1815  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1815]), .rdlo_in(a5_wr[1847]),  .coef_in(coef[736]), .rdup_out(a6_wr[1815]), .rdlo_out(a6_wr[1847]));
			radix2 #(.width(width)) rd_st5_1816  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1816]), .rdlo_in(a5_wr[1848]),  .coef_in(coef[768]), .rdup_out(a6_wr[1816]), .rdlo_out(a6_wr[1848]));
			radix2 #(.width(width)) rd_st5_1817  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1817]), .rdlo_in(a5_wr[1849]),  .coef_in(coef[800]), .rdup_out(a6_wr[1817]), .rdlo_out(a6_wr[1849]));
			radix2 #(.width(width)) rd_st5_1818  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1818]), .rdlo_in(a5_wr[1850]),  .coef_in(coef[832]), .rdup_out(a6_wr[1818]), .rdlo_out(a6_wr[1850]));
			radix2 #(.width(width)) rd_st5_1819  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1819]), .rdlo_in(a5_wr[1851]),  .coef_in(coef[864]), .rdup_out(a6_wr[1819]), .rdlo_out(a6_wr[1851]));
			radix2 #(.width(width)) rd_st5_1820  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1820]), .rdlo_in(a5_wr[1852]),  .coef_in(coef[896]), .rdup_out(a6_wr[1820]), .rdlo_out(a6_wr[1852]));
			radix2 #(.width(width)) rd_st5_1821  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1821]), .rdlo_in(a5_wr[1853]),  .coef_in(coef[928]), .rdup_out(a6_wr[1821]), .rdlo_out(a6_wr[1853]));
			radix2 #(.width(width)) rd_st5_1822  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1822]), .rdlo_in(a5_wr[1854]),  .coef_in(coef[960]), .rdup_out(a6_wr[1822]), .rdlo_out(a6_wr[1854]));
			radix2 #(.width(width)) rd_st5_1823  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1823]), .rdlo_in(a5_wr[1855]),  .coef_in(coef[992]), .rdup_out(a6_wr[1823]), .rdlo_out(a6_wr[1855]));
			radix2 #(.width(width)) rd_st5_1856  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1856]), .rdlo_in(a5_wr[1888]),  .coef_in(coef[0]), .rdup_out(a6_wr[1856]), .rdlo_out(a6_wr[1888]));
			radix2 #(.width(width)) rd_st5_1857  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1857]), .rdlo_in(a5_wr[1889]),  .coef_in(coef[32]), .rdup_out(a6_wr[1857]), .rdlo_out(a6_wr[1889]));
			radix2 #(.width(width)) rd_st5_1858  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1858]), .rdlo_in(a5_wr[1890]),  .coef_in(coef[64]), .rdup_out(a6_wr[1858]), .rdlo_out(a6_wr[1890]));
			radix2 #(.width(width)) rd_st5_1859  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1859]), .rdlo_in(a5_wr[1891]),  .coef_in(coef[96]), .rdup_out(a6_wr[1859]), .rdlo_out(a6_wr[1891]));
			radix2 #(.width(width)) rd_st5_1860  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1860]), .rdlo_in(a5_wr[1892]),  .coef_in(coef[128]), .rdup_out(a6_wr[1860]), .rdlo_out(a6_wr[1892]));
			radix2 #(.width(width)) rd_st5_1861  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1861]), .rdlo_in(a5_wr[1893]),  .coef_in(coef[160]), .rdup_out(a6_wr[1861]), .rdlo_out(a6_wr[1893]));
			radix2 #(.width(width)) rd_st5_1862  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1862]), .rdlo_in(a5_wr[1894]),  .coef_in(coef[192]), .rdup_out(a6_wr[1862]), .rdlo_out(a6_wr[1894]));
			radix2 #(.width(width)) rd_st5_1863  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1863]), .rdlo_in(a5_wr[1895]),  .coef_in(coef[224]), .rdup_out(a6_wr[1863]), .rdlo_out(a6_wr[1895]));
			radix2 #(.width(width)) rd_st5_1864  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1864]), .rdlo_in(a5_wr[1896]),  .coef_in(coef[256]), .rdup_out(a6_wr[1864]), .rdlo_out(a6_wr[1896]));
			radix2 #(.width(width)) rd_st5_1865  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1865]), .rdlo_in(a5_wr[1897]),  .coef_in(coef[288]), .rdup_out(a6_wr[1865]), .rdlo_out(a6_wr[1897]));
			radix2 #(.width(width)) rd_st5_1866  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1866]), .rdlo_in(a5_wr[1898]),  .coef_in(coef[320]), .rdup_out(a6_wr[1866]), .rdlo_out(a6_wr[1898]));
			radix2 #(.width(width)) rd_st5_1867  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1867]), .rdlo_in(a5_wr[1899]),  .coef_in(coef[352]), .rdup_out(a6_wr[1867]), .rdlo_out(a6_wr[1899]));
			radix2 #(.width(width)) rd_st5_1868  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1868]), .rdlo_in(a5_wr[1900]),  .coef_in(coef[384]), .rdup_out(a6_wr[1868]), .rdlo_out(a6_wr[1900]));
			radix2 #(.width(width)) rd_st5_1869  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1869]), .rdlo_in(a5_wr[1901]),  .coef_in(coef[416]), .rdup_out(a6_wr[1869]), .rdlo_out(a6_wr[1901]));
			radix2 #(.width(width)) rd_st5_1870  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1870]), .rdlo_in(a5_wr[1902]),  .coef_in(coef[448]), .rdup_out(a6_wr[1870]), .rdlo_out(a6_wr[1902]));
			radix2 #(.width(width)) rd_st5_1871  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1871]), .rdlo_in(a5_wr[1903]),  .coef_in(coef[480]), .rdup_out(a6_wr[1871]), .rdlo_out(a6_wr[1903]));
			radix2 #(.width(width)) rd_st5_1872  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1872]), .rdlo_in(a5_wr[1904]),  .coef_in(coef[512]), .rdup_out(a6_wr[1872]), .rdlo_out(a6_wr[1904]));
			radix2 #(.width(width)) rd_st5_1873  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1873]), .rdlo_in(a5_wr[1905]),  .coef_in(coef[544]), .rdup_out(a6_wr[1873]), .rdlo_out(a6_wr[1905]));
			radix2 #(.width(width)) rd_st5_1874  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1874]), .rdlo_in(a5_wr[1906]),  .coef_in(coef[576]), .rdup_out(a6_wr[1874]), .rdlo_out(a6_wr[1906]));
			radix2 #(.width(width)) rd_st5_1875  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1875]), .rdlo_in(a5_wr[1907]),  .coef_in(coef[608]), .rdup_out(a6_wr[1875]), .rdlo_out(a6_wr[1907]));
			radix2 #(.width(width)) rd_st5_1876  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1876]), .rdlo_in(a5_wr[1908]),  .coef_in(coef[640]), .rdup_out(a6_wr[1876]), .rdlo_out(a6_wr[1908]));
			radix2 #(.width(width)) rd_st5_1877  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1877]), .rdlo_in(a5_wr[1909]),  .coef_in(coef[672]), .rdup_out(a6_wr[1877]), .rdlo_out(a6_wr[1909]));
			radix2 #(.width(width)) rd_st5_1878  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1878]), .rdlo_in(a5_wr[1910]),  .coef_in(coef[704]), .rdup_out(a6_wr[1878]), .rdlo_out(a6_wr[1910]));
			radix2 #(.width(width)) rd_st5_1879  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1879]), .rdlo_in(a5_wr[1911]),  .coef_in(coef[736]), .rdup_out(a6_wr[1879]), .rdlo_out(a6_wr[1911]));
			radix2 #(.width(width)) rd_st5_1880  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1880]), .rdlo_in(a5_wr[1912]),  .coef_in(coef[768]), .rdup_out(a6_wr[1880]), .rdlo_out(a6_wr[1912]));
			radix2 #(.width(width)) rd_st5_1881  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1881]), .rdlo_in(a5_wr[1913]),  .coef_in(coef[800]), .rdup_out(a6_wr[1881]), .rdlo_out(a6_wr[1913]));
			radix2 #(.width(width)) rd_st5_1882  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1882]), .rdlo_in(a5_wr[1914]),  .coef_in(coef[832]), .rdup_out(a6_wr[1882]), .rdlo_out(a6_wr[1914]));
			radix2 #(.width(width)) rd_st5_1883  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1883]), .rdlo_in(a5_wr[1915]),  .coef_in(coef[864]), .rdup_out(a6_wr[1883]), .rdlo_out(a6_wr[1915]));
			radix2 #(.width(width)) rd_st5_1884  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1884]), .rdlo_in(a5_wr[1916]),  .coef_in(coef[896]), .rdup_out(a6_wr[1884]), .rdlo_out(a6_wr[1916]));
			radix2 #(.width(width)) rd_st5_1885  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1885]), .rdlo_in(a5_wr[1917]),  .coef_in(coef[928]), .rdup_out(a6_wr[1885]), .rdlo_out(a6_wr[1917]));
			radix2 #(.width(width)) rd_st5_1886  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1886]), .rdlo_in(a5_wr[1918]),  .coef_in(coef[960]), .rdup_out(a6_wr[1886]), .rdlo_out(a6_wr[1918]));
			radix2 #(.width(width)) rd_st5_1887  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1887]), .rdlo_in(a5_wr[1919]),  .coef_in(coef[992]), .rdup_out(a6_wr[1887]), .rdlo_out(a6_wr[1919]));
			radix2 #(.width(width)) rd_st5_1920  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1920]), .rdlo_in(a5_wr[1952]),  .coef_in(coef[0]), .rdup_out(a6_wr[1920]), .rdlo_out(a6_wr[1952]));
			radix2 #(.width(width)) rd_st5_1921  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1921]), .rdlo_in(a5_wr[1953]),  .coef_in(coef[32]), .rdup_out(a6_wr[1921]), .rdlo_out(a6_wr[1953]));
			radix2 #(.width(width)) rd_st5_1922  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1922]), .rdlo_in(a5_wr[1954]),  .coef_in(coef[64]), .rdup_out(a6_wr[1922]), .rdlo_out(a6_wr[1954]));
			radix2 #(.width(width)) rd_st5_1923  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1923]), .rdlo_in(a5_wr[1955]),  .coef_in(coef[96]), .rdup_out(a6_wr[1923]), .rdlo_out(a6_wr[1955]));
			radix2 #(.width(width)) rd_st5_1924  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1924]), .rdlo_in(a5_wr[1956]),  .coef_in(coef[128]), .rdup_out(a6_wr[1924]), .rdlo_out(a6_wr[1956]));
			radix2 #(.width(width)) rd_st5_1925  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1925]), .rdlo_in(a5_wr[1957]),  .coef_in(coef[160]), .rdup_out(a6_wr[1925]), .rdlo_out(a6_wr[1957]));
			radix2 #(.width(width)) rd_st5_1926  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1926]), .rdlo_in(a5_wr[1958]),  .coef_in(coef[192]), .rdup_out(a6_wr[1926]), .rdlo_out(a6_wr[1958]));
			radix2 #(.width(width)) rd_st5_1927  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1927]), .rdlo_in(a5_wr[1959]),  .coef_in(coef[224]), .rdup_out(a6_wr[1927]), .rdlo_out(a6_wr[1959]));
			radix2 #(.width(width)) rd_st5_1928  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1928]), .rdlo_in(a5_wr[1960]),  .coef_in(coef[256]), .rdup_out(a6_wr[1928]), .rdlo_out(a6_wr[1960]));
			radix2 #(.width(width)) rd_st5_1929  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1929]), .rdlo_in(a5_wr[1961]),  .coef_in(coef[288]), .rdup_out(a6_wr[1929]), .rdlo_out(a6_wr[1961]));
			radix2 #(.width(width)) rd_st5_1930  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1930]), .rdlo_in(a5_wr[1962]),  .coef_in(coef[320]), .rdup_out(a6_wr[1930]), .rdlo_out(a6_wr[1962]));
			radix2 #(.width(width)) rd_st5_1931  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1931]), .rdlo_in(a5_wr[1963]),  .coef_in(coef[352]), .rdup_out(a6_wr[1931]), .rdlo_out(a6_wr[1963]));
			radix2 #(.width(width)) rd_st5_1932  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1932]), .rdlo_in(a5_wr[1964]),  .coef_in(coef[384]), .rdup_out(a6_wr[1932]), .rdlo_out(a6_wr[1964]));
			radix2 #(.width(width)) rd_st5_1933  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1933]), .rdlo_in(a5_wr[1965]),  .coef_in(coef[416]), .rdup_out(a6_wr[1933]), .rdlo_out(a6_wr[1965]));
			radix2 #(.width(width)) rd_st5_1934  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1934]), .rdlo_in(a5_wr[1966]),  .coef_in(coef[448]), .rdup_out(a6_wr[1934]), .rdlo_out(a6_wr[1966]));
			radix2 #(.width(width)) rd_st5_1935  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1935]), .rdlo_in(a5_wr[1967]),  .coef_in(coef[480]), .rdup_out(a6_wr[1935]), .rdlo_out(a6_wr[1967]));
			radix2 #(.width(width)) rd_st5_1936  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1936]), .rdlo_in(a5_wr[1968]),  .coef_in(coef[512]), .rdup_out(a6_wr[1936]), .rdlo_out(a6_wr[1968]));
			radix2 #(.width(width)) rd_st5_1937  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1937]), .rdlo_in(a5_wr[1969]),  .coef_in(coef[544]), .rdup_out(a6_wr[1937]), .rdlo_out(a6_wr[1969]));
			radix2 #(.width(width)) rd_st5_1938  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1938]), .rdlo_in(a5_wr[1970]),  .coef_in(coef[576]), .rdup_out(a6_wr[1938]), .rdlo_out(a6_wr[1970]));
			radix2 #(.width(width)) rd_st5_1939  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1939]), .rdlo_in(a5_wr[1971]),  .coef_in(coef[608]), .rdup_out(a6_wr[1939]), .rdlo_out(a6_wr[1971]));
			radix2 #(.width(width)) rd_st5_1940  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1940]), .rdlo_in(a5_wr[1972]),  .coef_in(coef[640]), .rdup_out(a6_wr[1940]), .rdlo_out(a6_wr[1972]));
			radix2 #(.width(width)) rd_st5_1941  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1941]), .rdlo_in(a5_wr[1973]),  .coef_in(coef[672]), .rdup_out(a6_wr[1941]), .rdlo_out(a6_wr[1973]));
			radix2 #(.width(width)) rd_st5_1942  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1942]), .rdlo_in(a5_wr[1974]),  .coef_in(coef[704]), .rdup_out(a6_wr[1942]), .rdlo_out(a6_wr[1974]));
			radix2 #(.width(width)) rd_st5_1943  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1943]), .rdlo_in(a5_wr[1975]),  .coef_in(coef[736]), .rdup_out(a6_wr[1943]), .rdlo_out(a6_wr[1975]));
			radix2 #(.width(width)) rd_st5_1944  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1944]), .rdlo_in(a5_wr[1976]),  .coef_in(coef[768]), .rdup_out(a6_wr[1944]), .rdlo_out(a6_wr[1976]));
			radix2 #(.width(width)) rd_st5_1945  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1945]), .rdlo_in(a5_wr[1977]),  .coef_in(coef[800]), .rdup_out(a6_wr[1945]), .rdlo_out(a6_wr[1977]));
			radix2 #(.width(width)) rd_st5_1946  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1946]), .rdlo_in(a5_wr[1978]),  .coef_in(coef[832]), .rdup_out(a6_wr[1946]), .rdlo_out(a6_wr[1978]));
			radix2 #(.width(width)) rd_st5_1947  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1947]), .rdlo_in(a5_wr[1979]),  .coef_in(coef[864]), .rdup_out(a6_wr[1947]), .rdlo_out(a6_wr[1979]));
			radix2 #(.width(width)) rd_st5_1948  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1948]), .rdlo_in(a5_wr[1980]),  .coef_in(coef[896]), .rdup_out(a6_wr[1948]), .rdlo_out(a6_wr[1980]));
			radix2 #(.width(width)) rd_st5_1949  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1949]), .rdlo_in(a5_wr[1981]),  .coef_in(coef[928]), .rdup_out(a6_wr[1949]), .rdlo_out(a6_wr[1981]));
			radix2 #(.width(width)) rd_st5_1950  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1950]), .rdlo_in(a5_wr[1982]),  .coef_in(coef[960]), .rdup_out(a6_wr[1950]), .rdlo_out(a6_wr[1982]));
			radix2 #(.width(width)) rd_st5_1951  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1951]), .rdlo_in(a5_wr[1983]),  .coef_in(coef[992]), .rdup_out(a6_wr[1951]), .rdlo_out(a6_wr[1983]));
			radix2 #(.width(width)) rd_st5_1984  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1984]), .rdlo_in(a5_wr[2016]),  .coef_in(coef[0]), .rdup_out(a6_wr[1984]), .rdlo_out(a6_wr[2016]));
			radix2 #(.width(width)) rd_st5_1985  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1985]), .rdlo_in(a5_wr[2017]),  .coef_in(coef[32]), .rdup_out(a6_wr[1985]), .rdlo_out(a6_wr[2017]));
			radix2 #(.width(width)) rd_st5_1986  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1986]), .rdlo_in(a5_wr[2018]),  .coef_in(coef[64]), .rdup_out(a6_wr[1986]), .rdlo_out(a6_wr[2018]));
			radix2 #(.width(width)) rd_st5_1987  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1987]), .rdlo_in(a5_wr[2019]),  .coef_in(coef[96]), .rdup_out(a6_wr[1987]), .rdlo_out(a6_wr[2019]));
			radix2 #(.width(width)) rd_st5_1988  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1988]), .rdlo_in(a5_wr[2020]),  .coef_in(coef[128]), .rdup_out(a6_wr[1988]), .rdlo_out(a6_wr[2020]));
			radix2 #(.width(width)) rd_st5_1989  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1989]), .rdlo_in(a5_wr[2021]),  .coef_in(coef[160]), .rdup_out(a6_wr[1989]), .rdlo_out(a6_wr[2021]));
			radix2 #(.width(width)) rd_st5_1990  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1990]), .rdlo_in(a5_wr[2022]),  .coef_in(coef[192]), .rdup_out(a6_wr[1990]), .rdlo_out(a6_wr[2022]));
			radix2 #(.width(width)) rd_st5_1991  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1991]), .rdlo_in(a5_wr[2023]),  .coef_in(coef[224]), .rdup_out(a6_wr[1991]), .rdlo_out(a6_wr[2023]));
			radix2 #(.width(width)) rd_st5_1992  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1992]), .rdlo_in(a5_wr[2024]),  .coef_in(coef[256]), .rdup_out(a6_wr[1992]), .rdlo_out(a6_wr[2024]));
			radix2 #(.width(width)) rd_st5_1993  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1993]), .rdlo_in(a5_wr[2025]),  .coef_in(coef[288]), .rdup_out(a6_wr[1993]), .rdlo_out(a6_wr[2025]));
			radix2 #(.width(width)) rd_st5_1994  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1994]), .rdlo_in(a5_wr[2026]),  .coef_in(coef[320]), .rdup_out(a6_wr[1994]), .rdlo_out(a6_wr[2026]));
			radix2 #(.width(width)) rd_st5_1995  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1995]), .rdlo_in(a5_wr[2027]),  .coef_in(coef[352]), .rdup_out(a6_wr[1995]), .rdlo_out(a6_wr[2027]));
			radix2 #(.width(width)) rd_st5_1996  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1996]), .rdlo_in(a5_wr[2028]),  .coef_in(coef[384]), .rdup_out(a6_wr[1996]), .rdlo_out(a6_wr[2028]));
			radix2 #(.width(width)) rd_st5_1997  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1997]), .rdlo_in(a5_wr[2029]),  .coef_in(coef[416]), .rdup_out(a6_wr[1997]), .rdlo_out(a6_wr[2029]));
			radix2 #(.width(width)) rd_st5_1998  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1998]), .rdlo_in(a5_wr[2030]),  .coef_in(coef[448]), .rdup_out(a6_wr[1998]), .rdlo_out(a6_wr[2030]));
			radix2 #(.width(width)) rd_st5_1999  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[1999]), .rdlo_in(a5_wr[2031]),  .coef_in(coef[480]), .rdup_out(a6_wr[1999]), .rdlo_out(a6_wr[2031]));
			radix2 #(.width(width)) rd_st5_2000  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[2000]), .rdlo_in(a5_wr[2032]),  .coef_in(coef[512]), .rdup_out(a6_wr[2000]), .rdlo_out(a6_wr[2032]));
			radix2 #(.width(width)) rd_st5_2001  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[2001]), .rdlo_in(a5_wr[2033]),  .coef_in(coef[544]), .rdup_out(a6_wr[2001]), .rdlo_out(a6_wr[2033]));
			radix2 #(.width(width)) rd_st5_2002  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[2002]), .rdlo_in(a5_wr[2034]),  .coef_in(coef[576]), .rdup_out(a6_wr[2002]), .rdlo_out(a6_wr[2034]));
			radix2 #(.width(width)) rd_st5_2003  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[2003]), .rdlo_in(a5_wr[2035]),  .coef_in(coef[608]), .rdup_out(a6_wr[2003]), .rdlo_out(a6_wr[2035]));
			radix2 #(.width(width)) rd_st5_2004  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[2004]), .rdlo_in(a5_wr[2036]),  .coef_in(coef[640]), .rdup_out(a6_wr[2004]), .rdlo_out(a6_wr[2036]));
			radix2 #(.width(width)) rd_st5_2005  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[2005]), .rdlo_in(a5_wr[2037]),  .coef_in(coef[672]), .rdup_out(a6_wr[2005]), .rdlo_out(a6_wr[2037]));
			radix2 #(.width(width)) rd_st5_2006  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[2006]), .rdlo_in(a5_wr[2038]),  .coef_in(coef[704]), .rdup_out(a6_wr[2006]), .rdlo_out(a6_wr[2038]));
			radix2 #(.width(width)) rd_st5_2007  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[2007]), .rdlo_in(a5_wr[2039]),  .coef_in(coef[736]), .rdup_out(a6_wr[2007]), .rdlo_out(a6_wr[2039]));
			radix2 #(.width(width)) rd_st5_2008  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[2008]), .rdlo_in(a5_wr[2040]),  .coef_in(coef[768]), .rdup_out(a6_wr[2008]), .rdlo_out(a6_wr[2040]));
			radix2 #(.width(width)) rd_st5_2009  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[2009]), .rdlo_in(a5_wr[2041]),  .coef_in(coef[800]), .rdup_out(a6_wr[2009]), .rdlo_out(a6_wr[2041]));
			radix2 #(.width(width)) rd_st5_2010  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[2010]), .rdlo_in(a5_wr[2042]),  .coef_in(coef[832]), .rdup_out(a6_wr[2010]), .rdlo_out(a6_wr[2042]));
			radix2 #(.width(width)) rd_st5_2011  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[2011]), .rdlo_in(a5_wr[2043]),  .coef_in(coef[864]), .rdup_out(a6_wr[2011]), .rdlo_out(a6_wr[2043]));
			radix2 #(.width(width)) rd_st5_2012  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[2012]), .rdlo_in(a5_wr[2044]),  .coef_in(coef[896]), .rdup_out(a6_wr[2012]), .rdlo_out(a6_wr[2044]));
			radix2 #(.width(width)) rd_st5_2013  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[2013]), .rdlo_in(a5_wr[2045]),  .coef_in(coef[928]), .rdup_out(a6_wr[2013]), .rdlo_out(a6_wr[2045]));
			radix2 #(.width(width)) rd_st5_2014  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[2014]), .rdlo_in(a5_wr[2046]),  .coef_in(coef[960]), .rdup_out(a6_wr[2014]), .rdlo_out(a6_wr[2046]));
			radix2 #(.width(width)) rd_st5_2015  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a5_wr[2015]), .rdlo_in(a5_wr[2047]),  .coef_in(coef[992]), .rdup_out(a6_wr[2015]), .rdlo_out(a6_wr[2047]));

		//--- radix stage 6
			radix2 #(.width(width)) rd_st6_0   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[0]), .rdlo_in(a6_wr[16]),  .coef_in(coef[0]), .rdup_out(a7_wr[0]), .rdlo_out(a7_wr[16]));
			radix2 #(.width(width)) rd_st6_1   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1]), .rdlo_in(a6_wr[17]),  .coef_in(coef[64]), .rdup_out(a7_wr[1]), .rdlo_out(a7_wr[17]));
			radix2 #(.width(width)) rd_st6_2   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[2]), .rdlo_in(a6_wr[18]),  .coef_in(coef[128]), .rdup_out(a7_wr[2]), .rdlo_out(a7_wr[18]));
			radix2 #(.width(width)) rd_st6_3   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[3]), .rdlo_in(a6_wr[19]),  .coef_in(coef[192]), .rdup_out(a7_wr[3]), .rdlo_out(a7_wr[19]));
			radix2 #(.width(width)) rd_st6_4   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[4]), .rdlo_in(a6_wr[20]),  .coef_in(coef[256]), .rdup_out(a7_wr[4]), .rdlo_out(a7_wr[20]));
			radix2 #(.width(width)) rd_st6_5   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[5]), .rdlo_in(a6_wr[21]),  .coef_in(coef[320]), .rdup_out(a7_wr[5]), .rdlo_out(a7_wr[21]));
			radix2 #(.width(width)) rd_st6_6   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[6]), .rdlo_in(a6_wr[22]),  .coef_in(coef[384]), .rdup_out(a7_wr[6]), .rdlo_out(a7_wr[22]));
			radix2 #(.width(width)) rd_st6_7   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[7]), .rdlo_in(a6_wr[23]),  .coef_in(coef[448]), .rdup_out(a7_wr[7]), .rdlo_out(a7_wr[23]));
			radix2 #(.width(width)) rd_st6_8   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[8]), .rdlo_in(a6_wr[24]),  .coef_in(coef[512]), .rdup_out(a7_wr[8]), .rdlo_out(a7_wr[24]));
			radix2 #(.width(width)) rd_st6_9   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[9]), .rdlo_in(a6_wr[25]),  .coef_in(coef[576]), .rdup_out(a7_wr[9]), .rdlo_out(a7_wr[25]));
			radix2 #(.width(width)) rd_st6_10  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[10]), .rdlo_in(a6_wr[26]),  .coef_in(coef[640]), .rdup_out(a7_wr[10]), .rdlo_out(a7_wr[26]));
			radix2 #(.width(width)) rd_st6_11  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[11]), .rdlo_in(a6_wr[27]),  .coef_in(coef[704]), .rdup_out(a7_wr[11]), .rdlo_out(a7_wr[27]));
			radix2 #(.width(width)) rd_st6_12  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[12]), .rdlo_in(a6_wr[28]),  .coef_in(coef[768]), .rdup_out(a7_wr[12]), .rdlo_out(a7_wr[28]));
			radix2 #(.width(width)) rd_st6_13  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[13]), .rdlo_in(a6_wr[29]),  .coef_in(coef[832]), .rdup_out(a7_wr[13]), .rdlo_out(a7_wr[29]));
			radix2 #(.width(width)) rd_st6_14  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[14]), .rdlo_in(a6_wr[30]),  .coef_in(coef[896]), .rdup_out(a7_wr[14]), .rdlo_out(a7_wr[30]));
			radix2 #(.width(width)) rd_st6_15  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[15]), .rdlo_in(a6_wr[31]),  .coef_in(coef[960]), .rdup_out(a7_wr[15]), .rdlo_out(a7_wr[31]));
			radix2 #(.width(width)) rd_st6_32  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[32]), .rdlo_in(a6_wr[48]),  .coef_in(coef[0]), .rdup_out(a7_wr[32]), .rdlo_out(a7_wr[48]));
			radix2 #(.width(width)) rd_st6_33  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[33]), .rdlo_in(a6_wr[49]),  .coef_in(coef[64]), .rdup_out(a7_wr[33]), .rdlo_out(a7_wr[49]));
			radix2 #(.width(width)) rd_st6_34  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[34]), .rdlo_in(a6_wr[50]),  .coef_in(coef[128]), .rdup_out(a7_wr[34]), .rdlo_out(a7_wr[50]));
			radix2 #(.width(width)) rd_st6_35  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[35]), .rdlo_in(a6_wr[51]),  .coef_in(coef[192]), .rdup_out(a7_wr[35]), .rdlo_out(a7_wr[51]));
			radix2 #(.width(width)) rd_st6_36  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[36]), .rdlo_in(a6_wr[52]),  .coef_in(coef[256]), .rdup_out(a7_wr[36]), .rdlo_out(a7_wr[52]));
			radix2 #(.width(width)) rd_st6_37  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[37]), .rdlo_in(a6_wr[53]),  .coef_in(coef[320]), .rdup_out(a7_wr[37]), .rdlo_out(a7_wr[53]));
			radix2 #(.width(width)) rd_st6_38  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[38]), .rdlo_in(a6_wr[54]),  .coef_in(coef[384]), .rdup_out(a7_wr[38]), .rdlo_out(a7_wr[54]));
			radix2 #(.width(width)) rd_st6_39  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[39]), .rdlo_in(a6_wr[55]),  .coef_in(coef[448]), .rdup_out(a7_wr[39]), .rdlo_out(a7_wr[55]));
			radix2 #(.width(width)) rd_st6_40  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[40]), .rdlo_in(a6_wr[56]),  .coef_in(coef[512]), .rdup_out(a7_wr[40]), .rdlo_out(a7_wr[56]));
			radix2 #(.width(width)) rd_st6_41  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[41]), .rdlo_in(a6_wr[57]),  .coef_in(coef[576]), .rdup_out(a7_wr[41]), .rdlo_out(a7_wr[57]));
			radix2 #(.width(width)) rd_st6_42  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[42]), .rdlo_in(a6_wr[58]),  .coef_in(coef[640]), .rdup_out(a7_wr[42]), .rdlo_out(a7_wr[58]));
			radix2 #(.width(width)) rd_st6_43  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[43]), .rdlo_in(a6_wr[59]),  .coef_in(coef[704]), .rdup_out(a7_wr[43]), .rdlo_out(a7_wr[59]));
			radix2 #(.width(width)) rd_st6_44  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[44]), .rdlo_in(a6_wr[60]),  .coef_in(coef[768]), .rdup_out(a7_wr[44]), .rdlo_out(a7_wr[60]));
			radix2 #(.width(width)) rd_st6_45  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[45]), .rdlo_in(a6_wr[61]),  .coef_in(coef[832]), .rdup_out(a7_wr[45]), .rdlo_out(a7_wr[61]));
			radix2 #(.width(width)) rd_st6_46  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[46]), .rdlo_in(a6_wr[62]),  .coef_in(coef[896]), .rdup_out(a7_wr[46]), .rdlo_out(a7_wr[62]));
			radix2 #(.width(width)) rd_st6_47  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[47]), .rdlo_in(a6_wr[63]),  .coef_in(coef[960]), .rdup_out(a7_wr[47]), .rdlo_out(a7_wr[63]));
			radix2 #(.width(width)) rd_st6_64  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[64]), .rdlo_in(a6_wr[80]),  .coef_in(coef[0]), .rdup_out(a7_wr[64]), .rdlo_out(a7_wr[80]));
			radix2 #(.width(width)) rd_st6_65  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[65]), .rdlo_in(a6_wr[81]),  .coef_in(coef[64]), .rdup_out(a7_wr[65]), .rdlo_out(a7_wr[81]));
			radix2 #(.width(width)) rd_st6_66  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[66]), .rdlo_in(a6_wr[82]),  .coef_in(coef[128]), .rdup_out(a7_wr[66]), .rdlo_out(a7_wr[82]));
			radix2 #(.width(width)) rd_st6_67  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[67]), .rdlo_in(a6_wr[83]),  .coef_in(coef[192]), .rdup_out(a7_wr[67]), .rdlo_out(a7_wr[83]));
			radix2 #(.width(width)) rd_st6_68  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[68]), .rdlo_in(a6_wr[84]),  .coef_in(coef[256]), .rdup_out(a7_wr[68]), .rdlo_out(a7_wr[84]));
			radix2 #(.width(width)) rd_st6_69  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[69]), .rdlo_in(a6_wr[85]),  .coef_in(coef[320]), .rdup_out(a7_wr[69]), .rdlo_out(a7_wr[85]));
			radix2 #(.width(width)) rd_st6_70  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[70]), .rdlo_in(a6_wr[86]),  .coef_in(coef[384]), .rdup_out(a7_wr[70]), .rdlo_out(a7_wr[86]));
			radix2 #(.width(width)) rd_st6_71  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[71]), .rdlo_in(a6_wr[87]),  .coef_in(coef[448]), .rdup_out(a7_wr[71]), .rdlo_out(a7_wr[87]));
			radix2 #(.width(width)) rd_st6_72  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[72]), .rdlo_in(a6_wr[88]),  .coef_in(coef[512]), .rdup_out(a7_wr[72]), .rdlo_out(a7_wr[88]));
			radix2 #(.width(width)) rd_st6_73  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[73]), .rdlo_in(a6_wr[89]),  .coef_in(coef[576]), .rdup_out(a7_wr[73]), .rdlo_out(a7_wr[89]));
			radix2 #(.width(width)) rd_st6_74  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[74]), .rdlo_in(a6_wr[90]),  .coef_in(coef[640]), .rdup_out(a7_wr[74]), .rdlo_out(a7_wr[90]));
			radix2 #(.width(width)) rd_st6_75  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[75]), .rdlo_in(a6_wr[91]),  .coef_in(coef[704]), .rdup_out(a7_wr[75]), .rdlo_out(a7_wr[91]));
			radix2 #(.width(width)) rd_st6_76  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[76]), .rdlo_in(a6_wr[92]),  .coef_in(coef[768]), .rdup_out(a7_wr[76]), .rdlo_out(a7_wr[92]));
			radix2 #(.width(width)) rd_st6_77  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[77]), .rdlo_in(a6_wr[93]),  .coef_in(coef[832]), .rdup_out(a7_wr[77]), .rdlo_out(a7_wr[93]));
			radix2 #(.width(width)) rd_st6_78  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[78]), .rdlo_in(a6_wr[94]),  .coef_in(coef[896]), .rdup_out(a7_wr[78]), .rdlo_out(a7_wr[94]));
			radix2 #(.width(width)) rd_st6_79  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[79]), .rdlo_in(a6_wr[95]),  .coef_in(coef[960]), .rdup_out(a7_wr[79]), .rdlo_out(a7_wr[95]));
			radix2 #(.width(width)) rd_st6_96  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[96]), .rdlo_in(a6_wr[112]),  .coef_in(coef[0]), .rdup_out(a7_wr[96]), .rdlo_out(a7_wr[112]));
			radix2 #(.width(width)) rd_st6_97  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[97]), .rdlo_in(a6_wr[113]),  .coef_in(coef[64]), .rdup_out(a7_wr[97]), .rdlo_out(a7_wr[113]));
			radix2 #(.width(width)) rd_st6_98  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[98]), .rdlo_in(a6_wr[114]),  .coef_in(coef[128]), .rdup_out(a7_wr[98]), .rdlo_out(a7_wr[114]));
			radix2 #(.width(width)) rd_st6_99  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[99]), .rdlo_in(a6_wr[115]),  .coef_in(coef[192]), .rdup_out(a7_wr[99]), .rdlo_out(a7_wr[115]));
			radix2 #(.width(width)) rd_st6_100  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[100]), .rdlo_in(a6_wr[116]),  .coef_in(coef[256]), .rdup_out(a7_wr[100]), .rdlo_out(a7_wr[116]));
			radix2 #(.width(width)) rd_st6_101  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[101]), .rdlo_in(a6_wr[117]),  .coef_in(coef[320]), .rdup_out(a7_wr[101]), .rdlo_out(a7_wr[117]));
			radix2 #(.width(width)) rd_st6_102  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[102]), .rdlo_in(a6_wr[118]),  .coef_in(coef[384]), .rdup_out(a7_wr[102]), .rdlo_out(a7_wr[118]));
			radix2 #(.width(width)) rd_st6_103  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[103]), .rdlo_in(a6_wr[119]),  .coef_in(coef[448]), .rdup_out(a7_wr[103]), .rdlo_out(a7_wr[119]));
			radix2 #(.width(width)) rd_st6_104  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[104]), .rdlo_in(a6_wr[120]),  .coef_in(coef[512]), .rdup_out(a7_wr[104]), .rdlo_out(a7_wr[120]));
			radix2 #(.width(width)) rd_st6_105  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[105]), .rdlo_in(a6_wr[121]),  .coef_in(coef[576]), .rdup_out(a7_wr[105]), .rdlo_out(a7_wr[121]));
			radix2 #(.width(width)) rd_st6_106  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[106]), .rdlo_in(a6_wr[122]),  .coef_in(coef[640]), .rdup_out(a7_wr[106]), .rdlo_out(a7_wr[122]));
			radix2 #(.width(width)) rd_st6_107  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[107]), .rdlo_in(a6_wr[123]),  .coef_in(coef[704]), .rdup_out(a7_wr[107]), .rdlo_out(a7_wr[123]));
			radix2 #(.width(width)) rd_st6_108  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[108]), .rdlo_in(a6_wr[124]),  .coef_in(coef[768]), .rdup_out(a7_wr[108]), .rdlo_out(a7_wr[124]));
			radix2 #(.width(width)) rd_st6_109  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[109]), .rdlo_in(a6_wr[125]),  .coef_in(coef[832]), .rdup_out(a7_wr[109]), .rdlo_out(a7_wr[125]));
			radix2 #(.width(width)) rd_st6_110  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[110]), .rdlo_in(a6_wr[126]),  .coef_in(coef[896]), .rdup_out(a7_wr[110]), .rdlo_out(a7_wr[126]));
			radix2 #(.width(width)) rd_st6_111  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[111]), .rdlo_in(a6_wr[127]),  .coef_in(coef[960]), .rdup_out(a7_wr[111]), .rdlo_out(a7_wr[127]));
			radix2 #(.width(width)) rd_st6_128  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[128]), .rdlo_in(a6_wr[144]),  .coef_in(coef[0]), .rdup_out(a7_wr[128]), .rdlo_out(a7_wr[144]));
			radix2 #(.width(width)) rd_st6_129  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[129]), .rdlo_in(a6_wr[145]),  .coef_in(coef[64]), .rdup_out(a7_wr[129]), .rdlo_out(a7_wr[145]));
			radix2 #(.width(width)) rd_st6_130  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[130]), .rdlo_in(a6_wr[146]),  .coef_in(coef[128]), .rdup_out(a7_wr[130]), .rdlo_out(a7_wr[146]));
			radix2 #(.width(width)) rd_st6_131  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[131]), .rdlo_in(a6_wr[147]),  .coef_in(coef[192]), .rdup_out(a7_wr[131]), .rdlo_out(a7_wr[147]));
			radix2 #(.width(width)) rd_st6_132  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[132]), .rdlo_in(a6_wr[148]),  .coef_in(coef[256]), .rdup_out(a7_wr[132]), .rdlo_out(a7_wr[148]));
			radix2 #(.width(width)) rd_st6_133  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[133]), .rdlo_in(a6_wr[149]),  .coef_in(coef[320]), .rdup_out(a7_wr[133]), .rdlo_out(a7_wr[149]));
			radix2 #(.width(width)) rd_st6_134  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[134]), .rdlo_in(a6_wr[150]),  .coef_in(coef[384]), .rdup_out(a7_wr[134]), .rdlo_out(a7_wr[150]));
			radix2 #(.width(width)) rd_st6_135  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[135]), .rdlo_in(a6_wr[151]),  .coef_in(coef[448]), .rdup_out(a7_wr[135]), .rdlo_out(a7_wr[151]));
			radix2 #(.width(width)) rd_st6_136  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[136]), .rdlo_in(a6_wr[152]),  .coef_in(coef[512]), .rdup_out(a7_wr[136]), .rdlo_out(a7_wr[152]));
			radix2 #(.width(width)) rd_st6_137  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[137]), .rdlo_in(a6_wr[153]),  .coef_in(coef[576]), .rdup_out(a7_wr[137]), .rdlo_out(a7_wr[153]));
			radix2 #(.width(width)) rd_st6_138  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[138]), .rdlo_in(a6_wr[154]),  .coef_in(coef[640]), .rdup_out(a7_wr[138]), .rdlo_out(a7_wr[154]));
			radix2 #(.width(width)) rd_st6_139  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[139]), .rdlo_in(a6_wr[155]),  .coef_in(coef[704]), .rdup_out(a7_wr[139]), .rdlo_out(a7_wr[155]));
			radix2 #(.width(width)) rd_st6_140  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[140]), .rdlo_in(a6_wr[156]),  .coef_in(coef[768]), .rdup_out(a7_wr[140]), .rdlo_out(a7_wr[156]));
			radix2 #(.width(width)) rd_st6_141  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[141]), .rdlo_in(a6_wr[157]),  .coef_in(coef[832]), .rdup_out(a7_wr[141]), .rdlo_out(a7_wr[157]));
			radix2 #(.width(width)) rd_st6_142  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[142]), .rdlo_in(a6_wr[158]),  .coef_in(coef[896]), .rdup_out(a7_wr[142]), .rdlo_out(a7_wr[158]));
			radix2 #(.width(width)) rd_st6_143  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[143]), .rdlo_in(a6_wr[159]),  .coef_in(coef[960]), .rdup_out(a7_wr[143]), .rdlo_out(a7_wr[159]));
			radix2 #(.width(width)) rd_st6_160  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[160]), .rdlo_in(a6_wr[176]),  .coef_in(coef[0]), .rdup_out(a7_wr[160]), .rdlo_out(a7_wr[176]));
			radix2 #(.width(width)) rd_st6_161  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[161]), .rdlo_in(a6_wr[177]),  .coef_in(coef[64]), .rdup_out(a7_wr[161]), .rdlo_out(a7_wr[177]));
			radix2 #(.width(width)) rd_st6_162  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[162]), .rdlo_in(a6_wr[178]),  .coef_in(coef[128]), .rdup_out(a7_wr[162]), .rdlo_out(a7_wr[178]));
			radix2 #(.width(width)) rd_st6_163  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[163]), .rdlo_in(a6_wr[179]),  .coef_in(coef[192]), .rdup_out(a7_wr[163]), .rdlo_out(a7_wr[179]));
			radix2 #(.width(width)) rd_st6_164  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[164]), .rdlo_in(a6_wr[180]),  .coef_in(coef[256]), .rdup_out(a7_wr[164]), .rdlo_out(a7_wr[180]));
			radix2 #(.width(width)) rd_st6_165  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[165]), .rdlo_in(a6_wr[181]),  .coef_in(coef[320]), .rdup_out(a7_wr[165]), .rdlo_out(a7_wr[181]));
			radix2 #(.width(width)) rd_st6_166  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[166]), .rdlo_in(a6_wr[182]),  .coef_in(coef[384]), .rdup_out(a7_wr[166]), .rdlo_out(a7_wr[182]));
			radix2 #(.width(width)) rd_st6_167  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[167]), .rdlo_in(a6_wr[183]),  .coef_in(coef[448]), .rdup_out(a7_wr[167]), .rdlo_out(a7_wr[183]));
			radix2 #(.width(width)) rd_st6_168  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[168]), .rdlo_in(a6_wr[184]),  .coef_in(coef[512]), .rdup_out(a7_wr[168]), .rdlo_out(a7_wr[184]));
			radix2 #(.width(width)) rd_st6_169  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[169]), .rdlo_in(a6_wr[185]),  .coef_in(coef[576]), .rdup_out(a7_wr[169]), .rdlo_out(a7_wr[185]));
			radix2 #(.width(width)) rd_st6_170  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[170]), .rdlo_in(a6_wr[186]),  .coef_in(coef[640]), .rdup_out(a7_wr[170]), .rdlo_out(a7_wr[186]));
			radix2 #(.width(width)) rd_st6_171  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[171]), .rdlo_in(a6_wr[187]),  .coef_in(coef[704]), .rdup_out(a7_wr[171]), .rdlo_out(a7_wr[187]));
			radix2 #(.width(width)) rd_st6_172  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[172]), .rdlo_in(a6_wr[188]),  .coef_in(coef[768]), .rdup_out(a7_wr[172]), .rdlo_out(a7_wr[188]));
			radix2 #(.width(width)) rd_st6_173  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[173]), .rdlo_in(a6_wr[189]),  .coef_in(coef[832]), .rdup_out(a7_wr[173]), .rdlo_out(a7_wr[189]));
			radix2 #(.width(width)) rd_st6_174  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[174]), .rdlo_in(a6_wr[190]),  .coef_in(coef[896]), .rdup_out(a7_wr[174]), .rdlo_out(a7_wr[190]));
			radix2 #(.width(width)) rd_st6_175  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[175]), .rdlo_in(a6_wr[191]),  .coef_in(coef[960]), .rdup_out(a7_wr[175]), .rdlo_out(a7_wr[191]));
			radix2 #(.width(width)) rd_st6_192  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[192]), .rdlo_in(a6_wr[208]),  .coef_in(coef[0]), .rdup_out(a7_wr[192]), .rdlo_out(a7_wr[208]));
			radix2 #(.width(width)) rd_st6_193  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[193]), .rdlo_in(a6_wr[209]),  .coef_in(coef[64]), .rdup_out(a7_wr[193]), .rdlo_out(a7_wr[209]));
			radix2 #(.width(width)) rd_st6_194  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[194]), .rdlo_in(a6_wr[210]),  .coef_in(coef[128]), .rdup_out(a7_wr[194]), .rdlo_out(a7_wr[210]));
			radix2 #(.width(width)) rd_st6_195  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[195]), .rdlo_in(a6_wr[211]),  .coef_in(coef[192]), .rdup_out(a7_wr[195]), .rdlo_out(a7_wr[211]));
			radix2 #(.width(width)) rd_st6_196  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[196]), .rdlo_in(a6_wr[212]),  .coef_in(coef[256]), .rdup_out(a7_wr[196]), .rdlo_out(a7_wr[212]));
			radix2 #(.width(width)) rd_st6_197  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[197]), .rdlo_in(a6_wr[213]),  .coef_in(coef[320]), .rdup_out(a7_wr[197]), .rdlo_out(a7_wr[213]));
			radix2 #(.width(width)) rd_st6_198  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[198]), .rdlo_in(a6_wr[214]),  .coef_in(coef[384]), .rdup_out(a7_wr[198]), .rdlo_out(a7_wr[214]));
			radix2 #(.width(width)) rd_st6_199  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[199]), .rdlo_in(a6_wr[215]),  .coef_in(coef[448]), .rdup_out(a7_wr[199]), .rdlo_out(a7_wr[215]));
			radix2 #(.width(width)) rd_st6_200  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[200]), .rdlo_in(a6_wr[216]),  .coef_in(coef[512]), .rdup_out(a7_wr[200]), .rdlo_out(a7_wr[216]));
			radix2 #(.width(width)) rd_st6_201  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[201]), .rdlo_in(a6_wr[217]),  .coef_in(coef[576]), .rdup_out(a7_wr[201]), .rdlo_out(a7_wr[217]));
			radix2 #(.width(width)) rd_st6_202  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[202]), .rdlo_in(a6_wr[218]),  .coef_in(coef[640]), .rdup_out(a7_wr[202]), .rdlo_out(a7_wr[218]));
			radix2 #(.width(width)) rd_st6_203  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[203]), .rdlo_in(a6_wr[219]),  .coef_in(coef[704]), .rdup_out(a7_wr[203]), .rdlo_out(a7_wr[219]));
			radix2 #(.width(width)) rd_st6_204  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[204]), .rdlo_in(a6_wr[220]),  .coef_in(coef[768]), .rdup_out(a7_wr[204]), .rdlo_out(a7_wr[220]));
			radix2 #(.width(width)) rd_st6_205  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[205]), .rdlo_in(a6_wr[221]),  .coef_in(coef[832]), .rdup_out(a7_wr[205]), .rdlo_out(a7_wr[221]));
			radix2 #(.width(width)) rd_st6_206  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[206]), .rdlo_in(a6_wr[222]),  .coef_in(coef[896]), .rdup_out(a7_wr[206]), .rdlo_out(a7_wr[222]));
			radix2 #(.width(width)) rd_st6_207  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[207]), .rdlo_in(a6_wr[223]),  .coef_in(coef[960]), .rdup_out(a7_wr[207]), .rdlo_out(a7_wr[223]));
			radix2 #(.width(width)) rd_st6_224  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[224]), .rdlo_in(a6_wr[240]),  .coef_in(coef[0]), .rdup_out(a7_wr[224]), .rdlo_out(a7_wr[240]));
			radix2 #(.width(width)) rd_st6_225  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[225]), .rdlo_in(a6_wr[241]),  .coef_in(coef[64]), .rdup_out(a7_wr[225]), .rdlo_out(a7_wr[241]));
			radix2 #(.width(width)) rd_st6_226  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[226]), .rdlo_in(a6_wr[242]),  .coef_in(coef[128]), .rdup_out(a7_wr[226]), .rdlo_out(a7_wr[242]));
			radix2 #(.width(width)) rd_st6_227  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[227]), .rdlo_in(a6_wr[243]),  .coef_in(coef[192]), .rdup_out(a7_wr[227]), .rdlo_out(a7_wr[243]));
			radix2 #(.width(width)) rd_st6_228  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[228]), .rdlo_in(a6_wr[244]),  .coef_in(coef[256]), .rdup_out(a7_wr[228]), .rdlo_out(a7_wr[244]));
			radix2 #(.width(width)) rd_st6_229  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[229]), .rdlo_in(a6_wr[245]),  .coef_in(coef[320]), .rdup_out(a7_wr[229]), .rdlo_out(a7_wr[245]));
			radix2 #(.width(width)) rd_st6_230  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[230]), .rdlo_in(a6_wr[246]),  .coef_in(coef[384]), .rdup_out(a7_wr[230]), .rdlo_out(a7_wr[246]));
			radix2 #(.width(width)) rd_st6_231  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[231]), .rdlo_in(a6_wr[247]),  .coef_in(coef[448]), .rdup_out(a7_wr[231]), .rdlo_out(a7_wr[247]));
			radix2 #(.width(width)) rd_st6_232  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[232]), .rdlo_in(a6_wr[248]),  .coef_in(coef[512]), .rdup_out(a7_wr[232]), .rdlo_out(a7_wr[248]));
			radix2 #(.width(width)) rd_st6_233  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[233]), .rdlo_in(a6_wr[249]),  .coef_in(coef[576]), .rdup_out(a7_wr[233]), .rdlo_out(a7_wr[249]));
			radix2 #(.width(width)) rd_st6_234  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[234]), .rdlo_in(a6_wr[250]),  .coef_in(coef[640]), .rdup_out(a7_wr[234]), .rdlo_out(a7_wr[250]));
			radix2 #(.width(width)) rd_st6_235  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[235]), .rdlo_in(a6_wr[251]),  .coef_in(coef[704]), .rdup_out(a7_wr[235]), .rdlo_out(a7_wr[251]));
			radix2 #(.width(width)) rd_st6_236  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[236]), .rdlo_in(a6_wr[252]),  .coef_in(coef[768]), .rdup_out(a7_wr[236]), .rdlo_out(a7_wr[252]));
			radix2 #(.width(width)) rd_st6_237  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[237]), .rdlo_in(a6_wr[253]),  .coef_in(coef[832]), .rdup_out(a7_wr[237]), .rdlo_out(a7_wr[253]));
			radix2 #(.width(width)) rd_st6_238  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[238]), .rdlo_in(a6_wr[254]),  .coef_in(coef[896]), .rdup_out(a7_wr[238]), .rdlo_out(a7_wr[254]));
			radix2 #(.width(width)) rd_st6_239  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[239]), .rdlo_in(a6_wr[255]),  .coef_in(coef[960]), .rdup_out(a7_wr[239]), .rdlo_out(a7_wr[255]));
			radix2 #(.width(width)) rd_st6_256  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[256]), .rdlo_in(a6_wr[272]),  .coef_in(coef[0]), .rdup_out(a7_wr[256]), .rdlo_out(a7_wr[272]));
			radix2 #(.width(width)) rd_st6_257  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[257]), .rdlo_in(a6_wr[273]),  .coef_in(coef[64]), .rdup_out(a7_wr[257]), .rdlo_out(a7_wr[273]));
			radix2 #(.width(width)) rd_st6_258  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[258]), .rdlo_in(a6_wr[274]),  .coef_in(coef[128]), .rdup_out(a7_wr[258]), .rdlo_out(a7_wr[274]));
			radix2 #(.width(width)) rd_st6_259  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[259]), .rdlo_in(a6_wr[275]),  .coef_in(coef[192]), .rdup_out(a7_wr[259]), .rdlo_out(a7_wr[275]));
			radix2 #(.width(width)) rd_st6_260  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[260]), .rdlo_in(a6_wr[276]),  .coef_in(coef[256]), .rdup_out(a7_wr[260]), .rdlo_out(a7_wr[276]));
			radix2 #(.width(width)) rd_st6_261  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[261]), .rdlo_in(a6_wr[277]),  .coef_in(coef[320]), .rdup_out(a7_wr[261]), .rdlo_out(a7_wr[277]));
			radix2 #(.width(width)) rd_st6_262  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[262]), .rdlo_in(a6_wr[278]),  .coef_in(coef[384]), .rdup_out(a7_wr[262]), .rdlo_out(a7_wr[278]));
			radix2 #(.width(width)) rd_st6_263  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[263]), .rdlo_in(a6_wr[279]),  .coef_in(coef[448]), .rdup_out(a7_wr[263]), .rdlo_out(a7_wr[279]));
			radix2 #(.width(width)) rd_st6_264  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[264]), .rdlo_in(a6_wr[280]),  .coef_in(coef[512]), .rdup_out(a7_wr[264]), .rdlo_out(a7_wr[280]));
			radix2 #(.width(width)) rd_st6_265  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[265]), .rdlo_in(a6_wr[281]),  .coef_in(coef[576]), .rdup_out(a7_wr[265]), .rdlo_out(a7_wr[281]));
			radix2 #(.width(width)) rd_st6_266  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[266]), .rdlo_in(a6_wr[282]),  .coef_in(coef[640]), .rdup_out(a7_wr[266]), .rdlo_out(a7_wr[282]));
			radix2 #(.width(width)) rd_st6_267  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[267]), .rdlo_in(a6_wr[283]),  .coef_in(coef[704]), .rdup_out(a7_wr[267]), .rdlo_out(a7_wr[283]));
			radix2 #(.width(width)) rd_st6_268  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[268]), .rdlo_in(a6_wr[284]),  .coef_in(coef[768]), .rdup_out(a7_wr[268]), .rdlo_out(a7_wr[284]));
			radix2 #(.width(width)) rd_st6_269  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[269]), .rdlo_in(a6_wr[285]),  .coef_in(coef[832]), .rdup_out(a7_wr[269]), .rdlo_out(a7_wr[285]));
			radix2 #(.width(width)) rd_st6_270  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[270]), .rdlo_in(a6_wr[286]),  .coef_in(coef[896]), .rdup_out(a7_wr[270]), .rdlo_out(a7_wr[286]));
			radix2 #(.width(width)) rd_st6_271  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[271]), .rdlo_in(a6_wr[287]),  .coef_in(coef[960]), .rdup_out(a7_wr[271]), .rdlo_out(a7_wr[287]));
			radix2 #(.width(width)) rd_st6_288  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[288]), .rdlo_in(a6_wr[304]),  .coef_in(coef[0]), .rdup_out(a7_wr[288]), .rdlo_out(a7_wr[304]));
			radix2 #(.width(width)) rd_st6_289  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[289]), .rdlo_in(a6_wr[305]),  .coef_in(coef[64]), .rdup_out(a7_wr[289]), .rdlo_out(a7_wr[305]));
			radix2 #(.width(width)) rd_st6_290  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[290]), .rdlo_in(a6_wr[306]),  .coef_in(coef[128]), .rdup_out(a7_wr[290]), .rdlo_out(a7_wr[306]));
			radix2 #(.width(width)) rd_st6_291  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[291]), .rdlo_in(a6_wr[307]),  .coef_in(coef[192]), .rdup_out(a7_wr[291]), .rdlo_out(a7_wr[307]));
			radix2 #(.width(width)) rd_st6_292  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[292]), .rdlo_in(a6_wr[308]),  .coef_in(coef[256]), .rdup_out(a7_wr[292]), .rdlo_out(a7_wr[308]));
			radix2 #(.width(width)) rd_st6_293  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[293]), .rdlo_in(a6_wr[309]),  .coef_in(coef[320]), .rdup_out(a7_wr[293]), .rdlo_out(a7_wr[309]));
			radix2 #(.width(width)) rd_st6_294  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[294]), .rdlo_in(a6_wr[310]),  .coef_in(coef[384]), .rdup_out(a7_wr[294]), .rdlo_out(a7_wr[310]));
			radix2 #(.width(width)) rd_st6_295  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[295]), .rdlo_in(a6_wr[311]),  .coef_in(coef[448]), .rdup_out(a7_wr[295]), .rdlo_out(a7_wr[311]));
			radix2 #(.width(width)) rd_st6_296  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[296]), .rdlo_in(a6_wr[312]),  .coef_in(coef[512]), .rdup_out(a7_wr[296]), .rdlo_out(a7_wr[312]));
			radix2 #(.width(width)) rd_st6_297  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[297]), .rdlo_in(a6_wr[313]),  .coef_in(coef[576]), .rdup_out(a7_wr[297]), .rdlo_out(a7_wr[313]));
			radix2 #(.width(width)) rd_st6_298  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[298]), .rdlo_in(a6_wr[314]),  .coef_in(coef[640]), .rdup_out(a7_wr[298]), .rdlo_out(a7_wr[314]));
			radix2 #(.width(width)) rd_st6_299  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[299]), .rdlo_in(a6_wr[315]),  .coef_in(coef[704]), .rdup_out(a7_wr[299]), .rdlo_out(a7_wr[315]));
			radix2 #(.width(width)) rd_st6_300  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[300]), .rdlo_in(a6_wr[316]),  .coef_in(coef[768]), .rdup_out(a7_wr[300]), .rdlo_out(a7_wr[316]));
			radix2 #(.width(width)) rd_st6_301  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[301]), .rdlo_in(a6_wr[317]),  .coef_in(coef[832]), .rdup_out(a7_wr[301]), .rdlo_out(a7_wr[317]));
			radix2 #(.width(width)) rd_st6_302  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[302]), .rdlo_in(a6_wr[318]),  .coef_in(coef[896]), .rdup_out(a7_wr[302]), .rdlo_out(a7_wr[318]));
			radix2 #(.width(width)) rd_st6_303  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[303]), .rdlo_in(a6_wr[319]),  .coef_in(coef[960]), .rdup_out(a7_wr[303]), .rdlo_out(a7_wr[319]));
			radix2 #(.width(width)) rd_st6_320  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[320]), .rdlo_in(a6_wr[336]),  .coef_in(coef[0]), .rdup_out(a7_wr[320]), .rdlo_out(a7_wr[336]));
			radix2 #(.width(width)) rd_st6_321  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[321]), .rdlo_in(a6_wr[337]),  .coef_in(coef[64]), .rdup_out(a7_wr[321]), .rdlo_out(a7_wr[337]));
			radix2 #(.width(width)) rd_st6_322  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[322]), .rdlo_in(a6_wr[338]),  .coef_in(coef[128]), .rdup_out(a7_wr[322]), .rdlo_out(a7_wr[338]));
			radix2 #(.width(width)) rd_st6_323  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[323]), .rdlo_in(a6_wr[339]),  .coef_in(coef[192]), .rdup_out(a7_wr[323]), .rdlo_out(a7_wr[339]));
			radix2 #(.width(width)) rd_st6_324  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[324]), .rdlo_in(a6_wr[340]),  .coef_in(coef[256]), .rdup_out(a7_wr[324]), .rdlo_out(a7_wr[340]));
			radix2 #(.width(width)) rd_st6_325  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[325]), .rdlo_in(a6_wr[341]),  .coef_in(coef[320]), .rdup_out(a7_wr[325]), .rdlo_out(a7_wr[341]));
			radix2 #(.width(width)) rd_st6_326  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[326]), .rdlo_in(a6_wr[342]),  .coef_in(coef[384]), .rdup_out(a7_wr[326]), .rdlo_out(a7_wr[342]));
			radix2 #(.width(width)) rd_st6_327  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[327]), .rdlo_in(a6_wr[343]),  .coef_in(coef[448]), .rdup_out(a7_wr[327]), .rdlo_out(a7_wr[343]));
			radix2 #(.width(width)) rd_st6_328  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[328]), .rdlo_in(a6_wr[344]),  .coef_in(coef[512]), .rdup_out(a7_wr[328]), .rdlo_out(a7_wr[344]));
			radix2 #(.width(width)) rd_st6_329  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[329]), .rdlo_in(a6_wr[345]),  .coef_in(coef[576]), .rdup_out(a7_wr[329]), .rdlo_out(a7_wr[345]));
			radix2 #(.width(width)) rd_st6_330  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[330]), .rdlo_in(a6_wr[346]),  .coef_in(coef[640]), .rdup_out(a7_wr[330]), .rdlo_out(a7_wr[346]));
			radix2 #(.width(width)) rd_st6_331  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[331]), .rdlo_in(a6_wr[347]),  .coef_in(coef[704]), .rdup_out(a7_wr[331]), .rdlo_out(a7_wr[347]));
			radix2 #(.width(width)) rd_st6_332  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[332]), .rdlo_in(a6_wr[348]),  .coef_in(coef[768]), .rdup_out(a7_wr[332]), .rdlo_out(a7_wr[348]));
			radix2 #(.width(width)) rd_st6_333  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[333]), .rdlo_in(a6_wr[349]),  .coef_in(coef[832]), .rdup_out(a7_wr[333]), .rdlo_out(a7_wr[349]));
			radix2 #(.width(width)) rd_st6_334  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[334]), .rdlo_in(a6_wr[350]),  .coef_in(coef[896]), .rdup_out(a7_wr[334]), .rdlo_out(a7_wr[350]));
			radix2 #(.width(width)) rd_st6_335  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[335]), .rdlo_in(a6_wr[351]),  .coef_in(coef[960]), .rdup_out(a7_wr[335]), .rdlo_out(a7_wr[351]));
			radix2 #(.width(width)) rd_st6_352  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[352]), .rdlo_in(a6_wr[368]),  .coef_in(coef[0]), .rdup_out(a7_wr[352]), .rdlo_out(a7_wr[368]));
			radix2 #(.width(width)) rd_st6_353  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[353]), .rdlo_in(a6_wr[369]),  .coef_in(coef[64]), .rdup_out(a7_wr[353]), .rdlo_out(a7_wr[369]));
			radix2 #(.width(width)) rd_st6_354  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[354]), .rdlo_in(a6_wr[370]),  .coef_in(coef[128]), .rdup_out(a7_wr[354]), .rdlo_out(a7_wr[370]));
			radix2 #(.width(width)) rd_st6_355  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[355]), .rdlo_in(a6_wr[371]),  .coef_in(coef[192]), .rdup_out(a7_wr[355]), .rdlo_out(a7_wr[371]));
			radix2 #(.width(width)) rd_st6_356  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[356]), .rdlo_in(a6_wr[372]),  .coef_in(coef[256]), .rdup_out(a7_wr[356]), .rdlo_out(a7_wr[372]));
			radix2 #(.width(width)) rd_st6_357  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[357]), .rdlo_in(a6_wr[373]),  .coef_in(coef[320]), .rdup_out(a7_wr[357]), .rdlo_out(a7_wr[373]));
			radix2 #(.width(width)) rd_st6_358  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[358]), .rdlo_in(a6_wr[374]),  .coef_in(coef[384]), .rdup_out(a7_wr[358]), .rdlo_out(a7_wr[374]));
			radix2 #(.width(width)) rd_st6_359  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[359]), .rdlo_in(a6_wr[375]),  .coef_in(coef[448]), .rdup_out(a7_wr[359]), .rdlo_out(a7_wr[375]));
			radix2 #(.width(width)) rd_st6_360  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[360]), .rdlo_in(a6_wr[376]),  .coef_in(coef[512]), .rdup_out(a7_wr[360]), .rdlo_out(a7_wr[376]));
			radix2 #(.width(width)) rd_st6_361  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[361]), .rdlo_in(a6_wr[377]),  .coef_in(coef[576]), .rdup_out(a7_wr[361]), .rdlo_out(a7_wr[377]));
			radix2 #(.width(width)) rd_st6_362  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[362]), .rdlo_in(a6_wr[378]),  .coef_in(coef[640]), .rdup_out(a7_wr[362]), .rdlo_out(a7_wr[378]));
			radix2 #(.width(width)) rd_st6_363  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[363]), .rdlo_in(a6_wr[379]),  .coef_in(coef[704]), .rdup_out(a7_wr[363]), .rdlo_out(a7_wr[379]));
			radix2 #(.width(width)) rd_st6_364  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[364]), .rdlo_in(a6_wr[380]),  .coef_in(coef[768]), .rdup_out(a7_wr[364]), .rdlo_out(a7_wr[380]));
			radix2 #(.width(width)) rd_st6_365  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[365]), .rdlo_in(a6_wr[381]),  .coef_in(coef[832]), .rdup_out(a7_wr[365]), .rdlo_out(a7_wr[381]));
			radix2 #(.width(width)) rd_st6_366  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[366]), .rdlo_in(a6_wr[382]),  .coef_in(coef[896]), .rdup_out(a7_wr[366]), .rdlo_out(a7_wr[382]));
			radix2 #(.width(width)) rd_st6_367  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[367]), .rdlo_in(a6_wr[383]),  .coef_in(coef[960]), .rdup_out(a7_wr[367]), .rdlo_out(a7_wr[383]));
			radix2 #(.width(width)) rd_st6_384  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[384]), .rdlo_in(a6_wr[400]),  .coef_in(coef[0]), .rdup_out(a7_wr[384]), .rdlo_out(a7_wr[400]));
			radix2 #(.width(width)) rd_st6_385  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[385]), .rdlo_in(a6_wr[401]),  .coef_in(coef[64]), .rdup_out(a7_wr[385]), .rdlo_out(a7_wr[401]));
			radix2 #(.width(width)) rd_st6_386  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[386]), .rdlo_in(a6_wr[402]),  .coef_in(coef[128]), .rdup_out(a7_wr[386]), .rdlo_out(a7_wr[402]));
			radix2 #(.width(width)) rd_st6_387  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[387]), .rdlo_in(a6_wr[403]),  .coef_in(coef[192]), .rdup_out(a7_wr[387]), .rdlo_out(a7_wr[403]));
			radix2 #(.width(width)) rd_st6_388  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[388]), .rdlo_in(a6_wr[404]),  .coef_in(coef[256]), .rdup_out(a7_wr[388]), .rdlo_out(a7_wr[404]));
			radix2 #(.width(width)) rd_st6_389  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[389]), .rdlo_in(a6_wr[405]),  .coef_in(coef[320]), .rdup_out(a7_wr[389]), .rdlo_out(a7_wr[405]));
			radix2 #(.width(width)) rd_st6_390  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[390]), .rdlo_in(a6_wr[406]),  .coef_in(coef[384]), .rdup_out(a7_wr[390]), .rdlo_out(a7_wr[406]));
			radix2 #(.width(width)) rd_st6_391  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[391]), .rdlo_in(a6_wr[407]),  .coef_in(coef[448]), .rdup_out(a7_wr[391]), .rdlo_out(a7_wr[407]));
			radix2 #(.width(width)) rd_st6_392  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[392]), .rdlo_in(a6_wr[408]),  .coef_in(coef[512]), .rdup_out(a7_wr[392]), .rdlo_out(a7_wr[408]));
			radix2 #(.width(width)) rd_st6_393  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[393]), .rdlo_in(a6_wr[409]),  .coef_in(coef[576]), .rdup_out(a7_wr[393]), .rdlo_out(a7_wr[409]));
			radix2 #(.width(width)) rd_st6_394  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[394]), .rdlo_in(a6_wr[410]),  .coef_in(coef[640]), .rdup_out(a7_wr[394]), .rdlo_out(a7_wr[410]));
			radix2 #(.width(width)) rd_st6_395  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[395]), .rdlo_in(a6_wr[411]),  .coef_in(coef[704]), .rdup_out(a7_wr[395]), .rdlo_out(a7_wr[411]));
			radix2 #(.width(width)) rd_st6_396  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[396]), .rdlo_in(a6_wr[412]),  .coef_in(coef[768]), .rdup_out(a7_wr[396]), .rdlo_out(a7_wr[412]));
			radix2 #(.width(width)) rd_st6_397  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[397]), .rdlo_in(a6_wr[413]),  .coef_in(coef[832]), .rdup_out(a7_wr[397]), .rdlo_out(a7_wr[413]));
			radix2 #(.width(width)) rd_st6_398  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[398]), .rdlo_in(a6_wr[414]),  .coef_in(coef[896]), .rdup_out(a7_wr[398]), .rdlo_out(a7_wr[414]));
			radix2 #(.width(width)) rd_st6_399  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[399]), .rdlo_in(a6_wr[415]),  .coef_in(coef[960]), .rdup_out(a7_wr[399]), .rdlo_out(a7_wr[415]));
			radix2 #(.width(width)) rd_st6_416  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[416]), .rdlo_in(a6_wr[432]),  .coef_in(coef[0]), .rdup_out(a7_wr[416]), .rdlo_out(a7_wr[432]));
			radix2 #(.width(width)) rd_st6_417  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[417]), .rdlo_in(a6_wr[433]),  .coef_in(coef[64]), .rdup_out(a7_wr[417]), .rdlo_out(a7_wr[433]));
			radix2 #(.width(width)) rd_st6_418  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[418]), .rdlo_in(a6_wr[434]),  .coef_in(coef[128]), .rdup_out(a7_wr[418]), .rdlo_out(a7_wr[434]));
			radix2 #(.width(width)) rd_st6_419  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[419]), .rdlo_in(a6_wr[435]),  .coef_in(coef[192]), .rdup_out(a7_wr[419]), .rdlo_out(a7_wr[435]));
			radix2 #(.width(width)) rd_st6_420  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[420]), .rdlo_in(a6_wr[436]),  .coef_in(coef[256]), .rdup_out(a7_wr[420]), .rdlo_out(a7_wr[436]));
			radix2 #(.width(width)) rd_st6_421  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[421]), .rdlo_in(a6_wr[437]),  .coef_in(coef[320]), .rdup_out(a7_wr[421]), .rdlo_out(a7_wr[437]));
			radix2 #(.width(width)) rd_st6_422  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[422]), .rdlo_in(a6_wr[438]),  .coef_in(coef[384]), .rdup_out(a7_wr[422]), .rdlo_out(a7_wr[438]));
			radix2 #(.width(width)) rd_st6_423  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[423]), .rdlo_in(a6_wr[439]),  .coef_in(coef[448]), .rdup_out(a7_wr[423]), .rdlo_out(a7_wr[439]));
			radix2 #(.width(width)) rd_st6_424  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[424]), .rdlo_in(a6_wr[440]),  .coef_in(coef[512]), .rdup_out(a7_wr[424]), .rdlo_out(a7_wr[440]));
			radix2 #(.width(width)) rd_st6_425  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[425]), .rdlo_in(a6_wr[441]),  .coef_in(coef[576]), .rdup_out(a7_wr[425]), .rdlo_out(a7_wr[441]));
			radix2 #(.width(width)) rd_st6_426  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[426]), .rdlo_in(a6_wr[442]),  .coef_in(coef[640]), .rdup_out(a7_wr[426]), .rdlo_out(a7_wr[442]));
			radix2 #(.width(width)) rd_st6_427  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[427]), .rdlo_in(a6_wr[443]),  .coef_in(coef[704]), .rdup_out(a7_wr[427]), .rdlo_out(a7_wr[443]));
			radix2 #(.width(width)) rd_st6_428  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[428]), .rdlo_in(a6_wr[444]),  .coef_in(coef[768]), .rdup_out(a7_wr[428]), .rdlo_out(a7_wr[444]));
			radix2 #(.width(width)) rd_st6_429  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[429]), .rdlo_in(a6_wr[445]),  .coef_in(coef[832]), .rdup_out(a7_wr[429]), .rdlo_out(a7_wr[445]));
			radix2 #(.width(width)) rd_st6_430  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[430]), .rdlo_in(a6_wr[446]),  .coef_in(coef[896]), .rdup_out(a7_wr[430]), .rdlo_out(a7_wr[446]));
			radix2 #(.width(width)) rd_st6_431  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[431]), .rdlo_in(a6_wr[447]),  .coef_in(coef[960]), .rdup_out(a7_wr[431]), .rdlo_out(a7_wr[447]));
			radix2 #(.width(width)) rd_st6_448  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[448]), .rdlo_in(a6_wr[464]),  .coef_in(coef[0]), .rdup_out(a7_wr[448]), .rdlo_out(a7_wr[464]));
			radix2 #(.width(width)) rd_st6_449  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[449]), .rdlo_in(a6_wr[465]),  .coef_in(coef[64]), .rdup_out(a7_wr[449]), .rdlo_out(a7_wr[465]));
			radix2 #(.width(width)) rd_st6_450  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[450]), .rdlo_in(a6_wr[466]),  .coef_in(coef[128]), .rdup_out(a7_wr[450]), .rdlo_out(a7_wr[466]));
			radix2 #(.width(width)) rd_st6_451  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[451]), .rdlo_in(a6_wr[467]),  .coef_in(coef[192]), .rdup_out(a7_wr[451]), .rdlo_out(a7_wr[467]));
			radix2 #(.width(width)) rd_st6_452  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[452]), .rdlo_in(a6_wr[468]),  .coef_in(coef[256]), .rdup_out(a7_wr[452]), .rdlo_out(a7_wr[468]));
			radix2 #(.width(width)) rd_st6_453  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[453]), .rdlo_in(a6_wr[469]),  .coef_in(coef[320]), .rdup_out(a7_wr[453]), .rdlo_out(a7_wr[469]));
			radix2 #(.width(width)) rd_st6_454  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[454]), .rdlo_in(a6_wr[470]),  .coef_in(coef[384]), .rdup_out(a7_wr[454]), .rdlo_out(a7_wr[470]));
			radix2 #(.width(width)) rd_st6_455  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[455]), .rdlo_in(a6_wr[471]),  .coef_in(coef[448]), .rdup_out(a7_wr[455]), .rdlo_out(a7_wr[471]));
			radix2 #(.width(width)) rd_st6_456  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[456]), .rdlo_in(a6_wr[472]),  .coef_in(coef[512]), .rdup_out(a7_wr[456]), .rdlo_out(a7_wr[472]));
			radix2 #(.width(width)) rd_st6_457  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[457]), .rdlo_in(a6_wr[473]),  .coef_in(coef[576]), .rdup_out(a7_wr[457]), .rdlo_out(a7_wr[473]));
			radix2 #(.width(width)) rd_st6_458  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[458]), .rdlo_in(a6_wr[474]),  .coef_in(coef[640]), .rdup_out(a7_wr[458]), .rdlo_out(a7_wr[474]));
			radix2 #(.width(width)) rd_st6_459  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[459]), .rdlo_in(a6_wr[475]),  .coef_in(coef[704]), .rdup_out(a7_wr[459]), .rdlo_out(a7_wr[475]));
			radix2 #(.width(width)) rd_st6_460  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[460]), .rdlo_in(a6_wr[476]),  .coef_in(coef[768]), .rdup_out(a7_wr[460]), .rdlo_out(a7_wr[476]));
			radix2 #(.width(width)) rd_st6_461  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[461]), .rdlo_in(a6_wr[477]),  .coef_in(coef[832]), .rdup_out(a7_wr[461]), .rdlo_out(a7_wr[477]));
			radix2 #(.width(width)) rd_st6_462  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[462]), .rdlo_in(a6_wr[478]),  .coef_in(coef[896]), .rdup_out(a7_wr[462]), .rdlo_out(a7_wr[478]));
			radix2 #(.width(width)) rd_st6_463  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[463]), .rdlo_in(a6_wr[479]),  .coef_in(coef[960]), .rdup_out(a7_wr[463]), .rdlo_out(a7_wr[479]));
			radix2 #(.width(width)) rd_st6_480  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[480]), .rdlo_in(a6_wr[496]),  .coef_in(coef[0]), .rdup_out(a7_wr[480]), .rdlo_out(a7_wr[496]));
			radix2 #(.width(width)) rd_st6_481  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[481]), .rdlo_in(a6_wr[497]),  .coef_in(coef[64]), .rdup_out(a7_wr[481]), .rdlo_out(a7_wr[497]));
			radix2 #(.width(width)) rd_st6_482  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[482]), .rdlo_in(a6_wr[498]),  .coef_in(coef[128]), .rdup_out(a7_wr[482]), .rdlo_out(a7_wr[498]));
			radix2 #(.width(width)) rd_st6_483  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[483]), .rdlo_in(a6_wr[499]),  .coef_in(coef[192]), .rdup_out(a7_wr[483]), .rdlo_out(a7_wr[499]));
			radix2 #(.width(width)) rd_st6_484  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[484]), .rdlo_in(a6_wr[500]),  .coef_in(coef[256]), .rdup_out(a7_wr[484]), .rdlo_out(a7_wr[500]));
			radix2 #(.width(width)) rd_st6_485  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[485]), .rdlo_in(a6_wr[501]),  .coef_in(coef[320]), .rdup_out(a7_wr[485]), .rdlo_out(a7_wr[501]));
			radix2 #(.width(width)) rd_st6_486  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[486]), .rdlo_in(a6_wr[502]),  .coef_in(coef[384]), .rdup_out(a7_wr[486]), .rdlo_out(a7_wr[502]));
			radix2 #(.width(width)) rd_st6_487  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[487]), .rdlo_in(a6_wr[503]),  .coef_in(coef[448]), .rdup_out(a7_wr[487]), .rdlo_out(a7_wr[503]));
			radix2 #(.width(width)) rd_st6_488  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[488]), .rdlo_in(a6_wr[504]),  .coef_in(coef[512]), .rdup_out(a7_wr[488]), .rdlo_out(a7_wr[504]));
			radix2 #(.width(width)) rd_st6_489  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[489]), .rdlo_in(a6_wr[505]),  .coef_in(coef[576]), .rdup_out(a7_wr[489]), .rdlo_out(a7_wr[505]));
			radix2 #(.width(width)) rd_st6_490  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[490]), .rdlo_in(a6_wr[506]),  .coef_in(coef[640]), .rdup_out(a7_wr[490]), .rdlo_out(a7_wr[506]));
			radix2 #(.width(width)) rd_st6_491  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[491]), .rdlo_in(a6_wr[507]),  .coef_in(coef[704]), .rdup_out(a7_wr[491]), .rdlo_out(a7_wr[507]));
			radix2 #(.width(width)) rd_st6_492  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[492]), .rdlo_in(a6_wr[508]),  .coef_in(coef[768]), .rdup_out(a7_wr[492]), .rdlo_out(a7_wr[508]));
			radix2 #(.width(width)) rd_st6_493  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[493]), .rdlo_in(a6_wr[509]),  .coef_in(coef[832]), .rdup_out(a7_wr[493]), .rdlo_out(a7_wr[509]));
			radix2 #(.width(width)) rd_st6_494  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[494]), .rdlo_in(a6_wr[510]),  .coef_in(coef[896]), .rdup_out(a7_wr[494]), .rdlo_out(a7_wr[510]));
			radix2 #(.width(width)) rd_st6_495  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[495]), .rdlo_in(a6_wr[511]),  .coef_in(coef[960]), .rdup_out(a7_wr[495]), .rdlo_out(a7_wr[511]));
			radix2 #(.width(width)) rd_st6_512  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[512]), .rdlo_in(a6_wr[528]),  .coef_in(coef[0]), .rdup_out(a7_wr[512]), .rdlo_out(a7_wr[528]));
			radix2 #(.width(width)) rd_st6_513  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[513]), .rdlo_in(a6_wr[529]),  .coef_in(coef[64]), .rdup_out(a7_wr[513]), .rdlo_out(a7_wr[529]));
			radix2 #(.width(width)) rd_st6_514  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[514]), .rdlo_in(a6_wr[530]),  .coef_in(coef[128]), .rdup_out(a7_wr[514]), .rdlo_out(a7_wr[530]));
			radix2 #(.width(width)) rd_st6_515  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[515]), .rdlo_in(a6_wr[531]),  .coef_in(coef[192]), .rdup_out(a7_wr[515]), .rdlo_out(a7_wr[531]));
			radix2 #(.width(width)) rd_st6_516  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[516]), .rdlo_in(a6_wr[532]),  .coef_in(coef[256]), .rdup_out(a7_wr[516]), .rdlo_out(a7_wr[532]));
			radix2 #(.width(width)) rd_st6_517  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[517]), .rdlo_in(a6_wr[533]),  .coef_in(coef[320]), .rdup_out(a7_wr[517]), .rdlo_out(a7_wr[533]));
			radix2 #(.width(width)) rd_st6_518  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[518]), .rdlo_in(a6_wr[534]),  .coef_in(coef[384]), .rdup_out(a7_wr[518]), .rdlo_out(a7_wr[534]));
			radix2 #(.width(width)) rd_st6_519  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[519]), .rdlo_in(a6_wr[535]),  .coef_in(coef[448]), .rdup_out(a7_wr[519]), .rdlo_out(a7_wr[535]));
			radix2 #(.width(width)) rd_st6_520  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[520]), .rdlo_in(a6_wr[536]),  .coef_in(coef[512]), .rdup_out(a7_wr[520]), .rdlo_out(a7_wr[536]));
			radix2 #(.width(width)) rd_st6_521  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[521]), .rdlo_in(a6_wr[537]),  .coef_in(coef[576]), .rdup_out(a7_wr[521]), .rdlo_out(a7_wr[537]));
			radix2 #(.width(width)) rd_st6_522  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[522]), .rdlo_in(a6_wr[538]),  .coef_in(coef[640]), .rdup_out(a7_wr[522]), .rdlo_out(a7_wr[538]));
			radix2 #(.width(width)) rd_st6_523  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[523]), .rdlo_in(a6_wr[539]),  .coef_in(coef[704]), .rdup_out(a7_wr[523]), .rdlo_out(a7_wr[539]));
			radix2 #(.width(width)) rd_st6_524  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[524]), .rdlo_in(a6_wr[540]),  .coef_in(coef[768]), .rdup_out(a7_wr[524]), .rdlo_out(a7_wr[540]));
			radix2 #(.width(width)) rd_st6_525  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[525]), .rdlo_in(a6_wr[541]),  .coef_in(coef[832]), .rdup_out(a7_wr[525]), .rdlo_out(a7_wr[541]));
			radix2 #(.width(width)) rd_st6_526  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[526]), .rdlo_in(a6_wr[542]),  .coef_in(coef[896]), .rdup_out(a7_wr[526]), .rdlo_out(a7_wr[542]));
			radix2 #(.width(width)) rd_st6_527  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[527]), .rdlo_in(a6_wr[543]),  .coef_in(coef[960]), .rdup_out(a7_wr[527]), .rdlo_out(a7_wr[543]));
			radix2 #(.width(width)) rd_st6_544  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[544]), .rdlo_in(a6_wr[560]),  .coef_in(coef[0]), .rdup_out(a7_wr[544]), .rdlo_out(a7_wr[560]));
			radix2 #(.width(width)) rd_st6_545  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[545]), .rdlo_in(a6_wr[561]),  .coef_in(coef[64]), .rdup_out(a7_wr[545]), .rdlo_out(a7_wr[561]));
			radix2 #(.width(width)) rd_st6_546  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[546]), .rdlo_in(a6_wr[562]),  .coef_in(coef[128]), .rdup_out(a7_wr[546]), .rdlo_out(a7_wr[562]));
			radix2 #(.width(width)) rd_st6_547  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[547]), .rdlo_in(a6_wr[563]),  .coef_in(coef[192]), .rdup_out(a7_wr[547]), .rdlo_out(a7_wr[563]));
			radix2 #(.width(width)) rd_st6_548  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[548]), .rdlo_in(a6_wr[564]),  .coef_in(coef[256]), .rdup_out(a7_wr[548]), .rdlo_out(a7_wr[564]));
			radix2 #(.width(width)) rd_st6_549  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[549]), .rdlo_in(a6_wr[565]),  .coef_in(coef[320]), .rdup_out(a7_wr[549]), .rdlo_out(a7_wr[565]));
			radix2 #(.width(width)) rd_st6_550  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[550]), .rdlo_in(a6_wr[566]),  .coef_in(coef[384]), .rdup_out(a7_wr[550]), .rdlo_out(a7_wr[566]));
			radix2 #(.width(width)) rd_st6_551  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[551]), .rdlo_in(a6_wr[567]),  .coef_in(coef[448]), .rdup_out(a7_wr[551]), .rdlo_out(a7_wr[567]));
			radix2 #(.width(width)) rd_st6_552  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[552]), .rdlo_in(a6_wr[568]),  .coef_in(coef[512]), .rdup_out(a7_wr[552]), .rdlo_out(a7_wr[568]));
			radix2 #(.width(width)) rd_st6_553  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[553]), .rdlo_in(a6_wr[569]),  .coef_in(coef[576]), .rdup_out(a7_wr[553]), .rdlo_out(a7_wr[569]));
			radix2 #(.width(width)) rd_st6_554  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[554]), .rdlo_in(a6_wr[570]),  .coef_in(coef[640]), .rdup_out(a7_wr[554]), .rdlo_out(a7_wr[570]));
			radix2 #(.width(width)) rd_st6_555  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[555]), .rdlo_in(a6_wr[571]),  .coef_in(coef[704]), .rdup_out(a7_wr[555]), .rdlo_out(a7_wr[571]));
			radix2 #(.width(width)) rd_st6_556  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[556]), .rdlo_in(a6_wr[572]),  .coef_in(coef[768]), .rdup_out(a7_wr[556]), .rdlo_out(a7_wr[572]));
			radix2 #(.width(width)) rd_st6_557  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[557]), .rdlo_in(a6_wr[573]),  .coef_in(coef[832]), .rdup_out(a7_wr[557]), .rdlo_out(a7_wr[573]));
			radix2 #(.width(width)) rd_st6_558  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[558]), .rdlo_in(a6_wr[574]),  .coef_in(coef[896]), .rdup_out(a7_wr[558]), .rdlo_out(a7_wr[574]));
			radix2 #(.width(width)) rd_st6_559  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[559]), .rdlo_in(a6_wr[575]),  .coef_in(coef[960]), .rdup_out(a7_wr[559]), .rdlo_out(a7_wr[575]));
			radix2 #(.width(width)) rd_st6_576  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[576]), .rdlo_in(a6_wr[592]),  .coef_in(coef[0]), .rdup_out(a7_wr[576]), .rdlo_out(a7_wr[592]));
			radix2 #(.width(width)) rd_st6_577  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[577]), .rdlo_in(a6_wr[593]),  .coef_in(coef[64]), .rdup_out(a7_wr[577]), .rdlo_out(a7_wr[593]));
			radix2 #(.width(width)) rd_st6_578  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[578]), .rdlo_in(a6_wr[594]),  .coef_in(coef[128]), .rdup_out(a7_wr[578]), .rdlo_out(a7_wr[594]));
			radix2 #(.width(width)) rd_st6_579  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[579]), .rdlo_in(a6_wr[595]),  .coef_in(coef[192]), .rdup_out(a7_wr[579]), .rdlo_out(a7_wr[595]));
			radix2 #(.width(width)) rd_st6_580  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[580]), .rdlo_in(a6_wr[596]),  .coef_in(coef[256]), .rdup_out(a7_wr[580]), .rdlo_out(a7_wr[596]));
			radix2 #(.width(width)) rd_st6_581  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[581]), .rdlo_in(a6_wr[597]),  .coef_in(coef[320]), .rdup_out(a7_wr[581]), .rdlo_out(a7_wr[597]));
			radix2 #(.width(width)) rd_st6_582  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[582]), .rdlo_in(a6_wr[598]),  .coef_in(coef[384]), .rdup_out(a7_wr[582]), .rdlo_out(a7_wr[598]));
			radix2 #(.width(width)) rd_st6_583  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[583]), .rdlo_in(a6_wr[599]),  .coef_in(coef[448]), .rdup_out(a7_wr[583]), .rdlo_out(a7_wr[599]));
			radix2 #(.width(width)) rd_st6_584  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[584]), .rdlo_in(a6_wr[600]),  .coef_in(coef[512]), .rdup_out(a7_wr[584]), .rdlo_out(a7_wr[600]));
			radix2 #(.width(width)) rd_st6_585  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[585]), .rdlo_in(a6_wr[601]),  .coef_in(coef[576]), .rdup_out(a7_wr[585]), .rdlo_out(a7_wr[601]));
			radix2 #(.width(width)) rd_st6_586  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[586]), .rdlo_in(a6_wr[602]),  .coef_in(coef[640]), .rdup_out(a7_wr[586]), .rdlo_out(a7_wr[602]));
			radix2 #(.width(width)) rd_st6_587  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[587]), .rdlo_in(a6_wr[603]),  .coef_in(coef[704]), .rdup_out(a7_wr[587]), .rdlo_out(a7_wr[603]));
			radix2 #(.width(width)) rd_st6_588  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[588]), .rdlo_in(a6_wr[604]),  .coef_in(coef[768]), .rdup_out(a7_wr[588]), .rdlo_out(a7_wr[604]));
			radix2 #(.width(width)) rd_st6_589  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[589]), .rdlo_in(a6_wr[605]),  .coef_in(coef[832]), .rdup_out(a7_wr[589]), .rdlo_out(a7_wr[605]));
			radix2 #(.width(width)) rd_st6_590  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[590]), .rdlo_in(a6_wr[606]),  .coef_in(coef[896]), .rdup_out(a7_wr[590]), .rdlo_out(a7_wr[606]));
			radix2 #(.width(width)) rd_st6_591  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[591]), .rdlo_in(a6_wr[607]),  .coef_in(coef[960]), .rdup_out(a7_wr[591]), .rdlo_out(a7_wr[607]));
			radix2 #(.width(width)) rd_st6_608  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[608]), .rdlo_in(a6_wr[624]),  .coef_in(coef[0]), .rdup_out(a7_wr[608]), .rdlo_out(a7_wr[624]));
			radix2 #(.width(width)) rd_st6_609  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[609]), .rdlo_in(a6_wr[625]),  .coef_in(coef[64]), .rdup_out(a7_wr[609]), .rdlo_out(a7_wr[625]));
			radix2 #(.width(width)) rd_st6_610  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[610]), .rdlo_in(a6_wr[626]),  .coef_in(coef[128]), .rdup_out(a7_wr[610]), .rdlo_out(a7_wr[626]));
			radix2 #(.width(width)) rd_st6_611  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[611]), .rdlo_in(a6_wr[627]),  .coef_in(coef[192]), .rdup_out(a7_wr[611]), .rdlo_out(a7_wr[627]));
			radix2 #(.width(width)) rd_st6_612  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[612]), .rdlo_in(a6_wr[628]),  .coef_in(coef[256]), .rdup_out(a7_wr[612]), .rdlo_out(a7_wr[628]));
			radix2 #(.width(width)) rd_st6_613  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[613]), .rdlo_in(a6_wr[629]),  .coef_in(coef[320]), .rdup_out(a7_wr[613]), .rdlo_out(a7_wr[629]));
			radix2 #(.width(width)) rd_st6_614  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[614]), .rdlo_in(a6_wr[630]),  .coef_in(coef[384]), .rdup_out(a7_wr[614]), .rdlo_out(a7_wr[630]));
			radix2 #(.width(width)) rd_st6_615  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[615]), .rdlo_in(a6_wr[631]),  .coef_in(coef[448]), .rdup_out(a7_wr[615]), .rdlo_out(a7_wr[631]));
			radix2 #(.width(width)) rd_st6_616  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[616]), .rdlo_in(a6_wr[632]),  .coef_in(coef[512]), .rdup_out(a7_wr[616]), .rdlo_out(a7_wr[632]));
			radix2 #(.width(width)) rd_st6_617  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[617]), .rdlo_in(a6_wr[633]),  .coef_in(coef[576]), .rdup_out(a7_wr[617]), .rdlo_out(a7_wr[633]));
			radix2 #(.width(width)) rd_st6_618  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[618]), .rdlo_in(a6_wr[634]),  .coef_in(coef[640]), .rdup_out(a7_wr[618]), .rdlo_out(a7_wr[634]));
			radix2 #(.width(width)) rd_st6_619  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[619]), .rdlo_in(a6_wr[635]),  .coef_in(coef[704]), .rdup_out(a7_wr[619]), .rdlo_out(a7_wr[635]));
			radix2 #(.width(width)) rd_st6_620  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[620]), .rdlo_in(a6_wr[636]),  .coef_in(coef[768]), .rdup_out(a7_wr[620]), .rdlo_out(a7_wr[636]));
			radix2 #(.width(width)) rd_st6_621  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[621]), .rdlo_in(a6_wr[637]),  .coef_in(coef[832]), .rdup_out(a7_wr[621]), .rdlo_out(a7_wr[637]));
			radix2 #(.width(width)) rd_st6_622  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[622]), .rdlo_in(a6_wr[638]),  .coef_in(coef[896]), .rdup_out(a7_wr[622]), .rdlo_out(a7_wr[638]));
			radix2 #(.width(width)) rd_st6_623  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[623]), .rdlo_in(a6_wr[639]),  .coef_in(coef[960]), .rdup_out(a7_wr[623]), .rdlo_out(a7_wr[639]));
			radix2 #(.width(width)) rd_st6_640  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[640]), .rdlo_in(a6_wr[656]),  .coef_in(coef[0]), .rdup_out(a7_wr[640]), .rdlo_out(a7_wr[656]));
			radix2 #(.width(width)) rd_st6_641  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[641]), .rdlo_in(a6_wr[657]),  .coef_in(coef[64]), .rdup_out(a7_wr[641]), .rdlo_out(a7_wr[657]));
			radix2 #(.width(width)) rd_st6_642  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[642]), .rdlo_in(a6_wr[658]),  .coef_in(coef[128]), .rdup_out(a7_wr[642]), .rdlo_out(a7_wr[658]));
			radix2 #(.width(width)) rd_st6_643  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[643]), .rdlo_in(a6_wr[659]),  .coef_in(coef[192]), .rdup_out(a7_wr[643]), .rdlo_out(a7_wr[659]));
			radix2 #(.width(width)) rd_st6_644  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[644]), .rdlo_in(a6_wr[660]),  .coef_in(coef[256]), .rdup_out(a7_wr[644]), .rdlo_out(a7_wr[660]));
			radix2 #(.width(width)) rd_st6_645  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[645]), .rdlo_in(a6_wr[661]),  .coef_in(coef[320]), .rdup_out(a7_wr[645]), .rdlo_out(a7_wr[661]));
			radix2 #(.width(width)) rd_st6_646  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[646]), .rdlo_in(a6_wr[662]),  .coef_in(coef[384]), .rdup_out(a7_wr[646]), .rdlo_out(a7_wr[662]));
			radix2 #(.width(width)) rd_st6_647  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[647]), .rdlo_in(a6_wr[663]),  .coef_in(coef[448]), .rdup_out(a7_wr[647]), .rdlo_out(a7_wr[663]));
			radix2 #(.width(width)) rd_st6_648  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[648]), .rdlo_in(a6_wr[664]),  .coef_in(coef[512]), .rdup_out(a7_wr[648]), .rdlo_out(a7_wr[664]));
			radix2 #(.width(width)) rd_st6_649  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[649]), .rdlo_in(a6_wr[665]),  .coef_in(coef[576]), .rdup_out(a7_wr[649]), .rdlo_out(a7_wr[665]));
			radix2 #(.width(width)) rd_st6_650  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[650]), .rdlo_in(a6_wr[666]),  .coef_in(coef[640]), .rdup_out(a7_wr[650]), .rdlo_out(a7_wr[666]));
			radix2 #(.width(width)) rd_st6_651  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[651]), .rdlo_in(a6_wr[667]),  .coef_in(coef[704]), .rdup_out(a7_wr[651]), .rdlo_out(a7_wr[667]));
			radix2 #(.width(width)) rd_st6_652  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[652]), .rdlo_in(a6_wr[668]),  .coef_in(coef[768]), .rdup_out(a7_wr[652]), .rdlo_out(a7_wr[668]));
			radix2 #(.width(width)) rd_st6_653  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[653]), .rdlo_in(a6_wr[669]),  .coef_in(coef[832]), .rdup_out(a7_wr[653]), .rdlo_out(a7_wr[669]));
			radix2 #(.width(width)) rd_st6_654  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[654]), .rdlo_in(a6_wr[670]),  .coef_in(coef[896]), .rdup_out(a7_wr[654]), .rdlo_out(a7_wr[670]));
			radix2 #(.width(width)) rd_st6_655  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[655]), .rdlo_in(a6_wr[671]),  .coef_in(coef[960]), .rdup_out(a7_wr[655]), .rdlo_out(a7_wr[671]));
			radix2 #(.width(width)) rd_st6_672  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[672]), .rdlo_in(a6_wr[688]),  .coef_in(coef[0]), .rdup_out(a7_wr[672]), .rdlo_out(a7_wr[688]));
			radix2 #(.width(width)) rd_st6_673  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[673]), .rdlo_in(a6_wr[689]),  .coef_in(coef[64]), .rdup_out(a7_wr[673]), .rdlo_out(a7_wr[689]));
			radix2 #(.width(width)) rd_st6_674  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[674]), .rdlo_in(a6_wr[690]),  .coef_in(coef[128]), .rdup_out(a7_wr[674]), .rdlo_out(a7_wr[690]));
			radix2 #(.width(width)) rd_st6_675  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[675]), .rdlo_in(a6_wr[691]),  .coef_in(coef[192]), .rdup_out(a7_wr[675]), .rdlo_out(a7_wr[691]));
			radix2 #(.width(width)) rd_st6_676  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[676]), .rdlo_in(a6_wr[692]),  .coef_in(coef[256]), .rdup_out(a7_wr[676]), .rdlo_out(a7_wr[692]));
			radix2 #(.width(width)) rd_st6_677  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[677]), .rdlo_in(a6_wr[693]),  .coef_in(coef[320]), .rdup_out(a7_wr[677]), .rdlo_out(a7_wr[693]));
			radix2 #(.width(width)) rd_st6_678  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[678]), .rdlo_in(a6_wr[694]),  .coef_in(coef[384]), .rdup_out(a7_wr[678]), .rdlo_out(a7_wr[694]));
			radix2 #(.width(width)) rd_st6_679  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[679]), .rdlo_in(a6_wr[695]),  .coef_in(coef[448]), .rdup_out(a7_wr[679]), .rdlo_out(a7_wr[695]));
			radix2 #(.width(width)) rd_st6_680  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[680]), .rdlo_in(a6_wr[696]),  .coef_in(coef[512]), .rdup_out(a7_wr[680]), .rdlo_out(a7_wr[696]));
			radix2 #(.width(width)) rd_st6_681  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[681]), .rdlo_in(a6_wr[697]),  .coef_in(coef[576]), .rdup_out(a7_wr[681]), .rdlo_out(a7_wr[697]));
			radix2 #(.width(width)) rd_st6_682  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[682]), .rdlo_in(a6_wr[698]),  .coef_in(coef[640]), .rdup_out(a7_wr[682]), .rdlo_out(a7_wr[698]));
			radix2 #(.width(width)) rd_st6_683  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[683]), .rdlo_in(a6_wr[699]),  .coef_in(coef[704]), .rdup_out(a7_wr[683]), .rdlo_out(a7_wr[699]));
			radix2 #(.width(width)) rd_st6_684  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[684]), .rdlo_in(a6_wr[700]),  .coef_in(coef[768]), .rdup_out(a7_wr[684]), .rdlo_out(a7_wr[700]));
			radix2 #(.width(width)) rd_st6_685  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[685]), .rdlo_in(a6_wr[701]),  .coef_in(coef[832]), .rdup_out(a7_wr[685]), .rdlo_out(a7_wr[701]));
			radix2 #(.width(width)) rd_st6_686  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[686]), .rdlo_in(a6_wr[702]),  .coef_in(coef[896]), .rdup_out(a7_wr[686]), .rdlo_out(a7_wr[702]));
			radix2 #(.width(width)) rd_st6_687  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[687]), .rdlo_in(a6_wr[703]),  .coef_in(coef[960]), .rdup_out(a7_wr[687]), .rdlo_out(a7_wr[703]));
			radix2 #(.width(width)) rd_st6_704  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[704]), .rdlo_in(a6_wr[720]),  .coef_in(coef[0]), .rdup_out(a7_wr[704]), .rdlo_out(a7_wr[720]));
			radix2 #(.width(width)) rd_st6_705  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[705]), .rdlo_in(a6_wr[721]),  .coef_in(coef[64]), .rdup_out(a7_wr[705]), .rdlo_out(a7_wr[721]));
			radix2 #(.width(width)) rd_st6_706  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[706]), .rdlo_in(a6_wr[722]),  .coef_in(coef[128]), .rdup_out(a7_wr[706]), .rdlo_out(a7_wr[722]));
			radix2 #(.width(width)) rd_st6_707  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[707]), .rdlo_in(a6_wr[723]),  .coef_in(coef[192]), .rdup_out(a7_wr[707]), .rdlo_out(a7_wr[723]));
			radix2 #(.width(width)) rd_st6_708  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[708]), .rdlo_in(a6_wr[724]),  .coef_in(coef[256]), .rdup_out(a7_wr[708]), .rdlo_out(a7_wr[724]));
			radix2 #(.width(width)) rd_st6_709  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[709]), .rdlo_in(a6_wr[725]),  .coef_in(coef[320]), .rdup_out(a7_wr[709]), .rdlo_out(a7_wr[725]));
			radix2 #(.width(width)) rd_st6_710  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[710]), .rdlo_in(a6_wr[726]),  .coef_in(coef[384]), .rdup_out(a7_wr[710]), .rdlo_out(a7_wr[726]));
			radix2 #(.width(width)) rd_st6_711  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[711]), .rdlo_in(a6_wr[727]),  .coef_in(coef[448]), .rdup_out(a7_wr[711]), .rdlo_out(a7_wr[727]));
			radix2 #(.width(width)) rd_st6_712  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[712]), .rdlo_in(a6_wr[728]),  .coef_in(coef[512]), .rdup_out(a7_wr[712]), .rdlo_out(a7_wr[728]));
			radix2 #(.width(width)) rd_st6_713  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[713]), .rdlo_in(a6_wr[729]),  .coef_in(coef[576]), .rdup_out(a7_wr[713]), .rdlo_out(a7_wr[729]));
			radix2 #(.width(width)) rd_st6_714  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[714]), .rdlo_in(a6_wr[730]),  .coef_in(coef[640]), .rdup_out(a7_wr[714]), .rdlo_out(a7_wr[730]));
			radix2 #(.width(width)) rd_st6_715  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[715]), .rdlo_in(a6_wr[731]),  .coef_in(coef[704]), .rdup_out(a7_wr[715]), .rdlo_out(a7_wr[731]));
			radix2 #(.width(width)) rd_st6_716  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[716]), .rdlo_in(a6_wr[732]),  .coef_in(coef[768]), .rdup_out(a7_wr[716]), .rdlo_out(a7_wr[732]));
			radix2 #(.width(width)) rd_st6_717  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[717]), .rdlo_in(a6_wr[733]),  .coef_in(coef[832]), .rdup_out(a7_wr[717]), .rdlo_out(a7_wr[733]));
			radix2 #(.width(width)) rd_st6_718  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[718]), .rdlo_in(a6_wr[734]),  .coef_in(coef[896]), .rdup_out(a7_wr[718]), .rdlo_out(a7_wr[734]));
			radix2 #(.width(width)) rd_st6_719  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[719]), .rdlo_in(a6_wr[735]),  .coef_in(coef[960]), .rdup_out(a7_wr[719]), .rdlo_out(a7_wr[735]));
			radix2 #(.width(width)) rd_st6_736  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[736]), .rdlo_in(a6_wr[752]),  .coef_in(coef[0]), .rdup_out(a7_wr[736]), .rdlo_out(a7_wr[752]));
			radix2 #(.width(width)) rd_st6_737  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[737]), .rdlo_in(a6_wr[753]),  .coef_in(coef[64]), .rdup_out(a7_wr[737]), .rdlo_out(a7_wr[753]));
			radix2 #(.width(width)) rd_st6_738  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[738]), .rdlo_in(a6_wr[754]),  .coef_in(coef[128]), .rdup_out(a7_wr[738]), .rdlo_out(a7_wr[754]));
			radix2 #(.width(width)) rd_st6_739  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[739]), .rdlo_in(a6_wr[755]),  .coef_in(coef[192]), .rdup_out(a7_wr[739]), .rdlo_out(a7_wr[755]));
			radix2 #(.width(width)) rd_st6_740  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[740]), .rdlo_in(a6_wr[756]),  .coef_in(coef[256]), .rdup_out(a7_wr[740]), .rdlo_out(a7_wr[756]));
			radix2 #(.width(width)) rd_st6_741  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[741]), .rdlo_in(a6_wr[757]),  .coef_in(coef[320]), .rdup_out(a7_wr[741]), .rdlo_out(a7_wr[757]));
			radix2 #(.width(width)) rd_st6_742  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[742]), .rdlo_in(a6_wr[758]),  .coef_in(coef[384]), .rdup_out(a7_wr[742]), .rdlo_out(a7_wr[758]));
			radix2 #(.width(width)) rd_st6_743  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[743]), .rdlo_in(a6_wr[759]),  .coef_in(coef[448]), .rdup_out(a7_wr[743]), .rdlo_out(a7_wr[759]));
			radix2 #(.width(width)) rd_st6_744  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[744]), .rdlo_in(a6_wr[760]),  .coef_in(coef[512]), .rdup_out(a7_wr[744]), .rdlo_out(a7_wr[760]));
			radix2 #(.width(width)) rd_st6_745  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[745]), .rdlo_in(a6_wr[761]),  .coef_in(coef[576]), .rdup_out(a7_wr[745]), .rdlo_out(a7_wr[761]));
			radix2 #(.width(width)) rd_st6_746  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[746]), .rdlo_in(a6_wr[762]),  .coef_in(coef[640]), .rdup_out(a7_wr[746]), .rdlo_out(a7_wr[762]));
			radix2 #(.width(width)) rd_st6_747  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[747]), .rdlo_in(a6_wr[763]),  .coef_in(coef[704]), .rdup_out(a7_wr[747]), .rdlo_out(a7_wr[763]));
			radix2 #(.width(width)) rd_st6_748  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[748]), .rdlo_in(a6_wr[764]),  .coef_in(coef[768]), .rdup_out(a7_wr[748]), .rdlo_out(a7_wr[764]));
			radix2 #(.width(width)) rd_st6_749  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[749]), .rdlo_in(a6_wr[765]),  .coef_in(coef[832]), .rdup_out(a7_wr[749]), .rdlo_out(a7_wr[765]));
			radix2 #(.width(width)) rd_st6_750  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[750]), .rdlo_in(a6_wr[766]),  .coef_in(coef[896]), .rdup_out(a7_wr[750]), .rdlo_out(a7_wr[766]));
			radix2 #(.width(width)) rd_st6_751  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[751]), .rdlo_in(a6_wr[767]),  .coef_in(coef[960]), .rdup_out(a7_wr[751]), .rdlo_out(a7_wr[767]));
			radix2 #(.width(width)) rd_st6_768  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[768]), .rdlo_in(a6_wr[784]),  .coef_in(coef[0]), .rdup_out(a7_wr[768]), .rdlo_out(a7_wr[784]));
			radix2 #(.width(width)) rd_st6_769  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[769]), .rdlo_in(a6_wr[785]),  .coef_in(coef[64]), .rdup_out(a7_wr[769]), .rdlo_out(a7_wr[785]));
			radix2 #(.width(width)) rd_st6_770  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[770]), .rdlo_in(a6_wr[786]),  .coef_in(coef[128]), .rdup_out(a7_wr[770]), .rdlo_out(a7_wr[786]));
			radix2 #(.width(width)) rd_st6_771  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[771]), .rdlo_in(a6_wr[787]),  .coef_in(coef[192]), .rdup_out(a7_wr[771]), .rdlo_out(a7_wr[787]));
			radix2 #(.width(width)) rd_st6_772  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[772]), .rdlo_in(a6_wr[788]),  .coef_in(coef[256]), .rdup_out(a7_wr[772]), .rdlo_out(a7_wr[788]));
			radix2 #(.width(width)) rd_st6_773  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[773]), .rdlo_in(a6_wr[789]),  .coef_in(coef[320]), .rdup_out(a7_wr[773]), .rdlo_out(a7_wr[789]));
			radix2 #(.width(width)) rd_st6_774  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[774]), .rdlo_in(a6_wr[790]),  .coef_in(coef[384]), .rdup_out(a7_wr[774]), .rdlo_out(a7_wr[790]));
			radix2 #(.width(width)) rd_st6_775  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[775]), .rdlo_in(a6_wr[791]),  .coef_in(coef[448]), .rdup_out(a7_wr[775]), .rdlo_out(a7_wr[791]));
			radix2 #(.width(width)) rd_st6_776  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[776]), .rdlo_in(a6_wr[792]),  .coef_in(coef[512]), .rdup_out(a7_wr[776]), .rdlo_out(a7_wr[792]));
			radix2 #(.width(width)) rd_st6_777  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[777]), .rdlo_in(a6_wr[793]),  .coef_in(coef[576]), .rdup_out(a7_wr[777]), .rdlo_out(a7_wr[793]));
			radix2 #(.width(width)) rd_st6_778  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[778]), .rdlo_in(a6_wr[794]),  .coef_in(coef[640]), .rdup_out(a7_wr[778]), .rdlo_out(a7_wr[794]));
			radix2 #(.width(width)) rd_st6_779  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[779]), .rdlo_in(a6_wr[795]),  .coef_in(coef[704]), .rdup_out(a7_wr[779]), .rdlo_out(a7_wr[795]));
			radix2 #(.width(width)) rd_st6_780  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[780]), .rdlo_in(a6_wr[796]),  .coef_in(coef[768]), .rdup_out(a7_wr[780]), .rdlo_out(a7_wr[796]));
			radix2 #(.width(width)) rd_st6_781  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[781]), .rdlo_in(a6_wr[797]),  .coef_in(coef[832]), .rdup_out(a7_wr[781]), .rdlo_out(a7_wr[797]));
			radix2 #(.width(width)) rd_st6_782  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[782]), .rdlo_in(a6_wr[798]),  .coef_in(coef[896]), .rdup_out(a7_wr[782]), .rdlo_out(a7_wr[798]));
			radix2 #(.width(width)) rd_st6_783  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[783]), .rdlo_in(a6_wr[799]),  .coef_in(coef[960]), .rdup_out(a7_wr[783]), .rdlo_out(a7_wr[799]));
			radix2 #(.width(width)) rd_st6_800  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[800]), .rdlo_in(a6_wr[816]),  .coef_in(coef[0]), .rdup_out(a7_wr[800]), .rdlo_out(a7_wr[816]));
			radix2 #(.width(width)) rd_st6_801  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[801]), .rdlo_in(a6_wr[817]),  .coef_in(coef[64]), .rdup_out(a7_wr[801]), .rdlo_out(a7_wr[817]));
			radix2 #(.width(width)) rd_st6_802  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[802]), .rdlo_in(a6_wr[818]),  .coef_in(coef[128]), .rdup_out(a7_wr[802]), .rdlo_out(a7_wr[818]));
			radix2 #(.width(width)) rd_st6_803  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[803]), .rdlo_in(a6_wr[819]),  .coef_in(coef[192]), .rdup_out(a7_wr[803]), .rdlo_out(a7_wr[819]));
			radix2 #(.width(width)) rd_st6_804  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[804]), .rdlo_in(a6_wr[820]),  .coef_in(coef[256]), .rdup_out(a7_wr[804]), .rdlo_out(a7_wr[820]));
			radix2 #(.width(width)) rd_st6_805  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[805]), .rdlo_in(a6_wr[821]),  .coef_in(coef[320]), .rdup_out(a7_wr[805]), .rdlo_out(a7_wr[821]));
			radix2 #(.width(width)) rd_st6_806  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[806]), .rdlo_in(a6_wr[822]),  .coef_in(coef[384]), .rdup_out(a7_wr[806]), .rdlo_out(a7_wr[822]));
			radix2 #(.width(width)) rd_st6_807  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[807]), .rdlo_in(a6_wr[823]),  .coef_in(coef[448]), .rdup_out(a7_wr[807]), .rdlo_out(a7_wr[823]));
			radix2 #(.width(width)) rd_st6_808  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[808]), .rdlo_in(a6_wr[824]),  .coef_in(coef[512]), .rdup_out(a7_wr[808]), .rdlo_out(a7_wr[824]));
			radix2 #(.width(width)) rd_st6_809  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[809]), .rdlo_in(a6_wr[825]),  .coef_in(coef[576]), .rdup_out(a7_wr[809]), .rdlo_out(a7_wr[825]));
			radix2 #(.width(width)) rd_st6_810  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[810]), .rdlo_in(a6_wr[826]),  .coef_in(coef[640]), .rdup_out(a7_wr[810]), .rdlo_out(a7_wr[826]));
			radix2 #(.width(width)) rd_st6_811  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[811]), .rdlo_in(a6_wr[827]),  .coef_in(coef[704]), .rdup_out(a7_wr[811]), .rdlo_out(a7_wr[827]));
			radix2 #(.width(width)) rd_st6_812  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[812]), .rdlo_in(a6_wr[828]),  .coef_in(coef[768]), .rdup_out(a7_wr[812]), .rdlo_out(a7_wr[828]));
			radix2 #(.width(width)) rd_st6_813  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[813]), .rdlo_in(a6_wr[829]),  .coef_in(coef[832]), .rdup_out(a7_wr[813]), .rdlo_out(a7_wr[829]));
			radix2 #(.width(width)) rd_st6_814  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[814]), .rdlo_in(a6_wr[830]),  .coef_in(coef[896]), .rdup_out(a7_wr[814]), .rdlo_out(a7_wr[830]));
			radix2 #(.width(width)) rd_st6_815  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[815]), .rdlo_in(a6_wr[831]),  .coef_in(coef[960]), .rdup_out(a7_wr[815]), .rdlo_out(a7_wr[831]));
			radix2 #(.width(width)) rd_st6_832  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[832]), .rdlo_in(a6_wr[848]),  .coef_in(coef[0]), .rdup_out(a7_wr[832]), .rdlo_out(a7_wr[848]));
			radix2 #(.width(width)) rd_st6_833  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[833]), .rdlo_in(a6_wr[849]),  .coef_in(coef[64]), .rdup_out(a7_wr[833]), .rdlo_out(a7_wr[849]));
			radix2 #(.width(width)) rd_st6_834  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[834]), .rdlo_in(a6_wr[850]),  .coef_in(coef[128]), .rdup_out(a7_wr[834]), .rdlo_out(a7_wr[850]));
			radix2 #(.width(width)) rd_st6_835  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[835]), .rdlo_in(a6_wr[851]),  .coef_in(coef[192]), .rdup_out(a7_wr[835]), .rdlo_out(a7_wr[851]));
			radix2 #(.width(width)) rd_st6_836  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[836]), .rdlo_in(a6_wr[852]),  .coef_in(coef[256]), .rdup_out(a7_wr[836]), .rdlo_out(a7_wr[852]));
			radix2 #(.width(width)) rd_st6_837  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[837]), .rdlo_in(a6_wr[853]),  .coef_in(coef[320]), .rdup_out(a7_wr[837]), .rdlo_out(a7_wr[853]));
			radix2 #(.width(width)) rd_st6_838  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[838]), .rdlo_in(a6_wr[854]),  .coef_in(coef[384]), .rdup_out(a7_wr[838]), .rdlo_out(a7_wr[854]));
			radix2 #(.width(width)) rd_st6_839  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[839]), .rdlo_in(a6_wr[855]),  .coef_in(coef[448]), .rdup_out(a7_wr[839]), .rdlo_out(a7_wr[855]));
			radix2 #(.width(width)) rd_st6_840  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[840]), .rdlo_in(a6_wr[856]),  .coef_in(coef[512]), .rdup_out(a7_wr[840]), .rdlo_out(a7_wr[856]));
			radix2 #(.width(width)) rd_st6_841  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[841]), .rdlo_in(a6_wr[857]),  .coef_in(coef[576]), .rdup_out(a7_wr[841]), .rdlo_out(a7_wr[857]));
			radix2 #(.width(width)) rd_st6_842  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[842]), .rdlo_in(a6_wr[858]),  .coef_in(coef[640]), .rdup_out(a7_wr[842]), .rdlo_out(a7_wr[858]));
			radix2 #(.width(width)) rd_st6_843  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[843]), .rdlo_in(a6_wr[859]),  .coef_in(coef[704]), .rdup_out(a7_wr[843]), .rdlo_out(a7_wr[859]));
			radix2 #(.width(width)) rd_st6_844  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[844]), .rdlo_in(a6_wr[860]),  .coef_in(coef[768]), .rdup_out(a7_wr[844]), .rdlo_out(a7_wr[860]));
			radix2 #(.width(width)) rd_st6_845  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[845]), .rdlo_in(a6_wr[861]),  .coef_in(coef[832]), .rdup_out(a7_wr[845]), .rdlo_out(a7_wr[861]));
			radix2 #(.width(width)) rd_st6_846  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[846]), .rdlo_in(a6_wr[862]),  .coef_in(coef[896]), .rdup_out(a7_wr[846]), .rdlo_out(a7_wr[862]));
			radix2 #(.width(width)) rd_st6_847  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[847]), .rdlo_in(a6_wr[863]),  .coef_in(coef[960]), .rdup_out(a7_wr[847]), .rdlo_out(a7_wr[863]));
			radix2 #(.width(width)) rd_st6_864  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[864]), .rdlo_in(a6_wr[880]),  .coef_in(coef[0]), .rdup_out(a7_wr[864]), .rdlo_out(a7_wr[880]));
			radix2 #(.width(width)) rd_st6_865  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[865]), .rdlo_in(a6_wr[881]),  .coef_in(coef[64]), .rdup_out(a7_wr[865]), .rdlo_out(a7_wr[881]));
			radix2 #(.width(width)) rd_st6_866  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[866]), .rdlo_in(a6_wr[882]),  .coef_in(coef[128]), .rdup_out(a7_wr[866]), .rdlo_out(a7_wr[882]));
			radix2 #(.width(width)) rd_st6_867  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[867]), .rdlo_in(a6_wr[883]),  .coef_in(coef[192]), .rdup_out(a7_wr[867]), .rdlo_out(a7_wr[883]));
			radix2 #(.width(width)) rd_st6_868  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[868]), .rdlo_in(a6_wr[884]),  .coef_in(coef[256]), .rdup_out(a7_wr[868]), .rdlo_out(a7_wr[884]));
			radix2 #(.width(width)) rd_st6_869  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[869]), .rdlo_in(a6_wr[885]),  .coef_in(coef[320]), .rdup_out(a7_wr[869]), .rdlo_out(a7_wr[885]));
			radix2 #(.width(width)) rd_st6_870  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[870]), .rdlo_in(a6_wr[886]),  .coef_in(coef[384]), .rdup_out(a7_wr[870]), .rdlo_out(a7_wr[886]));
			radix2 #(.width(width)) rd_st6_871  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[871]), .rdlo_in(a6_wr[887]),  .coef_in(coef[448]), .rdup_out(a7_wr[871]), .rdlo_out(a7_wr[887]));
			radix2 #(.width(width)) rd_st6_872  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[872]), .rdlo_in(a6_wr[888]),  .coef_in(coef[512]), .rdup_out(a7_wr[872]), .rdlo_out(a7_wr[888]));
			radix2 #(.width(width)) rd_st6_873  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[873]), .rdlo_in(a6_wr[889]),  .coef_in(coef[576]), .rdup_out(a7_wr[873]), .rdlo_out(a7_wr[889]));
			radix2 #(.width(width)) rd_st6_874  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[874]), .rdlo_in(a6_wr[890]),  .coef_in(coef[640]), .rdup_out(a7_wr[874]), .rdlo_out(a7_wr[890]));
			radix2 #(.width(width)) rd_st6_875  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[875]), .rdlo_in(a6_wr[891]),  .coef_in(coef[704]), .rdup_out(a7_wr[875]), .rdlo_out(a7_wr[891]));
			radix2 #(.width(width)) rd_st6_876  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[876]), .rdlo_in(a6_wr[892]),  .coef_in(coef[768]), .rdup_out(a7_wr[876]), .rdlo_out(a7_wr[892]));
			radix2 #(.width(width)) rd_st6_877  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[877]), .rdlo_in(a6_wr[893]),  .coef_in(coef[832]), .rdup_out(a7_wr[877]), .rdlo_out(a7_wr[893]));
			radix2 #(.width(width)) rd_st6_878  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[878]), .rdlo_in(a6_wr[894]),  .coef_in(coef[896]), .rdup_out(a7_wr[878]), .rdlo_out(a7_wr[894]));
			radix2 #(.width(width)) rd_st6_879  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[879]), .rdlo_in(a6_wr[895]),  .coef_in(coef[960]), .rdup_out(a7_wr[879]), .rdlo_out(a7_wr[895]));
			radix2 #(.width(width)) rd_st6_896  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[896]), .rdlo_in(a6_wr[912]),  .coef_in(coef[0]), .rdup_out(a7_wr[896]), .rdlo_out(a7_wr[912]));
			radix2 #(.width(width)) rd_st6_897  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[897]), .rdlo_in(a6_wr[913]),  .coef_in(coef[64]), .rdup_out(a7_wr[897]), .rdlo_out(a7_wr[913]));
			radix2 #(.width(width)) rd_st6_898  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[898]), .rdlo_in(a6_wr[914]),  .coef_in(coef[128]), .rdup_out(a7_wr[898]), .rdlo_out(a7_wr[914]));
			radix2 #(.width(width)) rd_st6_899  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[899]), .rdlo_in(a6_wr[915]),  .coef_in(coef[192]), .rdup_out(a7_wr[899]), .rdlo_out(a7_wr[915]));
			radix2 #(.width(width)) rd_st6_900  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[900]), .rdlo_in(a6_wr[916]),  .coef_in(coef[256]), .rdup_out(a7_wr[900]), .rdlo_out(a7_wr[916]));
			radix2 #(.width(width)) rd_st6_901  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[901]), .rdlo_in(a6_wr[917]),  .coef_in(coef[320]), .rdup_out(a7_wr[901]), .rdlo_out(a7_wr[917]));
			radix2 #(.width(width)) rd_st6_902  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[902]), .rdlo_in(a6_wr[918]),  .coef_in(coef[384]), .rdup_out(a7_wr[902]), .rdlo_out(a7_wr[918]));
			radix2 #(.width(width)) rd_st6_903  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[903]), .rdlo_in(a6_wr[919]),  .coef_in(coef[448]), .rdup_out(a7_wr[903]), .rdlo_out(a7_wr[919]));
			radix2 #(.width(width)) rd_st6_904  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[904]), .rdlo_in(a6_wr[920]),  .coef_in(coef[512]), .rdup_out(a7_wr[904]), .rdlo_out(a7_wr[920]));
			radix2 #(.width(width)) rd_st6_905  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[905]), .rdlo_in(a6_wr[921]),  .coef_in(coef[576]), .rdup_out(a7_wr[905]), .rdlo_out(a7_wr[921]));
			radix2 #(.width(width)) rd_st6_906  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[906]), .rdlo_in(a6_wr[922]),  .coef_in(coef[640]), .rdup_out(a7_wr[906]), .rdlo_out(a7_wr[922]));
			radix2 #(.width(width)) rd_st6_907  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[907]), .rdlo_in(a6_wr[923]),  .coef_in(coef[704]), .rdup_out(a7_wr[907]), .rdlo_out(a7_wr[923]));
			radix2 #(.width(width)) rd_st6_908  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[908]), .rdlo_in(a6_wr[924]),  .coef_in(coef[768]), .rdup_out(a7_wr[908]), .rdlo_out(a7_wr[924]));
			radix2 #(.width(width)) rd_st6_909  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[909]), .rdlo_in(a6_wr[925]),  .coef_in(coef[832]), .rdup_out(a7_wr[909]), .rdlo_out(a7_wr[925]));
			radix2 #(.width(width)) rd_st6_910  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[910]), .rdlo_in(a6_wr[926]),  .coef_in(coef[896]), .rdup_out(a7_wr[910]), .rdlo_out(a7_wr[926]));
			radix2 #(.width(width)) rd_st6_911  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[911]), .rdlo_in(a6_wr[927]),  .coef_in(coef[960]), .rdup_out(a7_wr[911]), .rdlo_out(a7_wr[927]));
			radix2 #(.width(width)) rd_st6_928  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[928]), .rdlo_in(a6_wr[944]),  .coef_in(coef[0]), .rdup_out(a7_wr[928]), .rdlo_out(a7_wr[944]));
			radix2 #(.width(width)) rd_st6_929  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[929]), .rdlo_in(a6_wr[945]),  .coef_in(coef[64]), .rdup_out(a7_wr[929]), .rdlo_out(a7_wr[945]));
			radix2 #(.width(width)) rd_st6_930  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[930]), .rdlo_in(a6_wr[946]),  .coef_in(coef[128]), .rdup_out(a7_wr[930]), .rdlo_out(a7_wr[946]));
			radix2 #(.width(width)) rd_st6_931  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[931]), .rdlo_in(a6_wr[947]),  .coef_in(coef[192]), .rdup_out(a7_wr[931]), .rdlo_out(a7_wr[947]));
			radix2 #(.width(width)) rd_st6_932  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[932]), .rdlo_in(a6_wr[948]),  .coef_in(coef[256]), .rdup_out(a7_wr[932]), .rdlo_out(a7_wr[948]));
			radix2 #(.width(width)) rd_st6_933  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[933]), .rdlo_in(a6_wr[949]),  .coef_in(coef[320]), .rdup_out(a7_wr[933]), .rdlo_out(a7_wr[949]));
			radix2 #(.width(width)) rd_st6_934  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[934]), .rdlo_in(a6_wr[950]),  .coef_in(coef[384]), .rdup_out(a7_wr[934]), .rdlo_out(a7_wr[950]));
			radix2 #(.width(width)) rd_st6_935  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[935]), .rdlo_in(a6_wr[951]),  .coef_in(coef[448]), .rdup_out(a7_wr[935]), .rdlo_out(a7_wr[951]));
			radix2 #(.width(width)) rd_st6_936  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[936]), .rdlo_in(a6_wr[952]),  .coef_in(coef[512]), .rdup_out(a7_wr[936]), .rdlo_out(a7_wr[952]));
			radix2 #(.width(width)) rd_st6_937  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[937]), .rdlo_in(a6_wr[953]),  .coef_in(coef[576]), .rdup_out(a7_wr[937]), .rdlo_out(a7_wr[953]));
			radix2 #(.width(width)) rd_st6_938  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[938]), .rdlo_in(a6_wr[954]),  .coef_in(coef[640]), .rdup_out(a7_wr[938]), .rdlo_out(a7_wr[954]));
			radix2 #(.width(width)) rd_st6_939  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[939]), .rdlo_in(a6_wr[955]),  .coef_in(coef[704]), .rdup_out(a7_wr[939]), .rdlo_out(a7_wr[955]));
			radix2 #(.width(width)) rd_st6_940  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[940]), .rdlo_in(a6_wr[956]),  .coef_in(coef[768]), .rdup_out(a7_wr[940]), .rdlo_out(a7_wr[956]));
			radix2 #(.width(width)) rd_st6_941  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[941]), .rdlo_in(a6_wr[957]),  .coef_in(coef[832]), .rdup_out(a7_wr[941]), .rdlo_out(a7_wr[957]));
			radix2 #(.width(width)) rd_st6_942  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[942]), .rdlo_in(a6_wr[958]),  .coef_in(coef[896]), .rdup_out(a7_wr[942]), .rdlo_out(a7_wr[958]));
			radix2 #(.width(width)) rd_st6_943  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[943]), .rdlo_in(a6_wr[959]),  .coef_in(coef[960]), .rdup_out(a7_wr[943]), .rdlo_out(a7_wr[959]));
			radix2 #(.width(width)) rd_st6_960  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[960]), .rdlo_in(a6_wr[976]),  .coef_in(coef[0]), .rdup_out(a7_wr[960]), .rdlo_out(a7_wr[976]));
			radix2 #(.width(width)) rd_st6_961  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[961]), .rdlo_in(a6_wr[977]),  .coef_in(coef[64]), .rdup_out(a7_wr[961]), .rdlo_out(a7_wr[977]));
			radix2 #(.width(width)) rd_st6_962  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[962]), .rdlo_in(a6_wr[978]),  .coef_in(coef[128]), .rdup_out(a7_wr[962]), .rdlo_out(a7_wr[978]));
			radix2 #(.width(width)) rd_st6_963  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[963]), .rdlo_in(a6_wr[979]),  .coef_in(coef[192]), .rdup_out(a7_wr[963]), .rdlo_out(a7_wr[979]));
			radix2 #(.width(width)) rd_st6_964  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[964]), .rdlo_in(a6_wr[980]),  .coef_in(coef[256]), .rdup_out(a7_wr[964]), .rdlo_out(a7_wr[980]));
			radix2 #(.width(width)) rd_st6_965  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[965]), .rdlo_in(a6_wr[981]),  .coef_in(coef[320]), .rdup_out(a7_wr[965]), .rdlo_out(a7_wr[981]));
			radix2 #(.width(width)) rd_st6_966  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[966]), .rdlo_in(a6_wr[982]),  .coef_in(coef[384]), .rdup_out(a7_wr[966]), .rdlo_out(a7_wr[982]));
			radix2 #(.width(width)) rd_st6_967  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[967]), .rdlo_in(a6_wr[983]),  .coef_in(coef[448]), .rdup_out(a7_wr[967]), .rdlo_out(a7_wr[983]));
			radix2 #(.width(width)) rd_st6_968  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[968]), .rdlo_in(a6_wr[984]),  .coef_in(coef[512]), .rdup_out(a7_wr[968]), .rdlo_out(a7_wr[984]));
			radix2 #(.width(width)) rd_st6_969  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[969]), .rdlo_in(a6_wr[985]),  .coef_in(coef[576]), .rdup_out(a7_wr[969]), .rdlo_out(a7_wr[985]));
			radix2 #(.width(width)) rd_st6_970  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[970]), .rdlo_in(a6_wr[986]),  .coef_in(coef[640]), .rdup_out(a7_wr[970]), .rdlo_out(a7_wr[986]));
			radix2 #(.width(width)) rd_st6_971  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[971]), .rdlo_in(a6_wr[987]),  .coef_in(coef[704]), .rdup_out(a7_wr[971]), .rdlo_out(a7_wr[987]));
			radix2 #(.width(width)) rd_st6_972  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[972]), .rdlo_in(a6_wr[988]),  .coef_in(coef[768]), .rdup_out(a7_wr[972]), .rdlo_out(a7_wr[988]));
			radix2 #(.width(width)) rd_st6_973  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[973]), .rdlo_in(a6_wr[989]),  .coef_in(coef[832]), .rdup_out(a7_wr[973]), .rdlo_out(a7_wr[989]));
			radix2 #(.width(width)) rd_st6_974  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[974]), .rdlo_in(a6_wr[990]),  .coef_in(coef[896]), .rdup_out(a7_wr[974]), .rdlo_out(a7_wr[990]));
			radix2 #(.width(width)) rd_st6_975  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[975]), .rdlo_in(a6_wr[991]),  .coef_in(coef[960]), .rdup_out(a7_wr[975]), .rdlo_out(a7_wr[991]));
			radix2 #(.width(width)) rd_st6_992  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[992]), .rdlo_in(a6_wr[1008]),  .coef_in(coef[0]), .rdup_out(a7_wr[992]), .rdlo_out(a7_wr[1008]));
			radix2 #(.width(width)) rd_st6_993  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[993]), .rdlo_in(a6_wr[1009]),  .coef_in(coef[64]), .rdup_out(a7_wr[993]), .rdlo_out(a7_wr[1009]));
			radix2 #(.width(width)) rd_st6_994  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[994]), .rdlo_in(a6_wr[1010]),  .coef_in(coef[128]), .rdup_out(a7_wr[994]), .rdlo_out(a7_wr[1010]));
			radix2 #(.width(width)) rd_st6_995  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[995]), .rdlo_in(a6_wr[1011]),  .coef_in(coef[192]), .rdup_out(a7_wr[995]), .rdlo_out(a7_wr[1011]));
			radix2 #(.width(width)) rd_st6_996  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[996]), .rdlo_in(a6_wr[1012]),  .coef_in(coef[256]), .rdup_out(a7_wr[996]), .rdlo_out(a7_wr[1012]));
			radix2 #(.width(width)) rd_st6_997  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[997]), .rdlo_in(a6_wr[1013]),  .coef_in(coef[320]), .rdup_out(a7_wr[997]), .rdlo_out(a7_wr[1013]));
			radix2 #(.width(width)) rd_st6_998  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[998]), .rdlo_in(a6_wr[1014]),  .coef_in(coef[384]), .rdup_out(a7_wr[998]), .rdlo_out(a7_wr[1014]));
			radix2 #(.width(width)) rd_st6_999  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[999]), .rdlo_in(a6_wr[1015]),  .coef_in(coef[448]), .rdup_out(a7_wr[999]), .rdlo_out(a7_wr[1015]));
			radix2 #(.width(width)) rd_st6_1000  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1000]), .rdlo_in(a6_wr[1016]),  .coef_in(coef[512]), .rdup_out(a7_wr[1000]), .rdlo_out(a7_wr[1016]));
			radix2 #(.width(width)) rd_st6_1001  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1001]), .rdlo_in(a6_wr[1017]),  .coef_in(coef[576]), .rdup_out(a7_wr[1001]), .rdlo_out(a7_wr[1017]));
			radix2 #(.width(width)) rd_st6_1002  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1002]), .rdlo_in(a6_wr[1018]),  .coef_in(coef[640]), .rdup_out(a7_wr[1002]), .rdlo_out(a7_wr[1018]));
			radix2 #(.width(width)) rd_st6_1003  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1003]), .rdlo_in(a6_wr[1019]),  .coef_in(coef[704]), .rdup_out(a7_wr[1003]), .rdlo_out(a7_wr[1019]));
			radix2 #(.width(width)) rd_st6_1004  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1004]), .rdlo_in(a6_wr[1020]),  .coef_in(coef[768]), .rdup_out(a7_wr[1004]), .rdlo_out(a7_wr[1020]));
			radix2 #(.width(width)) rd_st6_1005  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1005]), .rdlo_in(a6_wr[1021]),  .coef_in(coef[832]), .rdup_out(a7_wr[1005]), .rdlo_out(a7_wr[1021]));
			radix2 #(.width(width)) rd_st6_1006  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1006]), .rdlo_in(a6_wr[1022]),  .coef_in(coef[896]), .rdup_out(a7_wr[1006]), .rdlo_out(a7_wr[1022]));
			radix2 #(.width(width)) rd_st6_1007  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1007]), .rdlo_in(a6_wr[1023]),  .coef_in(coef[960]), .rdup_out(a7_wr[1007]), .rdlo_out(a7_wr[1023]));
			radix2 #(.width(width)) rd_st6_1024  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1024]), .rdlo_in(a6_wr[1040]),  .coef_in(coef[0]), .rdup_out(a7_wr[1024]), .rdlo_out(a7_wr[1040]));
			radix2 #(.width(width)) rd_st6_1025  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1025]), .rdlo_in(a6_wr[1041]),  .coef_in(coef[64]), .rdup_out(a7_wr[1025]), .rdlo_out(a7_wr[1041]));
			radix2 #(.width(width)) rd_st6_1026  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1026]), .rdlo_in(a6_wr[1042]),  .coef_in(coef[128]), .rdup_out(a7_wr[1026]), .rdlo_out(a7_wr[1042]));
			radix2 #(.width(width)) rd_st6_1027  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1027]), .rdlo_in(a6_wr[1043]),  .coef_in(coef[192]), .rdup_out(a7_wr[1027]), .rdlo_out(a7_wr[1043]));
			radix2 #(.width(width)) rd_st6_1028  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1028]), .rdlo_in(a6_wr[1044]),  .coef_in(coef[256]), .rdup_out(a7_wr[1028]), .rdlo_out(a7_wr[1044]));
			radix2 #(.width(width)) rd_st6_1029  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1029]), .rdlo_in(a6_wr[1045]),  .coef_in(coef[320]), .rdup_out(a7_wr[1029]), .rdlo_out(a7_wr[1045]));
			radix2 #(.width(width)) rd_st6_1030  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1030]), .rdlo_in(a6_wr[1046]),  .coef_in(coef[384]), .rdup_out(a7_wr[1030]), .rdlo_out(a7_wr[1046]));
			radix2 #(.width(width)) rd_st6_1031  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1031]), .rdlo_in(a6_wr[1047]),  .coef_in(coef[448]), .rdup_out(a7_wr[1031]), .rdlo_out(a7_wr[1047]));
			radix2 #(.width(width)) rd_st6_1032  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1032]), .rdlo_in(a6_wr[1048]),  .coef_in(coef[512]), .rdup_out(a7_wr[1032]), .rdlo_out(a7_wr[1048]));
			radix2 #(.width(width)) rd_st6_1033  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1033]), .rdlo_in(a6_wr[1049]),  .coef_in(coef[576]), .rdup_out(a7_wr[1033]), .rdlo_out(a7_wr[1049]));
			radix2 #(.width(width)) rd_st6_1034  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1034]), .rdlo_in(a6_wr[1050]),  .coef_in(coef[640]), .rdup_out(a7_wr[1034]), .rdlo_out(a7_wr[1050]));
			radix2 #(.width(width)) rd_st6_1035  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1035]), .rdlo_in(a6_wr[1051]),  .coef_in(coef[704]), .rdup_out(a7_wr[1035]), .rdlo_out(a7_wr[1051]));
			radix2 #(.width(width)) rd_st6_1036  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1036]), .rdlo_in(a6_wr[1052]),  .coef_in(coef[768]), .rdup_out(a7_wr[1036]), .rdlo_out(a7_wr[1052]));
			radix2 #(.width(width)) rd_st6_1037  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1037]), .rdlo_in(a6_wr[1053]),  .coef_in(coef[832]), .rdup_out(a7_wr[1037]), .rdlo_out(a7_wr[1053]));
			radix2 #(.width(width)) rd_st6_1038  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1038]), .rdlo_in(a6_wr[1054]),  .coef_in(coef[896]), .rdup_out(a7_wr[1038]), .rdlo_out(a7_wr[1054]));
			radix2 #(.width(width)) rd_st6_1039  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1039]), .rdlo_in(a6_wr[1055]),  .coef_in(coef[960]), .rdup_out(a7_wr[1039]), .rdlo_out(a7_wr[1055]));
			radix2 #(.width(width)) rd_st6_1056  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1056]), .rdlo_in(a6_wr[1072]),  .coef_in(coef[0]), .rdup_out(a7_wr[1056]), .rdlo_out(a7_wr[1072]));
			radix2 #(.width(width)) rd_st6_1057  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1057]), .rdlo_in(a6_wr[1073]),  .coef_in(coef[64]), .rdup_out(a7_wr[1057]), .rdlo_out(a7_wr[1073]));
			radix2 #(.width(width)) rd_st6_1058  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1058]), .rdlo_in(a6_wr[1074]),  .coef_in(coef[128]), .rdup_out(a7_wr[1058]), .rdlo_out(a7_wr[1074]));
			radix2 #(.width(width)) rd_st6_1059  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1059]), .rdlo_in(a6_wr[1075]),  .coef_in(coef[192]), .rdup_out(a7_wr[1059]), .rdlo_out(a7_wr[1075]));
			radix2 #(.width(width)) rd_st6_1060  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1060]), .rdlo_in(a6_wr[1076]),  .coef_in(coef[256]), .rdup_out(a7_wr[1060]), .rdlo_out(a7_wr[1076]));
			radix2 #(.width(width)) rd_st6_1061  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1061]), .rdlo_in(a6_wr[1077]),  .coef_in(coef[320]), .rdup_out(a7_wr[1061]), .rdlo_out(a7_wr[1077]));
			radix2 #(.width(width)) rd_st6_1062  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1062]), .rdlo_in(a6_wr[1078]),  .coef_in(coef[384]), .rdup_out(a7_wr[1062]), .rdlo_out(a7_wr[1078]));
			radix2 #(.width(width)) rd_st6_1063  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1063]), .rdlo_in(a6_wr[1079]),  .coef_in(coef[448]), .rdup_out(a7_wr[1063]), .rdlo_out(a7_wr[1079]));
			radix2 #(.width(width)) rd_st6_1064  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1064]), .rdlo_in(a6_wr[1080]),  .coef_in(coef[512]), .rdup_out(a7_wr[1064]), .rdlo_out(a7_wr[1080]));
			radix2 #(.width(width)) rd_st6_1065  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1065]), .rdlo_in(a6_wr[1081]),  .coef_in(coef[576]), .rdup_out(a7_wr[1065]), .rdlo_out(a7_wr[1081]));
			radix2 #(.width(width)) rd_st6_1066  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1066]), .rdlo_in(a6_wr[1082]),  .coef_in(coef[640]), .rdup_out(a7_wr[1066]), .rdlo_out(a7_wr[1082]));
			radix2 #(.width(width)) rd_st6_1067  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1067]), .rdlo_in(a6_wr[1083]),  .coef_in(coef[704]), .rdup_out(a7_wr[1067]), .rdlo_out(a7_wr[1083]));
			radix2 #(.width(width)) rd_st6_1068  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1068]), .rdlo_in(a6_wr[1084]),  .coef_in(coef[768]), .rdup_out(a7_wr[1068]), .rdlo_out(a7_wr[1084]));
			radix2 #(.width(width)) rd_st6_1069  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1069]), .rdlo_in(a6_wr[1085]),  .coef_in(coef[832]), .rdup_out(a7_wr[1069]), .rdlo_out(a7_wr[1085]));
			radix2 #(.width(width)) rd_st6_1070  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1070]), .rdlo_in(a6_wr[1086]),  .coef_in(coef[896]), .rdup_out(a7_wr[1070]), .rdlo_out(a7_wr[1086]));
			radix2 #(.width(width)) rd_st6_1071  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1071]), .rdlo_in(a6_wr[1087]),  .coef_in(coef[960]), .rdup_out(a7_wr[1071]), .rdlo_out(a7_wr[1087]));
			radix2 #(.width(width)) rd_st6_1088  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1088]), .rdlo_in(a6_wr[1104]),  .coef_in(coef[0]), .rdup_out(a7_wr[1088]), .rdlo_out(a7_wr[1104]));
			radix2 #(.width(width)) rd_st6_1089  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1089]), .rdlo_in(a6_wr[1105]),  .coef_in(coef[64]), .rdup_out(a7_wr[1089]), .rdlo_out(a7_wr[1105]));
			radix2 #(.width(width)) rd_st6_1090  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1090]), .rdlo_in(a6_wr[1106]),  .coef_in(coef[128]), .rdup_out(a7_wr[1090]), .rdlo_out(a7_wr[1106]));
			radix2 #(.width(width)) rd_st6_1091  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1091]), .rdlo_in(a6_wr[1107]),  .coef_in(coef[192]), .rdup_out(a7_wr[1091]), .rdlo_out(a7_wr[1107]));
			radix2 #(.width(width)) rd_st6_1092  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1092]), .rdlo_in(a6_wr[1108]),  .coef_in(coef[256]), .rdup_out(a7_wr[1092]), .rdlo_out(a7_wr[1108]));
			radix2 #(.width(width)) rd_st6_1093  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1093]), .rdlo_in(a6_wr[1109]),  .coef_in(coef[320]), .rdup_out(a7_wr[1093]), .rdlo_out(a7_wr[1109]));
			radix2 #(.width(width)) rd_st6_1094  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1094]), .rdlo_in(a6_wr[1110]),  .coef_in(coef[384]), .rdup_out(a7_wr[1094]), .rdlo_out(a7_wr[1110]));
			radix2 #(.width(width)) rd_st6_1095  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1095]), .rdlo_in(a6_wr[1111]),  .coef_in(coef[448]), .rdup_out(a7_wr[1095]), .rdlo_out(a7_wr[1111]));
			radix2 #(.width(width)) rd_st6_1096  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1096]), .rdlo_in(a6_wr[1112]),  .coef_in(coef[512]), .rdup_out(a7_wr[1096]), .rdlo_out(a7_wr[1112]));
			radix2 #(.width(width)) rd_st6_1097  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1097]), .rdlo_in(a6_wr[1113]),  .coef_in(coef[576]), .rdup_out(a7_wr[1097]), .rdlo_out(a7_wr[1113]));
			radix2 #(.width(width)) rd_st6_1098  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1098]), .rdlo_in(a6_wr[1114]),  .coef_in(coef[640]), .rdup_out(a7_wr[1098]), .rdlo_out(a7_wr[1114]));
			radix2 #(.width(width)) rd_st6_1099  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1099]), .rdlo_in(a6_wr[1115]),  .coef_in(coef[704]), .rdup_out(a7_wr[1099]), .rdlo_out(a7_wr[1115]));
			radix2 #(.width(width)) rd_st6_1100  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1100]), .rdlo_in(a6_wr[1116]),  .coef_in(coef[768]), .rdup_out(a7_wr[1100]), .rdlo_out(a7_wr[1116]));
			radix2 #(.width(width)) rd_st6_1101  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1101]), .rdlo_in(a6_wr[1117]),  .coef_in(coef[832]), .rdup_out(a7_wr[1101]), .rdlo_out(a7_wr[1117]));
			radix2 #(.width(width)) rd_st6_1102  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1102]), .rdlo_in(a6_wr[1118]),  .coef_in(coef[896]), .rdup_out(a7_wr[1102]), .rdlo_out(a7_wr[1118]));
			radix2 #(.width(width)) rd_st6_1103  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1103]), .rdlo_in(a6_wr[1119]),  .coef_in(coef[960]), .rdup_out(a7_wr[1103]), .rdlo_out(a7_wr[1119]));
			radix2 #(.width(width)) rd_st6_1120  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1120]), .rdlo_in(a6_wr[1136]),  .coef_in(coef[0]), .rdup_out(a7_wr[1120]), .rdlo_out(a7_wr[1136]));
			radix2 #(.width(width)) rd_st6_1121  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1121]), .rdlo_in(a6_wr[1137]),  .coef_in(coef[64]), .rdup_out(a7_wr[1121]), .rdlo_out(a7_wr[1137]));
			radix2 #(.width(width)) rd_st6_1122  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1122]), .rdlo_in(a6_wr[1138]),  .coef_in(coef[128]), .rdup_out(a7_wr[1122]), .rdlo_out(a7_wr[1138]));
			radix2 #(.width(width)) rd_st6_1123  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1123]), .rdlo_in(a6_wr[1139]),  .coef_in(coef[192]), .rdup_out(a7_wr[1123]), .rdlo_out(a7_wr[1139]));
			radix2 #(.width(width)) rd_st6_1124  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1124]), .rdlo_in(a6_wr[1140]),  .coef_in(coef[256]), .rdup_out(a7_wr[1124]), .rdlo_out(a7_wr[1140]));
			radix2 #(.width(width)) rd_st6_1125  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1125]), .rdlo_in(a6_wr[1141]),  .coef_in(coef[320]), .rdup_out(a7_wr[1125]), .rdlo_out(a7_wr[1141]));
			radix2 #(.width(width)) rd_st6_1126  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1126]), .rdlo_in(a6_wr[1142]),  .coef_in(coef[384]), .rdup_out(a7_wr[1126]), .rdlo_out(a7_wr[1142]));
			radix2 #(.width(width)) rd_st6_1127  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1127]), .rdlo_in(a6_wr[1143]),  .coef_in(coef[448]), .rdup_out(a7_wr[1127]), .rdlo_out(a7_wr[1143]));
			radix2 #(.width(width)) rd_st6_1128  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1128]), .rdlo_in(a6_wr[1144]),  .coef_in(coef[512]), .rdup_out(a7_wr[1128]), .rdlo_out(a7_wr[1144]));
			radix2 #(.width(width)) rd_st6_1129  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1129]), .rdlo_in(a6_wr[1145]),  .coef_in(coef[576]), .rdup_out(a7_wr[1129]), .rdlo_out(a7_wr[1145]));
			radix2 #(.width(width)) rd_st6_1130  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1130]), .rdlo_in(a6_wr[1146]),  .coef_in(coef[640]), .rdup_out(a7_wr[1130]), .rdlo_out(a7_wr[1146]));
			radix2 #(.width(width)) rd_st6_1131  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1131]), .rdlo_in(a6_wr[1147]),  .coef_in(coef[704]), .rdup_out(a7_wr[1131]), .rdlo_out(a7_wr[1147]));
			radix2 #(.width(width)) rd_st6_1132  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1132]), .rdlo_in(a6_wr[1148]),  .coef_in(coef[768]), .rdup_out(a7_wr[1132]), .rdlo_out(a7_wr[1148]));
			radix2 #(.width(width)) rd_st6_1133  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1133]), .rdlo_in(a6_wr[1149]),  .coef_in(coef[832]), .rdup_out(a7_wr[1133]), .rdlo_out(a7_wr[1149]));
			radix2 #(.width(width)) rd_st6_1134  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1134]), .rdlo_in(a6_wr[1150]),  .coef_in(coef[896]), .rdup_out(a7_wr[1134]), .rdlo_out(a7_wr[1150]));
			radix2 #(.width(width)) rd_st6_1135  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1135]), .rdlo_in(a6_wr[1151]),  .coef_in(coef[960]), .rdup_out(a7_wr[1135]), .rdlo_out(a7_wr[1151]));
			radix2 #(.width(width)) rd_st6_1152  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1152]), .rdlo_in(a6_wr[1168]),  .coef_in(coef[0]), .rdup_out(a7_wr[1152]), .rdlo_out(a7_wr[1168]));
			radix2 #(.width(width)) rd_st6_1153  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1153]), .rdlo_in(a6_wr[1169]),  .coef_in(coef[64]), .rdup_out(a7_wr[1153]), .rdlo_out(a7_wr[1169]));
			radix2 #(.width(width)) rd_st6_1154  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1154]), .rdlo_in(a6_wr[1170]),  .coef_in(coef[128]), .rdup_out(a7_wr[1154]), .rdlo_out(a7_wr[1170]));
			radix2 #(.width(width)) rd_st6_1155  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1155]), .rdlo_in(a6_wr[1171]),  .coef_in(coef[192]), .rdup_out(a7_wr[1155]), .rdlo_out(a7_wr[1171]));
			radix2 #(.width(width)) rd_st6_1156  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1156]), .rdlo_in(a6_wr[1172]),  .coef_in(coef[256]), .rdup_out(a7_wr[1156]), .rdlo_out(a7_wr[1172]));
			radix2 #(.width(width)) rd_st6_1157  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1157]), .rdlo_in(a6_wr[1173]),  .coef_in(coef[320]), .rdup_out(a7_wr[1157]), .rdlo_out(a7_wr[1173]));
			radix2 #(.width(width)) rd_st6_1158  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1158]), .rdlo_in(a6_wr[1174]),  .coef_in(coef[384]), .rdup_out(a7_wr[1158]), .rdlo_out(a7_wr[1174]));
			radix2 #(.width(width)) rd_st6_1159  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1159]), .rdlo_in(a6_wr[1175]),  .coef_in(coef[448]), .rdup_out(a7_wr[1159]), .rdlo_out(a7_wr[1175]));
			radix2 #(.width(width)) rd_st6_1160  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1160]), .rdlo_in(a6_wr[1176]),  .coef_in(coef[512]), .rdup_out(a7_wr[1160]), .rdlo_out(a7_wr[1176]));
			radix2 #(.width(width)) rd_st6_1161  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1161]), .rdlo_in(a6_wr[1177]),  .coef_in(coef[576]), .rdup_out(a7_wr[1161]), .rdlo_out(a7_wr[1177]));
			radix2 #(.width(width)) rd_st6_1162  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1162]), .rdlo_in(a6_wr[1178]),  .coef_in(coef[640]), .rdup_out(a7_wr[1162]), .rdlo_out(a7_wr[1178]));
			radix2 #(.width(width)) rd_st6_1163  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1163]), .rdlo_in(a6_wr[1179]),  .coef_in(coef[704]), .rdup_out(a7_wr[1163]), .rdlo_out(a7_wr[1179]));
			radix2 #(.width(width)) rd_st6_1164  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1164]), .rdlo_in(a6_wr[1180]),  .coef_in(coef[768]), .rdup_out(a7_wr[1164]), .rdlo_out(a7_wr[1180]));
			radix2 #(.width(width)) rd_st6_1165  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1165]), .rdlo_in(a6_wr[1181]),  .coef_in(coef[832]), .rdup_out(a7_wr[1165]), .rdlo_out(a7_wr[1181]));
			radix2 #(.width(width)) rd_st6_1166  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1166]), .rdlo_in(a6_wr[1182]),  .coef_in(coef[896]), .rdup_out(a7_wr[1166]), .rdlo_out(a7_wr[1182]));
			radix2 #(.width(width)) rd_st6_1167  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1167]), .rdlo_in(a6_wr[1183]),  .coef_in(coef[960]), .rdup_out(a7_wr[1167]), .rdlo_out(a7_wr[1183]));
			radix2 #(.width(width)) rd_st6_1184  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1184]), .rdlo_in(a6_wr[1200]),  .coef_in(coef[0]), .rdup_out(a7_wr[1184]), .rdlo_out(a7_wr[1200]));
			radix2 #(.width(width)) rd_st6_1185  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1185]), .rdlo_in(a6_wr[1201]),  .coef_in(coef[64]), .rdup_out(a7_wr[1185]), .rdlo_out(a7_wr[1201]));
			radix2 #(.width(width)) rd_st6_1186  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1186]), .rdlo_in(a6_wr[1202]),  .coef_in(coef[128]), .rdup_out(a7_wr[1186]), .rdlo_out(a7_wr[1202]));
			radix2 #(.width(width)) rd_st6_1187  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1187]), .rdlo_in(a6_wr[1203]),  .coef_in(coef[192]), .rdup_out(a7_wr[1187]), .rdlo_out(a7_wr[1203]));
			radix2 #(.width(width)) rd_st6_1188  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1188]), .rdlo_in(a6_wr[1204]),  .coef_in(coef[256]), .rdup_out(a7_wr[1188]), .rdlo_out(a7_wr[1204]));
			radix2 #(.width(width)) rd_st6_1189  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1189]), .rdlo_in(a6_wr[1205]),  .coef_in(coef[320]), .rdup_out(a7_wr[1189]), .rdlo_out(a7_wr[1205]));
			radix2 #(.width(width)) rd_st6_1190  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1190]), .rdlo_in(a6_wr[1206]),  .coef_in(coef[384]), .rdup_out(a7_wr[1190]), .rdlo_out(a7_wr[1206]));
			radix2 #(.width(width)) rd_st6_1191  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1191]), .rdlo_in(a6_wr[1207]),  .coef_in(coef[448]), .rdup_out(a7_wr[1191]), .rdlo_out(a7_wr[1207]));
			radix2 #(.width(width)) rd_st6_1192  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1192]), .rdlo_in(a6_wr[1208]),  .coef_in(coef[512]), .rdup_out(a7_wr[1192]), .rdlo_out(a7_wr[1208]));
			radix2 #(.width(width)) rd_st6_1193  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1193]), .rdlo_in(a6_wr[1209]),  .coef_in(coef[576]), .rdup_out(a7_wr[1193]), .rdlo_out(a7_wr[1209]));
			radix2 #(.width(width)) rd_st6_1194  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1194]), .rdlo_in(a6_wr[1210]),  .coef_in(coef[640]), .rdup_out(a7_wr[1194]), .rdlo_out(a7_wr[1210]));
			radix2 #(.width(width)) rd_st6_1195  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1195]), .rdlo_in(a6_wr[1211]),  .coef_in(coef[704]), .rdup_out(a7_wr[1195]), .rdlo_out(a7_wr[1211]));
			radix2 #(.width(width)) rd_st6_1196  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1196]), .rdlo_in(a6_wr[1212]),  .coef_in(coef[768]), .rdup_out(a7_wr[1196]), .rdlo_out(a7_wr[1212]));
			radix2 #(.width(width)) rd_st6_1197  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1197]), .rdlo_in(a6_wr[1213]),  .coef_in(coef[832]), .rdup_out(a7_wr[1197]), .rdlo_out(a7_wr[1213]));
			radix2 #(.width(width)) rd_st6_1198  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1198]), .rdlo_in(a6_wr[1214]),  .coef_in(coef[896]), .rdup_out(a7_wr[1198]), .rdlo_out(a7_wr[1214]));
			radix2 #(.width(width)) rd_st6_1199  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1199]), .rdlo_in(a6_wr[1215]),  .coef_in(coef[960]), .rdup_out(a7_wr[1199]), .rdlo_out(a7_wr[1215]));
			radix2 #(.width(width)) rd_st6_1216  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1216]), .rdlo_in(a6_wr[1232]),  .coef_in(coef[0]), .rdup_out(a7_wr[1216]), .rdlo_out(a7_wr[1232]));
			radix2 #(.width(width)) rd_st6_1217  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1217]), .rdlo_in(a6_wr[1233]),  .coef_in(coef[64]), .rdup_out(a7_wr[1217]), .rdlo_out(a7_wr[1233]));
			radix2 #(.width(width)) rd_st6_1218  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1218]), .rdlo_in(a6_wr[1234]),  .coef_in(coef[128]), .rdup_out(a7_wr[1218]), .rdlo_out(a7_wr[1234]));
			radix2 #(.width(width)) rd_st6_1219  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1219]), .rdlo_in(a6_wr[1235]),  .coef_in(coef[192]), .rdup_out(a7_wr[1219]), .rdlo_out(a7_wr[1235]));
			radix2 #(.width(width)) rd_st6_1220  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1220]), .rdlo_in(a6_wr[1236]),  .coef_in(coef[256]), .rdup_out(a7_wr[1220]), .rdlo_out(a7_wr[1236]));
			radix2 #(.width(width)) rd_st6_1221  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1221]), .rdlo_in(a6_wr[1237]),  .coef_in(coef[320]), .rdup_out(a7_wr[1221]), .rdlo_out(a7_wr[1237]));
			radix2 #(.width(width)) rd_st6_1222  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1222]), .rdlo_in(a6_wr[1238]),  .coef_in(coef[384]), .rdup_out(a7_wr[1222]), .rdlo_out(a7_wr[1238]));
			radix2 #(.width(width)) rd_st6_1223  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1223]), .rdlo_in(a6_wr[1239]),  .coef_in(coef[448]), .rdup_out(a7_wr[1223]), .rdlo_out(a7_wr[1239]));
			radix2 #(.width(width)) rd_st6_1224  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1224]), .rdlo_in(a6_wr[1240]),  .coef_in(coef[512]), .rdup_out(a7_wr[1224]), .rdlo_out(a7_wr[1240]));
			radix2 #(.width(width)) rd_st6_1225  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1225]), .rdlo_in(a6_wr[1241]),  .coef_in(coef[576]), .rdup_out(a7_wr[1225]), .rdlo_out(a7_wr[1241]));
			radix2 #(.width(width)) rd_st6_1226  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1226]), .rdlo_in(a6_wr[1242]),  .coef_in(coef[640]), .rdup_out(a7_wr[1226]), .rdlo_out(a7_wr[1242]));
			radix2 #(.width(width)) rd_st6_1227  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1227]), .rdlo_in(a6_wr[1243]),  .coef_in(coef[704]), .rdup_out(a7_wr[1227]), .rdlo_out(a7_wr[1243]));
			radix2 #(.width(width)) rd_st6_1228  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1228]), .rdlo_in(a6_wr[1244]),  .coef_in(coef[768]), .rdup_out(a7_wr[1228]), .rdlo_out(a7_wr[1244]));
			radix2 #(.width(width)) rd_st6_1229  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1229]), .rdlo_in(a6_wr[1245]),  .coef_in(coef[832]), .rdup_out(a7_wr[1229]), .rdlo_out(a7_wr[1245]));
			radix2 #(.width(width)) rd_st6_1230  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1230]), .rdlo_in(a6_wr[1246]),  .coef_in(coef[896]), .rdup_out(a7_wr[1230]), .rdlo_out(a7_wr[1246]));
			radix2 #(.width(width)) rd_st6_1231  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1231]), .rdlo_in(a6_wr[1247]),  .coef_in(coef[960]), .rdup_out(a7_wr[1231]), .rdlo_out(a7_wr[1247]));
			radix2 #(.width(width)) rd_st6_1248  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1248]), .rdlo_in(a6_wr[1264]),  .coef_in(coef[0]), .rdup_out(a7_wr[1248]), .rdlo_out(a7_wr[1264]));
			radix2 #(.width(width)) rd_st6_1249  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1249]), .rdlo_in(a6_wr[1265]),  .coef_in(coef[64]), .rdup_out(a7_wr[1249]), .rdlo_out(a7_wr[1265]));
			radix2 #(.width(width)) rd_st6_1250  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1250]), .rdlo_in(a6_wr[1266]),  .coef_in(coef[128]), .rdup_out(a7_wr[1250]), .rdlo_out(a7_wr[1266]));
			radix2 #(.width(width)) rd_st6_1251  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1251]), .rdlo_in(a6_wr[1267]),  .coef_in(coef[192]), .rdup_out(a7_wr[1251]), .rdlo_out(a7_wr[1267]));
			radix2 #(.width(width)) rd_st6_1252  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1252]), .rdlo_in(a6_wr[1268]),  .coef_in(coef[256]), .rdup_out(a7_wr[1252]), .rdlo_out(a7_wr[1268]));
			radix2 #(.width(width)) rd_st6_1253  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1253]), .rdlo_in(a6_wr[1269]),  .coef_in(coef[320]), .rdup_out(a7_wr[1253]), .rdlo_out(a7_wr[1269]));
			radix2 #(.width(width)) rd_st6_1254  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1254]), .rdlo_in(a6_wr[1270]),  .coef_in(coef[384]), .rdup_out(a7_wr[1254]), .rdlo_out(a7_wr[1270]));
			radix2 #(.width(width)) rd_st6_1255  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1255]), .rdlo_in(a6_wr[1271]),  .coef_in(coef[448]), .rdup_out(a7_wr[1255]), .rdlo_out(a7_wr[1271]));
			radix2 #(.width(width)) rd_st6_1256  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1256]), .rdlo_in(a6_wr[1272]),  .coef_in(coef[512]), .rdup_out(a7_wr[1256]), .rdlo_out(a7_wr[1272]));
			radix2 #(.width(width)) rd_st6_1257  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1257]), .rdlo_in(a6_wr[1273]),  .coef_in(coef[576]), .rdup_out(a7_wr[1257]), .rdlo_out(a7_wr[1273]));
			radix2 #(.width(width)) rd_st6_1258  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1258]), .rdlo_in(a6_wr[1274]),  .coef_in(coef[640]), .rdup_out(a7_wr[1258]), .rdlo_out(a7_wr[1274]));
			radix2 #(.width(width)) rd_st6_1259  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1259]), .rdlo_in(a6_wr[1275]),  .coef_in(coef[704]), .rdup_out(a7_wr[1259]), .rdlo_out(a7_wr[1275]));
			radix2 #(.width(width)) rd_st6_1260  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1260]), .rdlo_in(a6_wr[1276]),  .coef_in(coef[768]), .rdup_out(a7_wr[1260]), .rdlo_out(a7_wr[1276]));
			radix2 #(.width(width)) rd_st6_1261  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1261]), .rdlo_in(a6_wr[1277]),  .coef_in(coef[832]), .rdup_out(a7_wr[1261]), .rdlo_out(a7_wr[1277]));
			radix2 #(.width(width)) rd_st6_1262  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1262]), .rdlo_in(a6_wr[1278]),  .coef_in(coef[896]), .rdup_out(a7_wr[1262]), .rdlo_out(a7_wr[1278]));
			radix2 #(.width(width)) rd_st6_1263  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1263]), .rdlo_in(a6_wr[1279]),  .coef_in(coef[960]), .rdup_out(a7_wr[1263]), .rdlo_out(a7_wr[1279]));
			radix2 #(.width(width)) rd_st6_1280  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1280]), .rdlo_in(a6_wr[1296]),  .coef_in(coef[0]), .rdup_out(a7_wr[1280]), .rdlo_out(a7_wr[1296]));
			radix2 #(.width(width)) rd_st6_1281  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1281]), .rdlo_in(a6_wr[1297]),  .coef_in(coef[64]), .rdup_out(a7_wr[1281]), .rdlo_out(a7_wr[1297]));
			radix2 #(.width(width)) rd_st6_1282  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1282]), .rdlo_in(a6_wr[1298]),  .coef_in(coef[128]), .rdup_out(a7_wr[1282]), .rdlo_out(a7_wr[1298]));
			radix2 #(.width(width)) rd_st6_1283  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1283]), .rdlo_in(a6_wr[1299]),  .coef_in(coef[192]), .rdup_out(a7_wr[1283]), .rdlo_out(a7_wr[1299]));
			radix2 #(.width(width)) rd_st6_1284  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1284]), .rdlo_in(a6_wr[1300]),  .coef_in(coef[256]), .rdup_out(a7_wr[1284]), .rdlo_out(a7_wr[1300]));
			radix2 #(.width(width)) rd_st6_1285  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1285]), .rdlo_in(a6_wr[1301]),  .coef_in(coef[320]), .rdup_out(a7_wr[1285]), .rdlo_out(a7_wr[1301]));
			radix2 #(.width(width)) rd_st6_1286  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1286]), .rdlo_in(a6_wr[1302]),  .coef_in(coef[384]), .rdup_out(a7_wr[1286]), .rdlo_out(a7_wr[1302]));
			radix2 #(.width(width)) rd_st6_1287  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1287]), .rdlo_in(a6_wr[1303]),  .coef_in(coef[448]), .rdup_out(a7_wr[1287]), .rdlo_out(a7_wr[1303]));
			radix2 #(.width(width)) rd_st6_1288  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1288]), .rdlo_in(a6_wr[1304]),  .coef_in(coef[512]), .rdup_out(a7_wr[1288]), .rdlo_out(a7_wr[1304]));
			radix2 #(.width(width)) rd_st6_1289  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1289]), .rdlo_in(a6_wr[1305]),  .coef_in(coef[576]), .rdup_out(a7_wr[1289]), .rdlo_out(a7_wr[1305]));
			radix2 #(.width(width)) rd_st6_1290  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1290]), .rdlo_in(a6_wr[1306]),  .coef_in(coef[640]), .rdup_out(a7_wr[1290]), .rdlo_out(a7_wr[1306]));
			radix2 #(.width(width)) rd_st6_1291  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1291]), .rdlo_in(a6_wr[1307]),  .coef_in(coef[704]), .rdup_out(a7_wr[1291]), .rdlo_out(a7_wr[1307]));
			radix2 #(.width(width)) rd_st6_1292  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1292]), .rdlo_in(a6_wr[1308]),  .coef_in(coef[768]), .rdup_out(a7_wr[1292]), .rdlo_out(a7_wr[1308]));
			radix2 #(.width(width)) rd_st6_1293  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1293]), .rdlo_in(a6_wr[1309]),  .coef_in(coef[832]), .rdup_out(a7_wr[1293]), .rdlo_out(a7_wr[1309]));
			radix2 #(.width(width)) rd_st6_1294  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1294]), .rdlo_in(a6_wr[1310]),  .coef_in(coef[896]), .rdup_out(a7_wr[1294]), .rdlo_out(a7_wr[1310]));
			radix2 #(.width(width)) rd_st6_1295  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1295]), .rdlo_in(a6_wr[1311]),  .coef_in(coef[960]), .rdup_out(a7_wr[1295]), .rdlo_out(a7_wr[1311]));
			radix2 #(.width(width)) rd_st6_1312  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1312]), .rdlo_in(a6_wr[1328]),  .coef_in(coef[0]), .rdup_out(a7_wr[1312]), .rdlo_out(a7_wr[1328]));
			radix2 #(.width(width)) rd_st6_1313  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1313]), .rdlo_in(a6_wr[1329]),  .coef_in(coef[64]), .rdup_out(a7_wr[1313]), .rdlo_out(a7_wr[1329]));
			radix2 #(.width(width)) rd_st6_1314  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1314]), .rdlo_in(a6_wr[1330]),  .coef_in(coef[128]), .rdup_out(a7_wr[1314]), .rdlo_out(a7_wr[1330]));
			radix2 #(.width(width)) rd_st6_1315  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1315]), .rdlo_in(a6_wr[1331]),  .coef_in(coef[192]), .rdup_out(a7_wr[1315]), .rdlo_out(a7_wr[1331]));
			radix2 #(.width(width)) rd_st6_1316  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1316]), .rdlo_in(a6_wr[1332]),  .coef_in(coef[256]), .rdup_out(a7_wr[1316]), .rdlo_out(a7_wr[1332]));
			radix2 #(.width(width)) rd_st6_1317  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1317]), .rdlo_in(a6_wr[1333]),  .coef_in(coef[320]), .rdup_out(a7_wr[1317]), .rdlo_out(a7_wr[1333]));
			radix2 #(.width(width)) rd_st6_1318  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1318]), .rdlo_in(a6_wr[1334]),  .coef_in(coef[384]), .rdup_out(a7_wr[1318]), .rdlo_out(a7_wr[1334]));
			radix2 #(.width(width)) rd_st6_1319  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1319]), .rdlo_in(a6_wr[1335]),  .coef_in(coef[448]), .rdup_out(a7_wr[1319]), .rdlo_out(a7_wr[1335]));
			radix2 #(.width(width)) rd_st6_1320  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1320]), .rdlo_in(a6_wr[1336]),  .coef_in(coef[512]), .rdup_out(a7_wr[1320]), .rdlo_out(a7_wr[1336]));
			radix2 #(.width(width)) rd_st6_1321  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1321]), .rdlo_in(a6_wr[1337]),  .coef_in(coef[576]), .rdup_out(a7_wr[1321]), .rdlo_out(a7_wr[1337]));
			radix2 #(.width(width)) rd_st6_1322  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1322]), .rdlo_in(a6_wr[1338]),  .coef_in(coef[640]), .rdup_out(a7_wr[1322]), .rdlo_out(a7_wr[1338]));
			radix2 #(.width(width)) rd_st6_1323  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1323]), .rdlo_in(a6_wr[1339]),  .coef_in(coef[704]), .rdup_out(a7_wr[1323]), .rdlo_out(a7_wr[1339]));
			radix2 #(.width(width)) rd_st6_1324  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1324]), .rdlo_in(a6_wr[1340]),  .coef_in(coef[768]), .rdup_out(a7_wr[1324]), .rdlo_out(a7_wr[1340]));
			radix2 #(.width(width)) rd_st6_1325  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1325]), .rdlo_in(a6_wr[1341]),  .coef_in(coef[832]), .rdup_out(a7_wr[1325]), .rdlo_out(a7_wr[1341]));
			radix2 #(.width(width)) rd_st6_1326  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1326]), .rdlo_in(a6_wr[1342]),  .coef_in(coef[896]), .rdup_out(a7_wr[1326]), .rdlo_out(a7_wr[1342]));
			radix2 #(.width(width)) rd_st6_1327  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1327]), .rdlo_in(a6_wr[1343]),  .coef_in(coef[960]), .rdup_out(a7_wr[1327]), .rdlo_out(a7_wr[1343]));
			radix2 #(.width(width)) rd_st6_1344  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1344]), .rdlo_in(a6_wr[1360]),  .coef_in(coef[0]), .rdup_out(a7_wr[1344]), .rdlo_out(a7_wr[1360]));
			radix2 #(.width(width)) rd_st6_1345  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1345]), .rdlo_in(a6_wr[1361]),  .coef_in(coef[64]), .rdup_out(a7_wr[1345]), .rdlo_out(a7_wr[1361]));
			radix2 #(.width(width)) rd_st6_1346  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1346]), .rdlo_in(a6_wr[1362]),  .coef_in(coef[128]), .rdup_out(a7_wr[1346]), .rdlo_out(a7_wr[1362]));
			radix2 #(.width(width)) rd_st6_1347  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1347]), .rdlo_in(a6_wr[1363]),  .coef_in(coef[192]), .rdup_out(a7_wr[1347]), .rdlo_out(a7_wr[1363]));
			radix2 #(.width(width)) rd_st6_1348  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1348]), .rdlo_in(a6_wr[1364]),  .coef_in(coef[256]), .rdup_out(a7_wr[1348]), .rdlo_out(a7_wr[1364]));
			radix2 #(.width(width)) rd_st6_1349  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1349]), .rdlo_in(a6_wr[1365]),  .coef_in(coef[320]), .rdup_out(a7_wr[1349]), .rdlo_out(a7_wr[1365]));
			radix2 #(.width(width)) rd_st6_1350  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1350]), .rdlo_in(a6_wr[1366]),  .coef_in(coef[384]), .rdup_out(a7_wr[1350]), .rdlo_out(a7_wr[1366]));
			radix2 #(.width(width)) rd_st6_1351  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1351]), .rdlo_in(a6_wr[1367]),  .coef_in(coef[448]), .rdup_out(a7_wr[1351]), .rdlo_out(a7_wr[1367]));
			radix2 #(.width(width)) rd_st6_1352  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1352]), .rdlo_in(a6_wr[1368]),  .coef_in(coef[512]), .rdup_out(a7_wr[1352]), .rdlo_out(a7_wr[1368]));
			radix2 #(.width(width)) rd_st6_1353  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1353]), .rdlo_in(a6_wr[1369]),  .coef_in(coef[576]), .rdup_out(a7_wr[1353]), .rdlo_out(a7_wr[1369]));
			radix2 #(.width(width)) rd_st6_1354  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1354]), .rdlo_in(a6_wr[1370]),  .coef_in(coef[640]), .rdup_out(a7_wr[1354]), .rdlo_out(a7_wr[1370]));
			radix2 #(.width(width)) rd_st6_1355  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1355]), .rdlo_in(a6_wr[1371]),  .coef_in(coef[704]), .rdup_out(a7_wr[1355]), .rdlo_out(a7_wr[1371]));
			radix2 #(.width(width)) rd_st6_1356  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1356]), .rdlo_in(a6_wr[1372]),  .coef_in(coef[768]), .rdup_out(a7_wr[1356]), .rdlo_out(a7_wr[1372]));
			radix2 #(.width(width)) rd_st6_1357  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1357]), .rdlo_in(a6_wr[1373]),  .coef_in(coef[832]), .rdup_out(a7_wr[1357]), .rdlo_out(a7_wr[1373]));
			radix2 #(.width(width)) rd_st6_1358  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1358]), .rdlo_in(a6_wr[1374]),  .coef_in(coef[896]), .rdup_out(a7_wr[1358]), .rdlo_out(a7_wr[1374]));
			radix2 #(.width(width)) rd_st6_1359  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1359]), .rdlo_in(a6_wr[1375]),  .coef_in(coef[960]), .rdup_out(a7_wr[1359]), .rdlo_out(a7_wr[1375]));
			radix2 #(.width(width)) rd_st6_1376  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1376]), .rdlo_in(a6_wr[1392]),  .coef_in(coef[0]), .rdup_out(a7_wr[1376]), .rdlo_out(a7_wr[1392]));
			radix2 #(.width(width)) rd_st6_1377  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1377]), .rdlo_in(a6_wr[1393]),  .coef_in(coef[64]), .rdup_out(a7_wr[1377]), .rdlo_out(a7_wr[1393]));
			radix2 #(.width(width)) rd_st6_1378  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1378]), .rdlo_in(a6_wr[1394]),  .coef_in(coef[128]), .rdup_out(a7_wr[1378]), .rdlo_out(a7_wr[1394]));
			radix2 #(.width(width)) rd_st6_1379  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1379]), .rdlo_in(a6_wr[1395]),  .coef_in(coef[192]), .rdup_out(a7_wr[1379]), .rdlo_out(a7_wr[1395]));
			radix2 #(.width(width)) rd_st6_1380  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1380]), .rdlo_in(a6_wr[1396]),  .coef_in(coef[256]), .rdup_out(a7_wr[1380]), .rdlo_out(a7_wr[1396]));
			radix2 #(.width(width)) rd_st6_1381  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1381]), .rdlo_in(a6_wr[1397]),  .coef_in(coef[320]), .rdup_out(a7_wr[1381]), .rdlo_out(a7_wr[1397]));
			radix2 #(.width(width)) rd_st6_1382  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1382]), .rdlo_in(a6_wr[1398]),  .coef_in(coef[384]), .rdup_out(a7_wr[1382]), .rdlo_out(a7_wr[1398]));
			radix2 #(.width(width)) rd_st6_1383  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1383]), .rdlo_in(a6_wr[1399]),  .coef_in(coef[448]), .rdup_out(a7_wr[1383]), .rdlo_out(a7_wr[1399]));
			radix2 #(.width(width)) rd_st6_1384  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1384]), .rdlo_in(a6_wr[1400]),  .coef_in(coef[512]), .rdup_out(a7_wr[1384]), .rdlo_out(a7_wr[1400]));
			radix2 #(.width(width)) rd_st6_1385  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1385]), .rdlo_in(a6_wr[1401]),  .coef_in(coef[576]), .rdup_out(a7_wr[1385]), .rdlo_out(a7_wr[1401]));
			radix2 #(.width(width)) rd_st6_1386  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1386]), .rdlo_in(a6_wr[1402]),  .coef_in(coef[640]), .rdup_out(a7_wr[1386]), .rdlo_out(a7_wr[1402]));
			radix2 #(.width(width)) rd_st6_1387  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1387]), .rdlo_in(a6_wr[1403]),  .coef_in(coef[704]), .rdup_out(a7_wr[1387]), .rdlo_out(a7_wr[1403]));
			radix2 #(.width(width)) rd_st6_1388  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1388]), .rdlo_in(a6_wr[1404]),  .coef_in(coef[768]), .rdup_out(a7_wr[1388]), .rdlo_out(a7_wr[1404]));
			radix2 #(.width(width)) rd_st6_1389  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1389]), .rdlo_in(a6_wr[1405]),  .coef_in(coef[832]), .rdup_out(a7_wr[1389]), .rdlo_out(a7_wr[1405]));
			radix2 #(.width(width)) rd_st6_1390  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1390]), .rdlo_in(a6_wr[1406]),  .coef_in(coef[896]), .rdup_out(a7_wr[1390]), .rdlo_out(a7_wr[1406]));
			radix2 #(.width(width)) rd_st6_1391  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1391]), .rdlo_in(a6_wr[1407]),  .coef_in(coef[960]), .rdup_out(a7_wr[1391]), .rdlo_out(a7_wr[1407]));
			radix2 #(.width(width)) rd_st6_1408  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1408]), .rdlo_in(a6_wr[1424]),  .coef_in(coef[0]), .rdup_out(a7_wr[1408]), .rdlo_out(a7_wr[1424]));
			radix2 #(.width(width)) rd_st6_1409  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1409]), .rdlo_in(a6_wr[1425]),  .coef_in(coef[64]), .rdup_out(a7_wr[1409]), .rdlo_out(a7_wr[1425]));
			radix2 #(.width(width)) rd_st6_1410  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1410]), .rdlo_in(a6_wr[1426]),  .coef_in(coef[128]), .rdup_out(a7_wr[1410]), .rdlo_out(a7_wr[1426]));
			radix2 #(.width(width)) rd_st6_1411  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1411]), .rdlo_in(a6_wr[1427]),  .coef_in(coef[192]), .rdup_out(a7_wr[1411]), .rdlo_out(a7_wr[1427]));
			radix2 #(.width(width)) rd_st6_1412  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1412]), .rdlo_in(a6_wr[1428]),  .coef_in(coef[256]), .rdup_out(a7_wr[1412]), .rdlo_out(a7_wr[1428]));
			radix2 #(.width(width)) rd_st6_1413  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1413]), .rdlo_in(a6_wr[1429]),  .coef_in(coef[320]), .rdup_out(a7_wr[1413]), .rdlo_out(a7_wr[1429]));
			radix2 #(.width(width)) rd_st6_1414  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1414]), .rdlo_in(a6_wr[1430]),  .coef_in(coef[384]), .rdup_out(a7_wr[1414]), .rdlo_out(a7_wr[1430]));
			radix2 #(.width(width)) rd_st6_1415  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1415]), .rdlo_in(a6_wr[1431]),  .coef_in(coef[448]), .rdup_out(a7_wr[1415]), .rdlo_out(a7_wr[1431]));
			radix2 #(.width(width)) rd_st6_1416  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1416]), .rdlo_in(a6_wr[1432]),  .coef_in(coef[512]), .rdup_out(a7_wr[1416]), .rdlo_out(a7_wr[1432]));
			radix2 #(.width(width)) rd_st6_1417  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1417]), .rdlo_in(a6_wr[1433]),  .coef_in(coef[576]), .rdup_out(a7_wr[1417]), .rdlo_out(a7_wr[1433]));
			radix2 #(.width(width)) rd_st6_1418  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1418]), .rdlo_in(a6_wr[1434]),  .coef_in(coef[640]), .rdup_out(a7_wr[1418]), .rdlo_out(a7_wr[1434]));
			radix2 #(.width(width)) rd_st6_1419  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1419]), .rdlo_in(a6_wr[1435]),  .coef_in(coef[704]), .rdup_out(a7_wr[1419]), .rdlo_out(a7_wr[1435]));
			radix2 #(.width(width)) rd_st6_1420  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1420]), .rdlo_in(a6_wr[1436]),  .coef_in(coef[768]), .rdup_out(a7_wr[1420]), .rdlo_out(a7_wr[1436]));
			radix2 #(.width(width)) rd_st6_1421  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1421]), .rdlo_in(a6_wr[1437]),  .coef_in(coef[832]), .rdup_out(a7_wr[1421]), .rdlo_out(a7_wr[1437]));
			radix2 #(.width(width)) rd_st6_1422  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1422]), .rdlo_in(a6_wr[1438]),  .coef_in(coef[896]), .rdup_out(a7_wr[1422]), .rdlo_out(a7_wr[1438]));
			radix2 #(.width(width)) rd_st6_1423  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1423]), .rdlo_in(a6_wr[1439]),  .coef_in(coef[960]), .rdup_out(a7_wr[1423]), .rdlo_out(a7_wr[1439]));
			radix2 #(.width(width)) rd_st6_1440  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1440]), .rdlo_in(a6_wr[1456]),  .coef_in(coef[0]), .rdup_out(a7_wr[1440]), .rdlo_out(a7_wr[1456]));
			radix2 #(.width(width)) rd_st6_1441  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1441]), .rdlo_in(a6_wr[1457]),  .coef_in(coef[64]), .rdup_out(a7_wr[1441]), .rdlo_out(a7_wr[1457]));
			radix2 #(.width(width)) rd_st6_1442  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1442]), .rdlo_in(a6_wr[1458]),  .coef_in(coef[128]), .rdup_out(a7_wr[1442]), .rdlo_out(a7_wr[1458]));
			radix2 #(.width(width)) rd_st6_1443  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1443]), .rdlo_in(a6_wr[1459]),  .coef_in(coef[192]), .rdup_out(a7_wr[1443]), .rdlo_out(a7_wr[1459]));
			radix2 #(.width(width)) rd_st6_1444  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1444]), .rdlo_in(a6_wr[1460]),  .coef_in(coef[256]), .rdup_out(a7_wr[1444]), .rdlo_out(a7_wr[1460]));
			radix2 #(.width(width)) rd_st6_1445  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1445]), .rdlo_in(a6_wr[1461]),  .coef_in(coef[320]), .rdup_out(a7_wr[1445]), .rdlo_out(a7_wr[1461]));
			radix2 #(.width(width)) rd_st6_1446  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1446]), .rdlo_in(a6_wr[1462]),  .coef_in(coef[384]), .rdup_out(a7_wr[1446]), .rdlo_out(a7_wr[1462]));
			radix2 #(.width(width)) rd_st6_1447  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1447]), .rdlo_in(a6_wr[1463]),  .coef_in(coef[448]), .rdup_out(a7_wr[1447]), .rdlo_out(a7_wr[1463]));
			radix2 #(.width(width)) rd_st6_1448  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1448]), .rdlo_in(a6_wr[1464]),  .coef_in(coef[512]), .rdup_out(a7_wr[1448]), .rdlo_out(a7_wr[1464]));
			radix2 #(.width(width)) rd_st6_1449  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1449]), .rdlo_in(a6_wr[1465]),  .coef_in(coef[576]), .rdup_out(a7_wr[1449]), .rdlo_out(a7_wr[1465]));
			radix2 #(.width(width)) rd_st6_1450  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1450]), .rdlo_in(a6_wr[1466]),  .coef_in(coef[640]), .rdup_out(a7_wr[1450]), .rdlo_out(a7_wr[1466]));
			radix2 #(.width(width)) rd_st6_1451  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1451]), .rdlo_in(a6_wr[1467]),  .coef_in(coef[704]), .rdup_out(a7_wr[1451]), .rdlo_out(a7_wr[1467]));
			radix2 #(.width(width)) rd_st6_1452  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1452]), .rdlo_in(a6_wr[1468]),  .coef_in(coef[768]), .rdup_out(a7_wr[1452]), .rdlo_out(a7_wr[1468]));
			radix2 #(.width(width)) rd_st6_1453  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1453]), .rdlo_in(a6_wr[1469]),  .coef_in(coef[832]), .rdup_out(a7_wr[1453]), .rdlo_out(a7_wr[1469]));
			radix2 #(.width(width)) rd_st6_1454  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1454]), .rdlo_in(a6_wr[1470]),  .coef_in(coef[896]), .rdup_out(a7_wr[1454]), .rdlo_out(a7_wr[1470]));
			radix2 #(.width(width)) rd_st6_1455  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1455]), .rdlo_in(a6_wr[1471]),  .coef_in(coef[960]), .rdup_out(a7_wr[1455]), .rdlo_out(a7_wr[1471]));
			radix2 #(.width(width)) rd_st6_1472  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1472]), .rdlo_in(a6_wr[1488]),  .coef_in(coef[0]), .rdup_out(a7_wr[1472]), .rdlo_out(a7_wr[1488]));
			radix2 #(.width(width)) rd_st6_1473  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1473]), .rdlo_in(a6_wr[1489]),  .coef_in(coef[64]), .rdup_out(a7_wr[1473]), .rdlo_out(a7_wr[1489]));
			radix2 #(.width(width)) rd_st6_1474  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1474]), .rdlo_in(a6_wr[1490]),  .coef_in(coef[128]), .rdup_out(a7_wr[1474]), .rdlo_out(a7_wr[1490]));
			radix2 #(.width(width)) rd_st6_1475  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1475]), .rdlo_in(a6_wr[1491]),  .coef_in(coef[192]), .rdup_out(a7_wr[1475]), .rdlo_out(a7_wr[1491]));
			radix2 #(.width(width)) rd_st6_1476  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1476]), .rdlo_in(a6_wr[1492]),  .coef_in(coef[256]), .rdup_out(a7_wr[1476]), .rdlo_out(a7_wr[1492]));
			radix2 #(.width(width)) rd_st6_1477  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1477]), .rdlo_in(a6_wr[1493]),  .coef_in(coef[320]), .rdup_out(a7_wr[1477]), .rdlo_out(a7_wr[1493]));
			radix2 #(.width(width)) rd_st6_1478  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1478]), .rdlo_in(a6_wr[1494]),  .coef_in(coef[384]), .rdup_out(a7_wr[1478]), .rdlo_out(a7_wr[1494]));
			radix2 #(.width(width)) rd_st6_1479  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1479]), .rdlo_in(a6_wr[1495]),  .coef_in(coef[448]), .rdup_out(a7_wr[1479]), .rdlo_out(a7_wr[1495]));
			radix2 #(.width(width)) rd_st6_1480  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1480]), .rdlo_in(a6_wr[1496]),  .coef_in(coef[512]), .rdup_out(a7_wr[1480]), .rdlo_out(a7_wr[1496]));
			radix2 #(.width(width)) rd_st6_1481  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1481]), .rdlo_in(a6_wr[1497]),  .coef_in(coef[576]), .rdup_out(a7_wr[1481]), .rdlo_out(a7_wr[1497]));
			radix2 #(.width(width)) rd_st6_1482  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1482]), .rdlo_in(a6_wr[1498]),  .coef_in(coef[640]), .rdup_out(a7_wr[1482]), .rdlo_out(a7_wr[1498]));
			radix2 #(.width(width)) rd_st6_1483  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1483]), .rdlo_in(a6_wr[1499]),  .coef_in(coef[704]), .rdup_out(a7_wr[1483]), .rdlo_out(a7_wr[1499]));
			radix2 #(.width(width)) rd_st6_1484  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1484]), .rdlo_in(a6_wr[1500]),  .coef_in(coef[768]), .rdup_out(a7_wr[1484]), .rdlo_out(a7_wr[1500]));
			radix2 #(.width(width)) rd_st6_1485  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1485]), .rdlo_in(a6_wr[1501]),  .coef_in(coef[832]), .rdup_out(a7_wr[1485]), .rdlo_out(a7_wr[1501]));
			radix2 #(.width(width)) rd_st6_1486  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1486]), .rdlo_in(a6_wr[1502]),  .coef_in(coef[896]), .rdup_out(a7_wr[1486]), .rdlo_out(a7_wr[1502]));
			radix2 #(.width(width)) rd_st6_1487  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1487]), .rdlo_in(a6_wr[1503]),  .coef_in(coef[960]), .rdup_out(a7_wr[1487]), .rdlo_out(a7_wr[1503]));
			radix2 #(.width(width)) rd_st6_1504  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1504]), .rdlo_in(a6_wr[1520]),  .coef_in(coef[0]), .rdup_out(a7_wr[1504]), .rdlo_out(a7_wr[1520]));
			radix2 #(.width(width)) rd_st6_1505  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1505]), .rdlo_in(a6_wr[1521]),  .coef_in(coef[64]), .rdup_out(a7_wr[1505]), .rdlo_out(a7_wr[1521]));
			radix2 #(.width(width)) rd_st6_1506  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1506]), .rdlo_in(a6_wr[1522]),  .coef_in(coef[128]), .rdup_out(a7_wr[1506]), .rdlo_out(a7_wr[1522]));
			radix2 #(.width(width)) rd_st6_1507  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1507]), .rdlo_in(a6_wr[1523]),  .coef_in(coef[192]), .rdup_out(a7_wr[1507]), .rdlo_out(a7_wr[1523]));
			radix2 #(.width(width)) rd_st6_1508  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1508]), .rdlo_in(a6_wr[1524]),  .coef_in(coef[256]), .rdup_out(a7_wr[1508]), .rdlo_out(a7_wr[1524]));
			radix2 #(.width(width)) rd_st6_1509  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1509]), .rdlo_in(a6_wr[1525]),  .coef_in(coef[320]), .rdup_out(a7_wr[1509]), .rdlo_out(a7_wr[1525]));
			radix2 #(.width(width)) rd_st6_1510  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1510]), .rdlo_in(a6_wr[1526]),  .coef_in(coef[384]), .rdup_out(a7_wr[1510]), .rdlo_out(a7_wr[1526]));
			radix2 #(.width(width)) rd_st6_1511  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1511]), .rdlo_in(a6_wr[1527]),  .coef_in(coef[448]), .rdup_out(a7_wr[1511]), .rdlo_out(a7_wr[1527]));
			radix2 #(.width(width)) rd_st6_1512  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1512]), .rdlo_in(a6_wr[1528]),  .coef_in(coef[512]), .rdup_out(a7_wr[1512]), .rdlo_out(a7_wr[1528]));
			radix2 #(.width(width)) rd_st6_1513  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1513]), .rdlo_in(a6_wr[1529]),  .coef_in(coef[576]), .rdup_out(a7_wr[1513]), .rdlo_out(a7_wr[1529]));
			radix2 #(.width(width)) rd_st6_1514  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1514]), .rdlo_in(a6_wr[1530]),  .coef_in(coef[640]), .rdup_out(a7_wr[1514]), .rdlo_out(a7_wr[1530]));
			radix2 #(.width(width)) rd_st6_1515  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1515]), .rdlo_in(a6_wr[1531]),  .coef_in(coef[704]), .rdup_out(a7_wr[1515]), .rdlo_out(a7_wr[1531]));
			radix2 #(.width(width)) rd_st6_1516  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1516]), .rdlo_in(a6_wr[1532]),  .coef_in(coef[768]), .rdup_out(a7_wr[1516]), .rdlo_out(a7_wr[1532]));
			radix2 #(.width(width)) rd_st6_1517  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1517]), .rdlo_in(a6_wr[1533]),  .coef_in(coef[832]), .rdup_out(a7_wr[1517]), .rdlo_out(a7_wr[1533]));
			radix2 #(.width(width)) rd_st6_1518  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1518]), .rdlo_in(a6_wr[1534]),  .coef_in(coef[896]), .rdup_out(a7_wr[1518]), .rdlo_out(a7_wr[1534]));
			radix2 #(.width(width)) rd_st6_1519  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1519]), .rdlo_in(a6_wr[1535]),  .coef_in(coef[960]), .rdup_out(a7_wr[1519]), .rdlo_out(a7_wr[1535]));
			radix2 #(.width(width)) rd_st6_1536  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1536]), .rdlo_in(a6_wr[1552]),  .coef_in(coef[0]), .rdup_out(a7_wr[1536]), .rdlo_out(a7_wr[1552]));
			radix2 #(.width(width)) rd_st6_1537  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1537]), .rdlo_in(a6_wr[1553]),  .coef_in(coef[64]), .rdup_out(a7_wr[1537]), .rdlo_out(a7_wr[1553]));
			radix2 #(.width(width)) rd_st6_1538  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1538]), .rdlo_in(a6_wr[1554]),  .coef_in(coef[128]), .rdup_out(a7_wr[1538]), .rdlo_out(a7_wr[1554]));
			radix2 #(.width(width)) rd_st6_1539  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1539]), .rdlo_in(a6_wr[1555]),  .coef_in(coef[192]), .rdup_out(a7_wr[1539]), .rdlo_out(a7_wr[1555]));
			radix2 #(.width(width)) rd_st6_1540  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1540]), .rdlo_in(a6_wr[1556]),  .coef_in(coef[256]), .rdup_out(a7_wr[1540]), .rdlo_out(a7_wr[1556]));
			radix2 #(.width(width)) rd_st6_1541  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1541]), .rdlo_in(a6_wr[1557]),  .coef_in(coef[320]), .rdup_out(a7_wr[1541]), .rdlo_out(a7_wr[1557]));
			radix2 #(.width(width)) rd_st6_1542  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1542]), .rdlo_in(a6_wr[1558]),  .coef_in(coef[384]), .rdup_out(a7_wr[1542]), .rdlo_out(a7_wr[1558]));
			radix2 #(.width(width)) rd_st6_1543  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1543]), .rdlo_in(a6_wr[1559]),  .coef_in(coef[448]), .rdup_out(a7_wr[1543]), .rdlo_out(a7_wr[1559]));
			radix2 #(.width(width)) rd_st6_1544  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1544]), .rdlo_in(a6_wr[1560]),  .coef_in(coef[512]), .rdup_out(a7_wr[1544]), .rdlo_out(a7_wr[1560]));
			radix2 #(.width(width)) rd_st6_1545  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1545]), .rdlo_in(a6_wr[1561]),  .coef_in(coef[576]), .rdup_out(a7_wr[1545]), .rdlo_out(a7_wr[1561]));
			radix2 #(.width(width)) rd_st6_1546  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1546]), .rdlo_in(a6_wr[1562]),  .coef_in(coef[640]), .rdup_out(a7_wr[1546]), .rdlo_out(a7_wr[1562]));
			radix2 #(.width(width)) rd_st6_1547  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1547]), .rdlo_in(a6_wr[1563]),  .coef_in(coef[704]), .rdup_out(a7_wr[1547]), .rdlo_out(a7_wr[1563]));
			radix2 #(.width(width)) rd_st6_1548  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1548]), .rdlo_in(a6_wr[1564]),  .coef_in(coef[768]), .rdup_out(a7_wr[1548]), .rdlo_out(a7_wr[1564]));
			radix2 #(.width(width)) rd_st6_1549  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1549]), .rdlo_in(a6_wr[1565]),  .coef_in(coef[832]), .rdup_out(a7_wr[1549]), .rdlo_out(a7_wr[1565]));
			radix2 #(.width(width)) rd_st6_1550  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1550]), .rdlo_in(a6_wr[1566]),  .coef_in(coef[896]), .rdup_out(a7_wr[1550]), .rdlo_out(a7_wr[1566]));
			radix2 #(.width(width)) rd_st6_1551  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1551]), .rdlo_in(a6_wr[1567]),  .coef_in(coef[960]), .rdup_out(a7_wr[1551]), .rdlo_out(a7_wr[1567]));
			radix2 #(.width(width)) rd_st6_1568  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1568]), .rdlo_in(a6_wr[1584]),  .coef_in(coef[0]), .rdup_out(a7_wr[1568]), .rdlo_out(a7_wr[1584]));
			radix2 #(.width(width)) rd_st6_1569  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1569]), .rdlo_in(a6_wr[1585]),  .coef_in(coef[64]), .rdup_out(a7_wr[1569]), .rdlo_out(a7_wr[1585]));
			radix2 #(.width(width)) rd_st6_1570  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1570]), .rdlo_in(a6_wr[1586]),  .coef_in(coef[128]), .rdup_out(a7_wr[1570]), .rdlo_out(a7_wr[1586]));
			radix2 #(.width(width)) rd_st6_1571  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1571]), .rdlo_in(a6_wr[1587]),  .coef_in(coef[192]), .rdup_out(a7_wr[1571]), .rdlo_out(a7_wr[1587]));
			radix2 #(.width(width)) rd_st6_1572  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1572]), .rdlo_in(a6_wr[1588]),  .coef_in(coef[256]), .rdup_out(a7_wr[1572]), .rdlo_out(a7_wr[1588]));
			radix2 #(.width(width)) rd_st6_1573  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1573]), .rdlo_in(a6_wr[1589]),  .coef_in(coef[320]), .rdup_out(a7_wr[1573]), .rdlo_out(a7_wr[1589]));
			radix2 #(.width(width)) rd_st6_1574  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1574]), .rdlo_in(a6_wr[1590]),  .coef_in(coef[384]), .rdup_out(a7_wr[1574]), .rdlo_out(a7_wr[1590]));
			radix2 #(.width(width)) rd_st6_1575  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1575]), .rdlo_in(a6_wr[1591]),  .coef_in(coef[448]), .rdup_out(a7_wr[1575]), .rdlo_out(a7_wr[1591]));
			radix2 #(.width(width)) rd_st6_1576  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1576]), .rdlo_in(a6_wr[1592]),  .coef_in(coef[512]), .rdup_out(a7_wr[1576]), .rdlo_out(a7_wr[1592]));
			radix2 #(.width(width)) rd_st6_1577  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1577]), .rdlo_in(a6_wr[1593]),  .coef_in(coef[576]), .rdup_out(a7_wr[1577]), .rdlo_out(a7_wr[1593]));
			radix2 #(.width(width)) rd_st6_1578  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1578]), .rdlo_in(a6_wr[1594]),  .coef_in(coef[640]), .rdup_out(a7_wr[1578]), .rdlo_out(a7_wr[1594]));
			radix2 #(.width(width)) rd_st6_1579  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1579]), .rdlo_in(a6_wr[1595]),  .coef_in(coef[704]), .rdup_out(a7_wr[1579]), .rdlo_out(a7_wr[1595]));
			radix2 #(.width(width)) rd_st6_1580  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1580]), .rdlo_in(a6_wr[1596]),  .coef_in(coef[768]), .rdup_out(a7_wr[1580]), .rdlo_out(a7_wr[1596]));
			radix2 #(.width(width)) rd_st6_1581  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1581]), .rdlo_in(a6_wr[1597]),  .coef_in(coef[832]), .rdup_out(a7_wr[1581]), .rdlo_out(a7_wr[1597]));
			radix2 #(.width(width)) rd_st6_1582  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1582]), .rdlo_in(a6_wr[1598]),  .coef_in(coef[896]), .rdup_out(a7_wr[1582]), .rdlo_out(a7_wr[1598]));
			radix2 #(.width(width)) rd_st6_1583  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1583]), .rdlo_in(a6_wr[1599]),  .coef_in(coef[960]), .rdup_out(a7_wr[1583]), .rdlo_out(a7_wr[1599]));
			radix2 #(.width(width)) rd_st6_1600  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1600]), .rdlo_in(a6_wr[1616]),  .coef_in(coef[0]), .rdup_out(a7_wr[1600]), .rdlo_out(a7_wr[1616]));
			radix2 #(.width(width)) rd_st6_1601  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1601]), .rdlo_in(a6_wr[1617]),  .coef_in(coef[64]), .rdup_out(a7_wr[1601]), .rdlo_out(a7_wr[1617]));
			radix2 #(.width(width)) rd_st6_1602  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1602]), .rdlo_in(a6_wr[1618]),  .coef_in(coef[128]), .rdup_out(a7_wr[1602]), .rdlo_out(a7_wr[1618]));
			radix2 #(.width(width)) rd_st6_1603  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1603]), .rdlo_in(a6_wr[1619]),  .coef_in(coef[192]), .rdup_out(a7_wr[1603]), .rdlo_out(a7_wr[1619]));
			radix2 #(.width(width)) rd_st6_1604  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1604]), .rdlo_in(a6_wr[1620]),  .coef_in(coef[256]), .rdup_out(a7_wr[1604]), .rdlo_out(a7_wr[1620]));
			radix2 #(.width(width)) rd_st6_1605  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1605]), .rdlo_in(a6_wr[1621]),  .coef_in(coef[320]), .rdup_out(a7_wr[1605]), .rdlo_out(a7_wr[1621]));
			radix2 #(.width(width)) rd_st6_1606  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1606]), .rdlo_in(a6_wr[1622]),  .coef_in(coef[384]), .rdup_out(a7_wr[1606]), .rdlo_out(a7_wr[1622]));
			radix2 #(.width(width)) rd_st6_1607  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1607]), .rdlo_in(a6_wr[1623]),  .coef_in(coef[448]), .rdup_out(a7_wr[1607]), .rdlo_out(a7_wr[1623]));
			radix2 #(.width(width)) rd_st6_1608  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1608]), .rdlo_in(a6_wr[1624]),  .coef_in(coef[512]), .rdup_out(a7_wr[1608]), .rdlo_out(a7_wr[1624]));
			radix2 #(.width(width)) rd_st6_1609  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1609]), .rdlo_in(a6_wr[1625]),  .coef_in(coef[576]), .rdup_out(a7_wr[1609]), .rdlo_out(a7_wr[1625]));
			radix2 #(.width(width)) rd_st6_1610  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1610]), .rdlo_in(a6_wr[1626]),  .coef_in(coef[640]), .rdup_out(a7_wr[1610]), .rdlo_out(a7_wr[1626]));
			radix2 #(.width(width)) rd_st6_1611  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1611]), .rdlo_in(a6_wr[1627]),  .coef_in(coef[704]), .rdup_out(a7_wr[1611]), .rdlo_out(a7_wr[1627]));
			radix2 #(.width(width)) rd_st6_1612  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1612]), .rdlo_in(a6_wr[1628]),  .coef_in(coef[768]), .rdup_out(a7_wr[1612]), .rdlo_out(a7_wr[1628]));
			radix2 #(.width(width)) rd_st6_1613  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1613]), .rdlo_in(a6_wr[1629]),  .coef_in(coef[832]), .rdup_out(a7_wr[1613]), .rdlo_out(a7_wr[1629]));
			radix2 #(.width(width)) rd_st6_1614  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1614]), .rdlo_in(a6_wr[1630]),  .coef_in(coef[896]), .rdup_out(a7_wr[1614]), .rdlo_out(a7_wr[1630]));
			radix2 #(.width(width)) rd_st6_1615  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1615]), .rdlo_in(a6_wr[1631]),  .coef_in(coef[960]), .rdup_out(a7_wr[1615]), .rdlo_out(a7_wr[1631]));
			radix2 #(.width(width)) rd_st6_1632  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1632]), .rdlo_in(a6_wr[1648]),  .coef_in(coef[0]), .rdup_out(a7_wr[1632]), .rdlo_out(a7_wr[1648]));
			radix2 #(.width(width)) rd_st6_1633  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1633]), .rdlo_in(a6_wr[1649]),  .coef_in(coef[64]), .rdup_out(a7_wr[1633]), .rdlo_out(a7_wr[1649]));
			radix2 #(.width(width)) rd_st6_1634  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1634]), .rdlo_in(a6_wr[1650]),  .coef_in(coef[128]), .rdup_out(a7_wr[1634]), .rdlo_out(a7_wr[1650]));
			radix2 #(.width(width)) rd_st6_1635  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1635]), .rdlo_in(a6_wr[1651]),  .coef_in(coef[192]), .rdup_out(a7_wr[1635]), .rdlo_out(a7_wr[1651]));
			radix2 #(.width(width)) rd_st6_1636  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1636]), .rdlo_in(a6_wr[1652]),  .coef_in(coef[256]), .rdup_out(a7_wr[1636]), .rdlo_out(a7_wr[1652]));
			radix2 #(.width(width)) rd_st6_1637  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1637]), .rdlo_in(a6_wr[1653]),  .coef_in(coef[320]), .rdup_out(a7_wr[1637]), .rdlo_out(a7_wr[1653]));
			radix2 #(.width(width)) rd_st6_1638  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1638]), .rdlo_in(a6_wr[1654]),  .coef_in(coef[384]), .rdup_out(a7_wr[1638]), .rdlo_out(a7_wr[1654]));
			radix2 #(.width(width)) rd_st6_1639  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1639]), .rdlo_in(a6_wr[1655]),  .coef_in(coef[448]), .rdup_out(a7_wr[1639]), .rdlo_out(a7_wr[1655]));
			radix2 #(.width(width)) rd_st6_1640  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1640]), .rdlo_in(a6_wr[1656]),  .coef_in(coef[512]), .rdup_out(a7_wr[1640]), .rdlo_out(a7_wr[1656]));
			radix2 #(.width(width)) rd_st6_1641  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1641]), .rdlo_in(a6_wr[1657]),  .coef_in(coef[576]), .rdup_out(a7_wr[1641]), .rdlo_out(a7_wr[1657]));
			radix2 #(.width(width)) rd_st6_1642  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1642]), .rdlo_in(a6_wr[1658]),  .coef_in(coef[640]), .rdup_out(a7_wr[1642]), .rdlo_out(a7_wr[1658]));
			radix2 #(.width(width)) rd_st6_1643  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1643]), .rdlo_in(a6_wr[1659]),  .coef_in(coef[704]), .rdup_out(a7_wr[1643]), .rdlo_out(a7_wr[1659]));
			radix2 #(.width(width)) rd_st6_1644  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1644]), .rdlo_in(a6_wr[1660]),  .coef_in(coef[768]), .rdup_out(a7_wr[1644]), .rdlo_out(a7_wr[1660]));
			radix2 #(.width(width)) rd_st6_1645  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1645]), .rdlo_in(a6_wr[1661]),  .coef_in(coef[832]), .rdup_out(a7_wr[1645]), .rdlo_out(a7_wr[1661]));
			radix2 #(.width(width)) rd_st6_1646  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1646]), .rdlo_in(a6_wr[1662]),  .coef_in(coef[896]), .rdup_out(a7_wr[1646]), .rdlo_out(a7_wr[1662]));
			radix2 #(.width(width)) rd_st6_1647  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1647]), .rdlo_in(a6_wr[1663]),  .coef_in(coef[960]), .rdup_out(a7_wr[1647]), .rdlo_out(a7_wr[1663]));
			radix2 #(.width(width)) rd_st6_1664  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1664]), .rdlo_in(a6_wr[1680]),  .coef_in(coef[0]), .rdup_out(a7_wr[1664]), .rdlo_out(a7_wr[1680]));
			radix2 #(.width(width)) rd_st6_1665  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1665]), .rdlo_in(a6_wr[1681]),  .coef_in(coef[64]), .rdup_out(a7_wr[1665]), .rdlo_out(a7_wr[1681]));
			radix2 #(.width(width)) rd_st6_1666  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1666]), .rdlo_in(a6_wr[1682]),  .coef_in(coef[128]), .rdup_out(a7_wr[1666]), .rdlo_out(a7_wr[1682]));
			radix2 #(.width(width)) rd_st6_1667  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1667]), .rdlo_in(a6_wr[1683]),  .coef_in(coef[192]), .rdup_out(a7_wr[1667]), .rdlo_out(a7_wr[1683]));
			radix2 #(.width(width)) rd_st6_1668  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1668]), .rdlo_in(a6_wr[1684]),  .coef_in(coef[256]), .rdup_out(a7_wr[1668]), .rdlo_out(a7_wr[1684]));
			radix2 #(.width(width)) rd_st6_1669  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1669]), .rdlo_in(a6_wr[1685]),  .coef_in(coef[320]), .rdup_out(a7_wr[1669]), .rdlo_out(a7_wr[1685]));
			radix2 #(.width(width)) rd_st6_1670  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1670]), .rdlo_in(a6_wr[1686]),  .coef_in(coef[384]), .rdup_out(a7_wr[1670]), .rdlo_out(a7_wr[1686]));
			radix2 #(.width(width)) rd_st6_1671  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1671]), .rdlo_in(a6_wr[1687]),  .coef_in(coef[448]), .rdup_out(a7_wr[1671]), .rdlo_out(a7_wr[1687]));
			radix2 #(.width(width)) rd_st6_1672  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1672]), .rdlo_in(a6_wr[1688]),  .coef_in(coef[512]), .rdup_out(a7_wr[1672]), .rdlo_out(a7_wr[1688]));
			radix2 #(.width(width)) rd_st6_1673  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1673]), .rdlo_in(a6_wr[1689]),  .coef_in(coef[576]), .rdup_out(a7_wr[1673]), .rdlo_out(a7_wr[1689]));
			radix2 #(.width(width)) rd_st6_1674  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1674]), .rdlo_in(a6_wr[1690]),  .coef_in(coef[640]), .rdup_out(a7_wr[1674]), .rdlo_out(a7_wr[1690]));
			radix2 #(.width(width)) rd_st6_1675  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1675]), .rdlo_in(a6_wr[1691]),  .coef_in(coef[704]), .rdup_out(a7_wr[1675]), .rdlo_out(a7_wr[1691]));
			radix2 #(.width(width)) rd_st6_1676  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1676]), .rdlo_in(a6_wr[1692]),  .coef_in(coef[768]), .rdup_out(a7_wr[1676]), .rdlo_out(a7_wr[1692]));
			radix2 #(.width(width)) rd_st6_1677  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1677]), .rdlo_in(a6_wr[1693]),  .coef_in(coef[832]), .rdup_out(a7_wr[1677]), .rdlo_out(a7_wr[1693]));
			radix2 #(.width(width)) rd_st6_1678  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1678]), .rdlo_in(a6_wr[1694]),  .coef_in(coef[896]), .rdup_out(a7_wr[1678]), .rdlo_out(a7_wr[1694]));
			radix2 #(.width(width)) rd_st6_1679  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1679]), .rdlo_in(a6_wr[1695]),  .coef_in(coef[960]), .rdup_out(a7_wr[1679]), .rdlo_out(a7_wr[1695]));
			radix2 #(.width(width)) rd_st6_1696  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1696]), .rdlo_in(a6_wr[1712]),  .coef_in(coef[0]), .rdup_out(a7_wr[1696]), .rdlo_out(a7_wr[1712]));
			radix2 #(.width(width)) rd_st6_1697  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1697]), .rdlo_in(a6_wr[1713]),  .coef_in(coef[64]), .rdup_out(a7_wr[1697]), .rdlo_out(a7_wr[1713]));
			radix2 #(.width(width)) rd_st6_1698  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1698]), .rdlo_in(a6_wr[1714]),  .coef_in(coef[128]), .rdup_out(a7_wr[1698]), .rdlo_out(a7_wr[1714]));
			radix2 #(.width(width)) rd_st6_1699  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1699]), .rdlo_in(a6_wr[1715]),  .coef_in(coef[192]), .rdup_out(a7_wr[1699]), .rdlo_out(a7_wr[1715]));
			radix2 #(.width(width)) rd_st6_1700  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1700]), .rdlo_in(a6_wr[1716]),  .coef_in(coef[256]), .rdup_out(a7_wr[1700]), .rdlo_out(a7_wr[1716]));
			radix2 #(.width(width)) rd_st6_1701  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1701]), .rdlo_in(a6_wr[1717]),  .coef_in(coef[320]), .rdup_out(a7_wr[1701]), .rdlo_out(a7_wr[1717]));
			radix2 #(.width(width)) rd_st6_1702  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1702]), .rdlo_in(a6_wr[1718]),  .coef_in(coef[384]), .rdup_out(a7_wr[1702]), .rdlo_out(a7_wr[1718]));
			radix2 #(.width(width)) rd_st6_1703  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1703]), .rdlo_in(a6_wr[1719]),  .coef_in(coef[448]), .rdup_out(a7_wr[1703]), .rdlo_out(a7_wr[1719]));
			radix2 #(.width(width)) rd_st6_1704  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1704]), .rdlo_in(a6_wr[1720]),  .coef_in(coef[512]), .rdup_out(a7_wr[1704]), .rdlo_out(a7_wr[1720]));
			radix2 #(.width(width)) rd_st6_1705  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1705]), .rdlo_in(a6_wr[1721]),  .coef_in(coef[576]), .rdup_out(a7_wr[1705]), .rdlo_out(a7_wr[1721]));
			radix2 #(.width(width)) rd_st6_1706  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1706]), .rdlo_in(a6_wr[1722]),  .coef_in(coef[640]), .rdup_out(a7_wr[1706]), .rdlo_out(a7_wr[1722]));
			radix2 #(.width(width)) rd_st6_1707  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1707]), .rdlo_in(a6_wr[1723]),  .coef_in(coef[704]), .rdup_out(a7_wr[1707]), .rdlo_out(a7_wr[1723]));
			radix2 #(.width(width)) rd_st6_1708  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1708]), .rdlo_in(a6_wr[1724]),  .coef_in(coef[768]), .rdup_out(a7_wr[1708]), .rdlo_out(a7_wr[1724]));
			radix2 #(.width(width)) rd_st6_1709  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1709]), .rdlo_in(a6_wr[1725]),  .coef_in(coef[832]), .rdup_out(a7_wr[1709]), .rdlo_out(a7_wr[1725]));
			radix2 #(.width(width)) rd_st6_1710  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1710]), .rdlo_in(a6_wr[1726]),  .coef_in(coef[896]), .rdup_out(a7_wr[1710]), .rdlo_out(a7_wr[1726]));
			radix2 #(.width(width)) rd_st6_1711  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1711]), .rdlo_in(a6_wr[1727]),  .coef_in(coef[960]), .rdup_out(a7_wr[1711]), .rdlo_out(a7_wr[1727]));
			radix2 #(.width(width)) rd_st6_1728  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1728]), .rdlo_in(a6_wr[1744]),  .coef_in(coef[0]), .rdup_out(a7_wr[1728]), .rdlo_out(a7_wr[1744]));
			radix2 #(.width(width)) rd_st6_1729  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1729]), .rdlo_in(a6_wr[1745]),  .coef_in(coef[64]), .rdup_out(a7_wr[1729]), .rdlo_out(a7_wr[1745]));
			radix2 #(.width(width)) rd_st6_1730  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1730]), .rdlo_in(a6_wr[1746]),  .coef_in(coef[128]), .rdup_out(a7_wr[1730]), .rdlo_out(a7_wr[1746]));
			radix2 #(.width(width)) rd_st6_1731  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1731]), .rdlo_in(a6_wr[1747]),  .coef_in(coef[192]), .rdup_out(a7_wr[1731]), .rdlo_out(a7_wr[1747]));
			radix2 #(.width(width)) rd_st6_1732  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1732]), .rdlo_in(a6_wr[1748]),  .coef_in(coef[256]), .rdup_out(a7_wr[1732]), .rdlo_out(a7_wr[1748]));
			radix2 #(.width(width)) rd_st6_1733  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1733]), .rdlo_in(a6_wr[1749]),  .coef_in(coef[320]), .rdup_out(a7_wr[1733]), .rdlo_out(a7_wr[1749]));
			radix2 #(.width(width)) rd_st6_1734  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1734]), .rdlo_in(a6_wr[1750]),  .coef_in(coef[384]), .rdup_out(a7_wr[1734]), .rdlo_out(a7_wr[1750]));
			radix2 #(.width(width)) rd_st6_1735  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1735]), .rdlo_in(a6_wr[1751]),  .coef_in(coef[448]), .rdup_out(a7_wr[1735]), .rdlo_out(a7_wr[1751]));
			radix2 #(.width(width)) rd_st6_1736  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1736]), .rdlo_in(a6_wr[1752]),  .coef_in(coef[512]), .rdup_out(a7_wr[1736]), .rdlo_out(a7_wr[1752]));
			radix2 #(.width(width)) rd_st6_1737  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1737]), .rdlo_in(a6_wr[1753]),  .coef_in(coef[576]), .rdup_out(a7_wr[1737]), .rdlo_out(a7_wr[1753]));
			radix2 #(.width(width)) rd_st6_1738  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1738]), .rdlo_in(a6_wr[1754]),  .coef_in(coef[640]), .rdup_out(a7_wr[1738]), .rdlo_out(a7_wr[1754]));
			radix2 #(.width(width)) rd_st6_1739  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1739]), .rdlo_in(a6_wr[1755]),  .coef_in(coef[704]), .rdup_out(a7_wr[1739]), .rdlo_out(a7_wr[1755]));
			radix2 #(.width(width)) rd_st6_1740  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1740]), .rdlo_in(a6_wr[1756]),  .coef_in(coef[768]), .rdup_out(a7_wr[1740]), .rdlo_out(a7_wr[1756]));
			radix2 #(.width(width)) rd_st6_1741  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1741]), .rdlo_in(a6_wr[1757]),  .coef_in(coef[832]), .rdup_out(a7_wr[1741]), .rdlo_out(a7_wr[1757]));
			radix2 #(.width(width)) rd_st6_1742  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1742]), .rdlo_in(a6_wr[1758]),  .coef_in(coef[896]), .rdup_out(a7_wr[1742]), .rdlo_out(a7_wr[1758]));
			radix2 #(.width(width)) rd_st6_1743  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1743]), .rdlo_in(a6_wr[1759]),  .coef_in(coef[960]), .rdup_out(a7_wr[1743]), .rdlo_out(a7_wr[1759]));
			radix2 #(.width(width)) rd_st6_1760  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1760]), .rdlo_in(a6_wr[1776]),  .coef_in(coef[0]), .rdup_out(a7_wr[1760]), .rdlo_out(a7_wr[1776]));
			radix2 #(.width(width)) rd_st6_1761  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1761]), .rdlo_in(a6_wr[1777]),  .coef_in(coef[64]), .rdup_out(a7_wr[1761]), .rdlo_out(a7_wr[1777]));
			radix2 #(.width(width)) rd_st6_1762  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1762]), .rdlo_in(a6_wr[1778]),  .coef_in(coef[128]), .rdup_out(a7_wr[1762]), .rdlo_out(a7_wr[1778]));
			radix2 #(.width(width)) rd_st6_1763  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1763]), .rdlo_in(a6_wr[1779]),  .coef_in(coef[192]), .rdup_out(a7_wr[1763]), .rdlo_out(a7_wr[1779]));
			radix2 #(.width(width)) rd_st6_1764  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1764]), .rdlo_in(a6_wr[1780]),  .coef_in(coef[256]), .rdup_out(a7_wr[1764]), .rdlo_out(a7_wr[1780]));
			radix2 #(.width(width)) rd_st6_1765  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1765]), .rdlo_in(a6_wr[1781]),  .coef_in(coef[320]), .rdup_out(a7_wr[1765]), .rdlo_out(a7_wr[1781]));
			radix2 #(.width(width)) rd_st6_1766  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1766]), .rdlo_in(a6_wr[1782]),  .coef_in(coef[384]), .rdup_out(a7_wr[1766]), .rdlo_out(a7_wr[1782]));
			radix2 #(.width(width)) rd_st6_1767  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1767]), .rdlo_in(a6_wr[1783]),  .coef_in(coef[448]), .rdup_out(a7_wr[1767]), .rdlo_out(a7_wr[1783]));
			radix2 #(.width(width)) rd_st6_1768  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1768]), .rdlo_in(a6_wr[1784]),  .coef_in(coef[512]), .rdup_out(a7_wr[1768]), .rdlo_out(a7_wr[1784]));
			radix2 #(.width(width)) rd_st6_1769  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1769]), .rdlo_in(a6_wr[1785]),  .coef_in(coef[576]), .rdup_out(a7_wr[1769]), .rdlo_out(a7_wr[1785]));
			radix2 #(.width(width)) rd_st6_1770  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1770]), .rdlo_in(a6_wr[1786]),  .coef_in(coef[640]), .rdup_out(a7_wr[1770]), .rdlo_out(a7_wr[1786]));
			radix2 #(.width(width)) rd_st6_1771  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1771]), .rdlo_in(a6_wr[1787]),  .coef_in(coef[704]), .rdup_out(a7_wr[1771]), .rdlo_out(a7_wr[1787]));
			radix2 #(.width(width)) rd_st6_1772  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1772]), .rdlo_in(a6_wr[1788]),  .coef_in(coef[768]), .rdup_out(a7_wr[1772]), .rdlo_out(a7_wr[1788]));
			radix2 #(.width(width)) rd_st6_1773  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1773]), .rdlo_in(a6_wr[1789]),  .coef_in(coef[832]), .rdup_out(a7_wr[1773]), .rdlo_out(a7_wr[1789]));
			radix2 #(.width(width)) rd_st6_1774  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1774]), .rdlo_in(a6_wr[1790]),  .coef_in(coef[896]), .rdup_out(a7_wr[1774]), .rdlo_out(a7_wr[1790]));
			radix2 #(.width(width)) rd_st6_1775  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1775]), .rdlo_in(a6_wr[1791]),  .coef_in(coef[960]), .rdup_out(a7_wr[1775]), .rdlo_out(a7_wr[1791]));
			radix2 #(.width(width)) rd_st6_1792  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1792]), .rdlo_in(a6_wr[1808]),  .coef_in(coef[0]), .rdup_out(a7_wr[1792]), .rdlo_out(a7_wr[1808]));
			radix2 #(.width(width)) rd_st6_1793  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1793]), .rdlo_in(a6_wr[1809]),  .coef_in(coef[64]), .rdup_out(a7_wr[1793]), .rdlo_out(a7_wr[1809]));
			radix2 #(.width(width)) rd_st6_1794  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1794]), .rdlo_in(a6_wr[1810]),  .coef_in(coef[128]), .rdup_out(a7_wr[1794]), .rdlo_out(a7_wr[1810]));
			radix2 #(.width(width)) rd_st6_1795  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1795]), .rdlo_in(a6_wr[1811]),  .coef_in(coef[192]), .rdup_out(a7_wr[1795]), .rdlo_out(a7_wr[1811]));
			radix2 #(.width(width)) rd_st6_1796  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1796]), .rdlo_in(a6_wr[1812]),  .coef_in(coef[256]), .rdup_out(a7_wr[1796]), .rdlo_out(a7_wr[1812]));
			radix2 #(.width(width)) rd_st6_1797  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1797]), .rdlo_in(a6_wr[1813]),  .coef_in(coef[320]), .rdup_out(a7_wr[1797]), .rdlo_out(a7_wr[1813]));
			radix2 #(.width(width)) rd_st6_1798  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1798]), .rdlo_in(a6_wr[1814]),  .coef_in(coef[384]), .rdup_out(a7_wr[1798]), .rdlo_out(a7_wr[1814]));
			radix2 #(.width(width)) rd_st6_1799  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1799]), .rdlo_in(a6_wr[1815]),  .coef_in(coef[448]), .rdup_out(a7_wr[1799]), .rdlo_out(a7_wr[1815]));
			radix2 #(.width(width)) rd_st6_1800  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1800]), .rdlo_in(a6_wr[1816]),  .coef_in(coef[512]), .rdup_out(a7_wr[1800]), .rdlo_out(a7_wr[1816]));
			radix2 #(.width(width)) rd_st6_1801  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1801]), .rdlo_in(a6_wr[1817]),  .coef_in(coef[576]), .rdup_out(a7_wr[1801]), .rdlo_out(a7_wr[1817]));
			radix2 #(.width(width)) rd_st6_1802  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1802]), .rdlo_in(a6_wr[1818]),  .coef_in(coef[640]), .rdup_out(a7_wr[1802]), .rdlo_out(a7_wr[1818]));
			radix2 #(.width(width)) rd_st6_1803  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1803]), .rdlo_in(a6_wr[1819]),  .coef_in(coef[704]), .rdup_out(a7_wr[1803]), .rdlo_out(a7_wr[1819]));
			radix2 #(.width(width)) rd_st6_1804  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1804]), .rdlo_in(a6_wr[1820]),  .coef_in(coef[768]), .rdup_out(a7_wr[1804]), .rdlo_out(a7_wr[1820]));
			radix2 #(.width(width)) rd_st6_1805  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1805]), .rdlo_in(a6_wr[1821]),  .coef_in(coef[832]), .rdup_out(a7_wr[1805]), .rdlo_out(a7_wr[1821]));
			radix2 #(.width(width)) rd_st6_1806  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1806]), .rdlo_in(a6_wr[1822]),  .coef_in(coef[896]), .rdup_out(a7_wr[1806]), .rdlo_out(a7_wr[1822]));
			radix2 #(.width(width)) rd_st6_1807  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1807]), .rdlo_in(a6_wr[1823]),  .coef_in(coef[960]), .rdup_out(a7_wr[1807]), .rdlo_out(a7_wr[1823]));
			radix2 #(.width(width)) rd_st6_1824  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1824]), .rdlo_in(a6_wr[1840]),  .coef_in(coef[0]), .rdup_out(a7_wr[1824]), .rdlo_out(a7_wr[1840]));
			radix2 #(.width(width)) rd_st6_1825  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1825]), .rdlo_in(a6_wr[1841]),  .coef_in(coef[64]), .rdup_out(a7_wr[1825]), .rdlo_out(a7_wr[1841]));
			radix2 #(.width(width)) rd_st6_1826  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1826]), .rdlo_in(a6_wr[1842]),  .coef_in(coef[128]), .rdup_out(a7_wr[1826]), .rdlo_out(a7_wr[1842]));
			radix2 #(.width(width)) rd_st6_1827  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1827]), .rdlo_in(a6_wr[1843]),  .coef_in(coef[192]), .rdup_out(a7_wr[1827]), .rdlo_out(a7_wr[1843]));
			radix2 #(.width(width)) rd_st6_1828  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1828]), .rdlo_in(a6_wr[1844]),  .coef_in(coef[256]), .rdup_out(a7_wr[1828]), .rdlo_out(a7_wr[1844]));
			radix2 #(.width(width)) rd_st6_1829  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1829]), .rdlo_in(a6_wr[1845]),  .coef_in(coef[320]), .rdup_out(a7_wr[1829]), .rdlo_out(a7_wr[1845]));
			radix2 #(.width(width)) rd_st6_1830  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1830]), .rdlo_in(a6_wr[1846]),  .coef_in(coef[384]), .rdup_out(a7_wr[1830]), .rdlo_out(a7_wr[1846]));
			radix2 #(.width(width)) rd_st6_1831  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1831]), .rdlo_in(a6_wr[1847]),  .coef_in(coef[448]), .rdup_out(a7_wr[1831]), .rdlo_out(a7_wr[1847]));
			radix2 #(.width(width)) rd_st6_1832  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1832]), .rdlo_in(a6_wr[1848]),  .coef_in(coef[512]), .rdup_out(a7_wr[1832]), .rdlo_out(a7_wr[1848]));
			radix2 #(.width(width)) rd_st6_1833  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1833]), .rdlo_in(a6_wr[1849]),  .coef_in(coef[576]), .rdup_out(a7_wr[1833]), .rdlo_out(a7_wr[1849]));
			radix2 #(.width(width)) rd_st6_1834  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1834]), .rdlo_in(a6_wr[1850]),  .coef_in(coef[640]), .rdup_out(a7_wr[1834]), .rdlo_out(a7_wr[1850]));
			radix2 #(.width(width)) rd_st6_1835  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1835]), .rdlo_in(a6_wr[1851]),  .coef_in(coef[704]), .rdup_out(a7_wr[1835]), .rdlo_out(a7_wr[1851]));
			radix2 #(.width(width)) rd_st6_1836  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1836]), .rdlo_in(a6_wr[1852]),  .coef_in(coef[768]), .rdup_out(a7_wr[1836]), .rdlo_out(a7_wr[1852]));
			radix2 #(.width(width)) rd_st6_1837  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1837]), .rdlo_in(a6_wr[1853]),  .coef_in(coef[832]), .rdup_out(a7_wr[1837]), .rdlo_out(a7_wr[1853]));
			radix2 #(.width(width)) rd_st6_1838  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1838]), .rdlo_in(a6_wr[1854]),  .coef_in(coef[896]), .rdup_out(a7_wr[1838]), .rdlo_out(a7_wr[1854]));
			radix2 #(.width(width)) rd_st6_1839  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1839]), .rdlo_in(a6_wr[1855]),  .coef_in(coef[960]), .rdup_out(a7_wr[1839]), .rdlo_out(a7_wr[1855]));
			radix2 #(.width(width)) rd_st6_1856  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1856]), .rdlo_in(a6_wr[1872]),  .coef_in(coef[0]), .rdup_out(a7_wr[1856]), .rdlo_out(a7_wr[1872]));
			radix2 #(.width(width)) rd_st6_1857  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1857]), .rdlo_in(a6_wr[1873]),  .coef_in(coef[64]), .rdup_out(a7_wr[1857]), .rdlo_out(a7_wr[1873]));
			radix2 #(.width(width)) rd_st6_1858  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1858]), .rdlo_in(a6_wr[1874]),  .coef_in(coef[128]), .rdup_out(a7_wr[1858]), .rdlo_out(a7_wr[1874]));
			radix2 #(.width(width)) rd_st6_1859  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1859]), .rdlo_in(a6_wr[1875]),  .coef_in(coef[192]), .rdup_out(a7_wr[1859]), .rdlo_out(a7_wr[1875]));
			radix2 #(.width(width)) rd_st6_1860  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1860]), .rdlo_in(a6_wr[1876]),  .coef_in(coef[256]), .rdup_out(a7_wr[1860]), .rdlo_out(a7_wr[1876]));
			radix2 #(.width(width)) rd_st6_1861  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1861]), .rdlo_in(a6_wr[1877]),  .coef_in(coef[320]), .rdup_out(a7_wr[1861]), .rdlo_out(a7_wr[1877]));
			radix2 #(.width(width)) rd_st6_1862  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1862]), .rdlo_in(a6_wr[1878]),  .coef_in(coef[384]), .rdup_out(a7_wr[1862]), .rdlo_out(a7_wr[1878]));
			radix2 #(.width(width)) rd_st6_1863  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1863]), .rdlo_in(a6_wr[1879]),  .coef_in(coef[448]), .rdup_out(a7_wr[1863]), .rdlo_out(a7_wr[1879]));
			radix2 #(.width(width)) rd_st6_1864  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1864]), .rdlo_in(a6_wr[1880]),  .coef_in(coef[512]), .rdup_out(a7_wr[1864]), .rdlo_out(a7_wr[1880]));
			radix2 #(.width(width)) rd_st6_1865  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1865]), .rdlo_in(a6_wr[1881]),  .coef_in(coef[576]), .rdup_out(a7_wr[1865]), .rdlo_out(a7_wr[1881]));
			radix2 #(.width(width)) rd_st6_1866  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1866]), .rdlo_in(a6_wr[1882]),  .coef_in(coef[640]), .rdup_out(a7_wr[1866]), .rdlo_out(a7_wr[1882]));
			radix2 #(.width(width)) rd_st6_1867  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1867]), .rdlo_in(a6_wr[1883]),  .coef_in(coef[704]), .rdup_out(a7_wr[1867]), .rdlo_out(a7_wr[1883]));
			radix2 #(.width(width)) rd_st6_1868  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1868]), .rdlo_in(a6_wr[1884]),  .coef_in(coef[768]), .rdup_out(a7_wr[1868]), .rdlo_out(a7_wr[1884]));
			radix2 #(.width(width)) rd_st6_1869  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1869]), .rdlo_in(a6_wr[1885]),  .coef_in(coef[832]), .rdup_out(a7_wr[1869]), .rdlo_out(a7_wr[1885]));
			radix2 #(.width(width)) rd_st6_1870  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1870]), .rdlo_in(a6_wr[1886]),  .coef_in(coef[896]), .rdup_out(a7_wr[1870]), .rdlo_out(a7_wr[1886]));
			radix2 #(.width(width)) rd_st6_1871  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1871]), .rdlo_in(a6_wr[1887]),  .coef_in(coef[960]), .rdup_out(a7_wr[1871]), .rdlo_out(a7_wr[1887]));
			radix2 #(.width(width)) rd_st6_1888  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1888]), .rdlo_in(a6_wr[1904]),  .coef_in(coef[0]), .rdup_out(a7_wr[1888]), .rdlo_out(a7_wr[1904]));
			radix2 #(.width(width)) rd_st6_1889  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1889]), .rdlo_in(a6_wr[1905]),  .coef_in(coef[64]), .rdup_out(a7_wr[1889]), .rdlo_out(a7_wr[1905]));
			radix2 #(.width(width)) rd_st6_1890  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1890]), .rdlo_in(a6_wr[1906]),  .coef_in(coef[128]), .rdup_out(a7_wr[1890]), .rdlo_out(a7_wr[1906]));
			radix2 #(.width(width)) rd_st6_1891  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1891]), .rdlo_in(a6_wr[1907]),  .coef_in(coef[192]), .rdup_out(a7_wr[1891]), .rdlo_out(a7_wr[1907]));
			radix2 #(.width(width)) rd_st6_1892  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1892]), .rdlo_in(a6_wr[1908]),  .coef_in(coef[256]), .rdup_out(a7_wr[1892]), .rdlo_out(a7_wr[1908]));
			radix2 #(.width(width)) rd_st6_1893  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1893]), .rdlo_in(a6_wr[1909]),  .coef_in(coef[320]), .rdup_out(a7_wr[1893]), .rdlo_out(a7_wr[1909]));
			radix2 #(.width(width)) rd_st6_1894  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1894]), .rdlo_in(a6_wr[1910]),  .coef_in(coef[384]), .rdup_out(a7_wr[1894]), .rdlo_out(a7_wr[1910]));
			radix2 #(.width(width)) rd_st6_1895  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1895]), .rdlo_in(a6_wr[1911]),  .coef_in(coef[448]), .rdup_out(a7_wr[1895]), .rdlo_out(a7_wr[1911]));
			radix2 #(.width(width)) rd_st6_1896  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1896]), .rdlo_in(a6_wr[1912]),  .coef_in(coef[512]), .rdup_out(a7_wr[1896]), .rdlo_out(a7_wr[1912]));
			radix2 #(.width(width)) rd_st6_1897  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1897]), .rdlo_in(a6_wr[1913]),  .coef_in(coef[576]), .rdup_out(a7_wr[1897]), .rdlo_out(a7_wr[1913]));
			radix2 #(.width(width)) rd_st6_1898  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1898]), .rdlo_in(a6_wr[1914]),  .coef_in(coef[640]), .rdup_out(a7_wr[1898]), .rdlo_out(a7_wr[1914]));
			radix2 #(.width(width)) rd_st6_1899  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1899]), .rdlo_in(a6_wr[1915]),  .coef_in(coef[704]), .rdup_out(a7_wr[1899]), .rdlo_out(a7_wr[1915]));
			radix2 #(.width(width)) rd_st6_1900  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1900]), .rdlo_in(a6_wr[1916]),  .coef_in(coef[768]), .rdup_out(a7_wr[1900]), .rdlo_out(a7_wr[1916]));
			radix2 #(.width(width)) rd_st6_1901  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1901]), .rdlo_in(a6_wr[1917]),  .coef_in(coef[832]), .rdup_out(a7_wr[1901]), .rdlo_out(a7_wr[1917]));
			radix2 #(.width(width)) rd_st6_1902  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1902]), .rdlo_in(a6_wr[1918]),  .coef_in(coef[896]), .rdup_out(a7_wr[1902]), .rdlo_out(a7_wr[1918]));
			radix2 #(.width(width)) rd_st6_1903  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1903]), .rdlo_in(a6_wr[1919]),  .coef_in(coef[960]), .rdup_out(a7_wr[1903]), .rdlo_out(a7_wr[1919]));
			radix2 #(.width(width)) rd_st6_1920  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1920]), .rdlo_in(a6_wr[1936]),  .coef_in(coef[0]), .rdup_out(a7_wr[1920]), .rdlo_out(a7_wr[1936]));
			radix2 #(.width(width)) rd_st6_1921  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1921]), .rdlo_in(a6_wr[1937]),  .coef_in(coef[64]), .rdup_out(a7_wr[1921]), .rdlo_out(a7_wr[1937]));
			radix2 #(.width(width)) rd_st6_1922  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1922]), .rdlo_in(a6_wr[1938]),  .coef_in(coef[128]), .rdup_out(a7_wr[1922]), .rdlo_out(a7_wr[1938]));
			radix2 #(.width(width)) rd_st6_1923  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1923]), .rdlo_in(a6_wr[1939]),  .coef_in(coef[192]), .rdup_out(a7_wr[1923]), .rdlo_out(a7_wr[1939]));
			radix2 #(.width(width)) rd_st6_1924  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1924]), .rdlo_in(a6_wr[1940]),  .coef_in(coef[256]), .rdup_out(a7_wr[1924]), .rdlo_out(a7_wr[1940]));
			radix2 #(.width(width)) rd_st6_1925  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1925]), .rdlo_in(a6_wr[1941]),  .coef_in(coef[320]), .rdup_out(a7_wr[1925]), .rdlo_out(a7_wr[1941]));
			radix2 #(.width(width)) rd_st6_1926  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1926]), .rdlo_in(a6_wr[1942]),  .coef_in(coef[384]), .rdup_out(a7_wr[1926]), .rdlo_out(a7_wr[1942]));
			radix2 #(.width(width)) rd_st6_1927  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1927]), .rdlo_in(a6_wr[1943]),  .coef_in(coef[448]), .rdup_out(a7_wr[1927]), .rdlo_out(a7_wr[1943]));
			radix2 #(.width(width)) rd_st6_1928  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1928]), .rdlo_in(a6_wr[1944]),  .coef_in(coef[512]), .rdup_out(a7_wr[1928]), .rdlo_out(a7_wr[1944]));
			radix2 #(.width(width)) rd_st6_1929  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1929]), .rdlo_in(a6_wr[1945]),  .coef_in(coef[576]), .rdup_out(a7_wr[1929]), .rdlo_out(a7_wr[1945]));
			radix2 #(.width(width)) rd_st6_1930  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1930]), .rdlo_in(a6_wr[1946]),  .coef_in(coef[640]), .rdup_out(a7_wr[1930]), .rdlo_out(a7_wr[1946]));
			radix2 #(.width(width)) rd_st6_1931  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1931]), .rdlo_in(a6_wr[1947]),  .coef_in(coef[704]), .rdup_out(a7_wr[1931]), .rdlo_out(a7_wr[1947]));
			radix2 #(.width(width)) rd_st6_1932  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1932]), .rdlo_in(a6_wr[1948]),  .coef_in(coef[768]), .rdup_out(a7_wr[1932]), .rdlo_out(a7_wr[1948]));
			radix2 #(.width(width)) rd_st6_1933  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1933]), .rdlo_in(a6_wr[1949]),  .coef_in(coef[832]), .rdup_out(a7_wr[1933]), .rdlo_out(a7_wr[1949]));
			radix2 #(.width(width)) rd_st6_1934  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1934]), .rdlo_in(a6_wr[1950]),  .coef_in(coef[896]), .rdup_out(a7_wr[1934]), .rdlo_out(a7_wr[1950]));
			radix2 #(.width(width)) rd_st6_1935  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1935]), .rdlo_in(a6_wr[1951]),  .coef_in(coef[960]), .rdup_out(a7_wr[1935]), .rdlo_out(a7_wr[1951]));
			radix2 #(.width(width)) rd_st6_1952  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1952]), .rdlo_in(a6_wr[1968]),  .coef_in(coef[0]), .rdup_out(a7_wr[1952]), .rdlo_out(a7_wr[1968]));
			radix2 #(.width(width)) rd_st6_1953  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1953]), .rdlo_in(a6_wr[1969]),  .coef_in(coef[64]), .rdup_out(a7_wr[1953]), .rdlo_out(a7_wr[1969]));
			radix2 #(.width(width)) rd_st6_1954  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1954]), .rdlo_in(a6_wr[1970]),  .coef_in(coef[128]), .rdup_out(a7_wr[1954]), .rdlo_out(a7_wr[1970]));
			radix2 #(.width(width)) rd_st6_1955  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1955]), .rdlo_in(a6_wr[1971]),  .coef_in(coef[192]), .rdup_out(a7_wr[1955]), .rdlo_out(a7_wr[1971]));
			radix2 #(.width(width)) rd_st6_1956  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1956]), .rdlo_in(a6_wr[1972]),  .coef_in(coef[256]), .rdup_out(a7_wr[1956]), .rdlo_out(a7_wr[1972]));
			radix2 #(.width(width)) rd_st6_1957  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1957]), .rdlo_in(a6_wr[1973]),  .coef_in(coef[320]), .rdup_out(a7_wr[1957]), .rdlo_out(a7_wr[1973]));
			radix2 #(.width(width)) rd_st6_1958  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1958]), .rdlo_in(a6_wr[1974]),  .coef_in(coef[384]), .rdup_out(a7_wr[1958]), .rdlo_out(a7_wr[1974]));
			radix2 #(.width(width)) rd_st6_1959  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1959]), .rdlo_in(a6_wr[1975]),  .coef_in(coef[448]), .rdup_out(a7_wr[1959]), .rdlo_out(a7_wr[1975]));
			radix2 #(.width(width)) rd_st6_1960  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1960]), .rdlo_in(a6_wr[1976]),  .coef_in(coef[512]), .rdup_out(a7_wr[1960]), .rdlo_out(a7_wr[1976]));
			radix2 #(.width(width)) rd_st6_1961  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1961]), .rdlo_in(a6_wr[1977]),  .coef_in(coef[576]), .rdup_out(a7_wr[1961]), .rdlo_out(a7_wr[1977]));
			radix2 #(.width(width)) rd_st6_1962  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1962]), .rdlo_in(a6_wr[1978]),  .coef_in(coef[640]), .rdup_out(a7_wr[1962]), .rdlo_out(a7_wr[1978]));
			radix2 #(.width(width)) rd_st6_1963  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1963]), .rdlo_in(a6_wr[1979]),  .coef_in(coef[704]), .rdup_out(a7_wr[1963]), .rdlo_out(a7_wr[1979]));
			radix2 #(.width(width)) rd_st6_1964  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1964]), .rdlo_in(a6_wr[1980]),  .coef_in(coef[768]), .rdup_out(a7_wr[1964]), .rdlo_out(a7_wr[1980]));
			radix2 #(.width(width)) rd_st6_1965  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1965]), .rdlo_in(a6_wr[1981]),  .coef_in(coef[832]), .rdup_out(a7_wr[1965]), .rdlo_out(a7_wr[1981]));
			radix2 #(.width(width)) rd_st6_1966  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1966]), .rdlo_in(a6_wr[1982]),  .coef_in(coef[896]), .rdup_out(a7_wr[1966]), .rdlo_out(a7_wr[1982]));
			radix2 #(.width(width)) rd_st6_1967  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1967]), .rdlo_in(a6_wr[1983]),  .coef_in(coef[960]), .rdup_out(a7_wr[1967]), .rdlo_out(a7_wr[1983]));
			radix2 #(.width(width)) rd_st6_1984  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1984]), .rdlo_in(a6_wr[2000]),  .coef_in(coef[0]), .rdup_out(a7_wr[1984]), .rdlo_out(a7_wr[2000]));
			radix2 #(.width(width)) rd_st6_1985  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1985]), .rdlo_in(a6_wr[2001]),  .coef_in(coef[64]), .rdup_out(a7_wr[1985]), .rdlo_out(a7_wr[2001]));
			radix2 #(.width(width)) rd_st6_1986  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1986]), .rdlo_in(a6_wr[2002]),  .coef_in(coef[128]), .rdup_out(a7_wr[1986]), .rdlo_out(a7_wr[2002]));
			radix2 #(.width(width)) rd_st6_1987  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1987]), .rdlo_in(a6_wr[2003]),  .coef_in(coef[192]), .rdup_out(a7_wr[1987]), .rdlo_out(a7_wr[2003]));
			radix2 #(.width(width)) rd_st6_1988  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1988]), .rdlo_in(a6_wr[2004]),  .coef_in(coef[256]), .rdup_out(a7_wr[1988]), .rdlo_out(a7_wr[2004]));
			radix2 #(.width(width)) rd_st6_1989  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1989]), .rdlo_in(a6_wr[2005]),  .coef_in(coef[320]), .rdup_out(a7_wr[1989]), .rdlo_out(a7_wr[2005]));
			radix2 #(.width(width)) rd_st6_1990  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1990]), .rdlo_in(a6_wr[2006]),  .coef_in(coef[384]), .rdup_out(a7_wr[1990]), .rdlo_out(a7_wr[2006]));
			radix2 #(.width(width)) rd_st6_1991  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1991]), .rdlo_in(a6_wr[2007]),  .coef_in(coef[448]), .rdup_out(a7_wr[1991]), .rdlo_out(a7_wr[2007]));
			radix2 #(.width(width)) rd_st6_1992  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1992]), .rdlo_in(a6_wr[2008]),  .coef_in(coef[512]), .rdup_out(a7_wr[1992]), .rdlo_out(a7_wr[2008]));
			radix2 #(.width(width)) rd_st6_1993  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1993]), .rdlo_in(a6_wr[2009]),  .coef_in(coef[576]), .rdup_out(a7_wr[1993]), .rdlo_out(a7_wr[2009]));
			radix2 #(.width(width)) rd_st6_1994  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1994]), .rdlo_in(a6_wr[2010]),  .coef_in(coef[640]), .rdup_out(a7_wr[1994]), .rdlo_out(a7_wr[2010]));
			radix2 #(.width(width)) rd_st6_1995  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1995]), .rdlo_in(a6_wr[2011]),  .coef_in(coef[704]), .rdup_out(a7_wr[1995]), .rdlo_out(a7_wr[2011]));
			radix2 #(.width(width)) rd_st6_1996  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1996]), .rdlo_in(a6_wr[2012]),  .coef_in(coef[768]), .rdup_out(a7_wr[1996]), .rdlo_out(a7_wr[2012]));
			radix2 #(.width(width)) rd_st6_1997  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1997]), .rdlo_in(a6_wr[2013]),  .coef_in(coef[832]), .rdup_out(a7_wr[1997]), .rdlo_out(a7_wr[2013]));
			radix2 #(.width(width)) rd_st6_1998  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1998]), .rdlo_in(a6_wr[2014]),  .coef_in(coef[896]), .rdup_out(a7_wr[1998]), .rdlo_out(a7_wr[2014]));
			radix2 #(.width(width)) rd_st6_1999  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[1999]), .rdlo_in(a6_wr[2015]),  .coef_in(coef[960]), .rdup_out(a7_wr[1999]), .rdlo_out(a7_wr[2015]));
			radix2 #(.width(width)) rd_st6_2016  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[2016]), .rdlo_in(a6_wr[2032]),  .coef_in(coef[0]), .rdup_out(a7_wr[2016]), .rdlo_out(a7_wr[2032]));
			radix2 #(.width(width)) rd_st6_2017  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[2017]), .rdlo_in(a6_wr[2033]),  .coef_in(coef[64]), .rdup_out(a7_wr[2017]), .rdlo_out(a7_wr[2033]));
			radix2 #(.width(width)) rd_st6_2018  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[2018]), .rdlo_in(a6_wr[2034]),  .coef_in(coef[128]), .rdup_out(a7_wr[2018]), .rdlo_out(a7_wr[2034]));
			radix2 #(.width(width)) rd_st6_2019  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[2019]), .rdlo_in(a6_wr[2035]),  .coef_in(coef[192]), .rdup_out(a7_wr[2019]), .rdlo_out(a7_wr[2035]));
			radix2 #(.width(width)) rd_st6_2020  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[2020]), .rdlo_in(a6_wr[2036]),  .coef_in(coef[256]), .rdup_out(a7_wr[2020]), .rdlo_out(a7_wr[2036]));
			radix2 #(.width(width)) rd_st6_2021  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[2021]), .rdlo_in(a6_wr[2037]),  .coef_in(coef[320]), .rdup_out(a7_wr[2021]), .rdlo_out(a7_wr[2037]));
			radix2 #(.width(width)) rd_st6_2022  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[2022]), .rdlo_in(a6_wr[2038]),  .coef_in(coef[384]), .rdup_out(a7_wr[2022]), .rdlo_out(a7_wr[2038]));
			radix2 #(.width(width)) rd_st6_2023  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[2023]), .rdlo_in(a6_wr[2039]),  .coef_in(coef[448]), .rdup_out(a7_wr[2023]), .rdlo_out(a7_wr[2039]));
			radix2 #(.width(width)) rd_st6_2024  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[2024]), .rdlo_in(a6_wr[2040]),  .coef_in(coef[512]), .rdup_out(a7_wr[2024]), .rdlo_out(a7_wr[2040]));
			radix2 #(.width(width)) rd_st6_2025  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[2025]), .rdlo_in(a6_wr[2041]),  .coef_in(coef[576]), .rdup_out(a7_wr[2025]), .rdlo_out(a7_wr[2041]));
			radix2 #(.width(width)) rd_st6_2026  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[2026]), .rdlo_in(a6_wr[2042]),  .coef_in(coef[640]), .rdup_out(a7_wr[2026]), .rdlo_out(a7_wr[2042]));
			radix2 #(.width(width)) rd_st6_2027  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[2027]), .rdlo_in(a6_wr[2043]),  .coef_in(coef[704]), .rdup_out(a7_wr[2027]), .rdlo_out(a7_wr[2043]));
			radix2 #(.width(width)) rd_st6_2028  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[2028]), .rdlo_in(a6_wr[2044]),  .coef_in(coef[768]), .rdup_out(a7_wr[2028]), .rdlo_out(a7_wr[2044]));
			radix2 #(.width(width)) rd_st6_2029  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[2029]), .rdlo_in(a6_wr[2045]),  .coef_in(coef[832]), .rdup_out(a7_wr[2029]), .rdlo_out(a7_wr[2045]));
			radix2 #(.width(width)) rd_st6_2030  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[2030]), .rdlo_in(a6_wr[2046]),  .coef_in(coef[896]), .rdup_out(a7_wr[2030]), .rdlo_out(a7_wr[2046]));
			radix2 #(.width(width)) rd_st6_2031  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a6_wr[2031]), .rdlo_in(a6_wr[2047]),  .coef_in(coef[960]), .rdup_out(a7_wr[2031]), .rdlo_out(a7_wr[2047]));

		//--- radix stage 7
			radix2 #(.width(width)) rd_st7_0   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[0]), .rdlo_in(a7_wr[8]),  .coef_in(coef[0]), .rdup_out(a8_wr[0]), .rdlo_out(a8_wr[8]));
			radix2 #(.width(width)) rd_st7_1   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1]), .rdlo_in(a7_wr[9]),  .coef_in(coef[128]), .rdup_out(a8_wr[1]), .rdlo_out(a8_wr[9]));
			radix2 #(.width(width)) rd_st7_2   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[2]), .rdlo_in(a7_wr[10]),  .coef_in(coef[256]), .rdup_out(a8_wr[2]), .rdlo_out(a8_wr[10]));
			radix2 #(.width(width)) rd_st7_3   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[3]), .rdlo_in(a7_wr[11]),  .coef_in(coef[384]), .rdup_out(a8_wr[3]), .rdlo_out(a8_wr[11]));
			radix2 #(.width(width)) rd_st7_4   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[4]), .rdlo_in(a7_wr[12]),  .coef_in(coef[512]), .rdup_out(a8_wr[4]), .rdlo_out(a8_wr[12]));
			radix2 #(.width(width)) rd_st7_5   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[5]), .rdlo_in(a7_wr[13]),  .coef_in(coef[640]), .rdup_out(a8_wr[5]), .rdlo_out(a8_wr[13]));
			radix2 #(.width(width)) rd_st7_6   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[6]), .rdlo_in(a7_wr[14]),  .coef_in(coef[768]), .rdup_out(a8_wr[6]), .rdlo_out(a8_wr[14]));
			radix2 #(.width(width)) rd_st7_7   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[7]), .rdlo_in(a7_wr[15]),  .coef_in(coef[896]), .rdup_out(a8_wr[7]), .rdlo_out(a8_wr[15]));
			radix2 #(.width(width)) rd_st7_16  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[16]), .rdlo_in(a7_wr[24]),  .coef_in(coef[0]), .rdup_out(a8_wr[16]), .rdlo_out(a8_wr[24]));
			radix2 #(.width(width)) rd_st7_17  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[17]), .rdlo_in(a7_wr[25]),  .coef_in(coef[128]), .rdup_out(a8_wr[17]), .rdlo_out(a8_wr[25]));
			radix2 #(.width(width)) rd_st7_18  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[18]), .rdlo_in(a7_wr[26]),  .coef_in(coef[256]), .rdup_out(a8_wr[18]), .rdlo_out(a8_wr[26]));
			radix2 #(.width(width)) rd_st7_19  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[19]), .rdlo_in(a7_wr[27]),  .coef_in(coef[384]), .rdup_out(a8_wr[19]), .rdlo_out(a8_wr[27]));
			radix2 #(.width(width)) rd_st7_20  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[20]), .rdlo_in(a7_wr[28]),  .coef_in(coef[512]), .rdup_out(a8_wr[20]), .rdlo_out(a8_wr[28]));
			radix2 #(.width(width)) rd_st7_21  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[21]), .rdlo_in(a7_wr[29]),  .coef_in(coef[640]), .rdup_out(a8_wr[21]), .rdlo_out(a8_wr[29]));
			radix2 #(.width(width)) rd_st7_22  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[22]), .rdlo_in(a7_wr[30]),  .coef_in(coef[768]), .rdup_out(a8_wr[22]), .rdlo_out(a8_wr[30]));
			radix2 #(.width(width)) rd_st7_23  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[23]), .rdlo_in(a7_wr[31]),  .coef_in(coef[896]), .rdup_out(a8_wr[23]), .rdlo_out(a8_wr[31]));
			radix2 #(.width(width)) rd_st7_32  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[32]), .rdlo_in(a7_wr[40]),  .coef_in(coef[0]), .rdup_out(a8_wr[32]), .rdlo_out(a8_wr[40]));
			radix2 #(.width(width)) rd_st7_33  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[33]), .rdlo_in(a7_wr[41]),  .coef_in(coef[128]), .rdup_out(a8_wr[33]), .rdlo_out(a8_wr[41]));
			radix2 #(.width(width)) rd_st7_34  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[34]), .rdlo_in(a7_wr[42]),  .coef_in(coef[256]), .rdup_out(a8_wr[34]), .rdlo_out(a8_wr[42]));
			radix2 #(.width(width)) rd_st7_35  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[35]), .rdlo_in(a7_wr[43]),  .coef_in(coef[384]), .rdup_out(a8_wr[35]), .rdlo_out(a8_wr[43]));
			radix2 #(.width(width)) rd_st7_36  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[36]), .rdlo_in(a7_wr[44]),  .coef_in(coef[512]), .rdup_out(a8_wr[36]), .rdlo_out(a8_wr[44]));
			radix2 #(.width(width)) rd_st7_37  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[37]), .rdlo_in(a7_wr[45]),  .coef_in(coef[640]), .rdup_out(a8_wr[37]), .rdlo_out(a8_wr[45]));
			radix2 #(.width(width)) rd_st7_38  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[38]), .rdlo_in(a7_wr[46]),  .coef_in(coef[768]), .rdup_out(a8_wr[38]), .rdlo_out(a8_wr[46]));
			radix2 #(.width(width)) rd_st7_39  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[39]), .rdlo_in(a7_wr[47]),  .coef_in(coef[896]), .rdup_out(a8_wr[39]), .rdlo_out(a8_wr[47]));
			radix2 #(.width(width)) rd_st7_48  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[48]), .rdlo_in(a7_wr[56]),  .coef_in(coef[0]), .rdup_out(a8_wr[48]), .rdlo_out(a8_wr[56]));
			radix2 #(.width(width)) rd_st7_49  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[49]), .rdlo_in(a7_wr[57]),  .coef_in(coef[128]), .rdup_out(a8_wr[49]), .rdlo_out(a8_wr[57]));
			radix2 #(.width(width)) rd_st7_50  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[50]), .rdlo_in(a7_wr[58]),  .coef_in(coef[256]), .rdup_out(a8_wr[50]), .rdlo_out(a8_wr[58]));
			radix2 #(.width(width)) rd_st7_51  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[51]), .rdlo_in(a7_wr[59]),  .coef_in(coef[384]), .rdup_out(a8_wr[51]), .rdlo_out(a8_wr[59]));
			radix2 #(.width(width)) rd_st7_52  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[52]), .rdlo_in(a7_wr[60]),  .coef_in(coef[512]), .rdup_out(a8_wr[52]), .rdlo_out(a8_wr[60]));
			radix2 #(.width(width)) rd_st7_53  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[53]), .rdlo_in(a7_wr[61]),  .coef_in(coef[640]), .rdup_out(a8_wr[53]), .rdlo_out(a8_wr[61]));
			radix2 #(.width(width)) rd_st7_54  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[54]), .rdlo_in(a7_wr[62]),  .coef_in(coef[768]), .rdup_out(a8_wr[54]), .rdlo_out(a8_wr[62]));
			radix2 #(.width(width)) rd_st7_55  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[55]), .rdlo_in(a7_wr[63]),  .coef_in(coef[896]), .rdup_out(a8_wr[55]), .rdlo_out(a8_wr[63]));
			radix2 #(.width(width)) rd_st7_64  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[64]), .rdlo_in(a7_wr[72]),  .coef_in(coef[0]), .rdup_out(a8_wr[64]), .rdlo_out(a8_wr[72]));
			radix2 #(.width(width)) rd_st7_65  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[65]), .rdlo_in(a7_wr[73]),  .coef_in(coef[128]), .rdup_out(a8_wr[65]), .rdlo_out(a8_wr[73]));
			radix2 #(.width(width)) rd_st7_66  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[66]), .rdlo_in(a7_wr[74]),  .coef_in(coef[256]), .rdup_out(a8_wr[66]), .rdlo_out(a8_wr[74]));
			radix2 #(.width(width)) rd_st7_67  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[67]), .rdlo_in(a7_wr[75]),  .coef_in(coef[384]), .rdup_out(a8_wr[67]), .rdlo_out(a8_wr[75]));
			radix2 #(.width(width)) rd_st7_68  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[68]), .rdlo_in(a7_wr[76]),  .coef_in(coef[512]), .rdup_out(a8_wr[68]), .rdlo_out(a8_wr[76]));
			radix2 #(.width(width)) rd_st7_69  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[69]), .rdlo_in(a7_wr[77]),  .coef_in(coef[640]), .rdup_out(a8_wr[69]), .rdlo_out(a8_wr[77]));
			radix2 #(.width(width)) rd_st7_70  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[70]), .rdlo_in(a7_wr[78]),  .coef_in(coef[768]), .rdup_out(a8_wr[70]), .rdlo_out(a8_wr[78]));
			radix2 #(.width(width)) rd_st7_71  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[71]), .rdlo_in(a7_wr[79]),  .coef_in(coef[896]), .rdup_out(a8_wr[71]), .rdlo_out(a8_wr[79]));
			radix2 #(.width(width)) rd_st7_80  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[80]), .rdlo_in(a7_wr[88]),  .coef_in(coef[0]), .rdup_out(a8_wr[80]), .rdlo_out(a8_wr[88]));
			radix2 #(.width(width)) rd_st7_81  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[81]), .rdlo_in(a7_wr[89]),  .coef_in(coef[128]), .rdup_out(a8_wr[81]), .rdlo_out(a8_wr[89]));
			radix2 #(.width(width)) rd_st7_82  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[82]), .rdlo_in(a7_wr[90]),  .coef_in(coef[256]), .rdup_out(a8_wr[82]), .rdlo_out(a8_wr[90]));
			radix2 #(.width(width)) rd_st7_83  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[83]), .rdlo_in(a7_wr[91]),  .coef_in(coef[384]), .rdup_out(a8_wr[83]), .rdlo_out(a8_wr[91]));
			radix2 #(.width(width)) rd_st7_84  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[84]), .rdlo_in(a7_wr[92]),  .coef_in(coef[512]), .rdup_out(a8_wr[84]), .rdlo_out(a8_wr[92]));
			radix2 #(.width(width)) rd_st7_85  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[85]), .rdlo_in(a7_wr[93]),  .coef_in(coef[640]), .rdup_out(a8_wr[85]), .rdlo_out(a8_wr[93]));
			radix2 #(.width(width)) rd_st7_86  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[86]), .rdlo_in(a7_wr[94]),  .coef_in(coef[768]), .rdup_out(a8_wr[86]), .rdlo_out(a8_wr[94]));
			radix2 #(.width(width)) rd_st7_87  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[87]), .rdlo_in(a7_wr[95]),  .coef_in(coef[896]), .rdup_out(a8_wr[87]), .rdlo_out(a8_wr[95]));
			radix2 #(.width(width)) rd_st7_96  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[96]), .rdlo_in(a7_wr[104]),  .coef_in(coef[0]), .rdup_out(a8_wr[96]), .rdlo_out(a8_wr[104]));
			radix2 #(.width(width)) rd_st7_97  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[97]), .rdlo_in(a7_wr[105]),  .coef_in(coef[128]), .rdup_out(a8_wr[97]), .rdlo_out(a8_wr[105]));
			radix2 #(.width(width)) rd_st7_98  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[98]), .rdlo_in(a7_wr[106]),  .coef_in(coef[256]), .rdup_out(a8_wr[98]), .rdlo_out(a8_wr[106]));
			radix2 #(.width(width)) rd_st7_99  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[99]), .rdlo_in(a7_wr[107]),  .coef_in(coef[384]), .rdup_out(a8_wr[99]), .rdlo_out(a8_wr[107]));
			radix2 #(.width(width)) rd_st7_100  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[100]), .rdlo_in(a7_wr[108]),  .coef_in(coef[512]), .rdup_out(a8_wr[100]), .rdlo_out(a8_wr[108]));
			radix2 #(.width(width)) rd_st7_101  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[101]), .rdlo_in(a7_wr[109]),  .coef_in(coef[640]), .rdup_out(a8_wr[101]), .rdlo_out(a8_wr[109]));
			radix2 #(.width(width)) rd_st7_102  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[102]), .rdlo_in(a7_wr[110]),  .coef_in(coef[768]), .rdup_out(a8_wr[102]), .rdlo_out(a8_wr[110]));
			radix2 #(.width(width)) rd_st7_103  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[103]), .rdlo_in(a7_wr[111]),  .coef_in(coef[896]), .rdup_out(a8_wr[103]), .rdlo_out(a8_wr[111]));
			radix2 #(.width(width)) rd_st7_112  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[112]), .rdlo_in(a7_wr[120]),  .coef_in(coef[0]), .rdup_out(a8_wr[112]), .rdlo_out(a8_wr[120]));
			radix2 #(.width(width)) rd_st7_113  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[113]), .rdlo_in(a7_wr[121]),  .coef_in(coef[128]), .rdup_out(a8_wr[113]), .rdlo_out(a8_wr[121]));
			radix2 #(.width(width)) rd_st7_114  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[114]), .rdlo_in(a7_wr[122]),  .coef_in(coef[256]), .rdup_out(a8_wr[114]), .rdlo_out(a8_wr[122]));
			radix2 #(.width(width)) rd_st7_115  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[115]), .rdlo_in(a7_wr[123]),  .coef_in(coef[384]), .rdup_out(a8_wr[115]), .rdlo_out(a8_wr[123]));
			radix2 #(.width(width)) rd_st7_116  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[116]), .rdlo_in(a7_wr[124]),  .coef_in(coef[512]), .rdup_out(a8_wr[116]), .rdlo_out(a8_wr[124]));
			radix2 #(.width(width)) rd_st7_117  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[117]), .rdlo_in(a7_wr[125]),  .coef_in(coef[640]), .rdup_out(a8_wr[117]), .rdlo_out(a8_wr[125]));
			radix2 #(.width(width)) rd_st7_118  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[118]), .rdlo_in(a7_wr[126]),  .coef_in(coef[768]), .rdup_out(a8_wr[118]), .rdlo_out(a8_wr[126]));
			radix2 #(.width(width)) rd_st7_119  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[119]), .rdlo_in(a7_wr[127]),  .coef_in(coef[896]), .rdup_out(a8_wr[119]), .rdlo_out(a8_wr[127]));
			radix2 #(.width(width)) rd_st7_128  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[128]), .rdlo_in(a7_wr[136]),  .coef_in(coef[0]), .rdup_out(a8_wr[128]), .rdlo_out(a8_wr[136]));
			radix2 #(.width(width)) rd_st7_129  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[129]), .rdlo_in(a7_wr[137]),  .coef_in(coef[128]), .rdup_out(a8_wr[129]), .rdlo_out(a8_wr[137]));
			radix2 #(.width(width)) rd_st7_130  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[130]), .rdlo_in(a7_wr[138]),  .coef_in(coef[256]), .rdup_out(a8_wr[130]), .rdlo_out(a8_wr[138]));
			radix2 #(.width(width)) rd_st7_131  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[131]), .rdlo_in(a7_wr[139]),  .coef_in(coef[384]), .rdup_out(a8_wr[131]), .rdlo_out(a8_wr[139]));
			radix2 #(.width(width)) rd_st7_132  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[132]), .rdlo_in(a7_wr[140]),  .coef_in(coef[512]), .rdup_out(a8_wr[132]), .rdlo_out(a8_wr[140]));
			radix2 #(.width(width)) rd_st7_133  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[133]), .rdlo_in(a7_wr[141]),  .coef_in(coef[640]), .rdup_out(a8_wr[133]), .rdlo_out(a8_wr[141]));
			radix2 #(.width(width)) rd_st7_134  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[134]), .rdlo_in(a7_wr[142]),  .coef_in(coef[768]), .rdup_out(a8_wr[134]), .rdlo_out(a8_wr[142]));
			radix2 #(.width(width)) rd_st7_135  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[135]), .rdlo_in(a7_wr[143]),  .coef_in(coef[896]), .rdup_out(a8_wr[135]), .rdlo_out(a8_wr[143]));
			radix2 #(.width(width)) rd_st7_144  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[144]), .rdlo_in(a7_wr[152]),  .coef_in(coef[0]), .rdup_out(a8_wr[144]), .rdlo_out(a8_wr[152]));
			radix2 #(.width(width)) rd_st7_145  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[145]), .rdlo_in(a7_wr[153]),  .coef_in(coef[128]), .rdup_out(a8_wr[145]), .rdlo_out(a8_wr[153]));
			radix2 #(.width(width)) rd_st7_146  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[146]), .rdlo_in(a7_wr[154]),  .coef_in(coef[256]), .rdup_out(a8_wr[146]), .rdlo_out(a8_wr[154]));
			radix2 #(.width(width)) rd_st7_147  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[147]), .rdlo_in(a7_wr[155]),  .coef_in(coef[384]), .rdup_out(a8_wr[147]), .rdlo_out(a8_wr[155]));
			radix2 #(.width(width)) rd_st7_148  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[148]), .rdlo_in(a7_wr[156]),  .coef_in(coef[512]), .rdup_out(a8_wr[148]), .rdlo_out(a8_wr[156]));
			radix2 #(.width(width)) rd_st7_149  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[149]), .rdlo_in(a7_wr[157]),  .coef_in(coef[640]), .rdup_out(a8_wr[149]), .rdlo_out(a8_wr[157]));
			radix2 #(.width(width)) rd_st7_150  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[150]), .rdlo_in(a7_wr[158]),  .coef_in(coef[768]), .rdup_out(a8_wr[150]), .rdlo_out(a8_wr[158]));
			radix2 #(.width(width)) rd_st7_151  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[151]), .rdlo_in(a7_wr[159]),  .coef_in(coef[896]), .rdup_out(a8_wr[151]), .rdlo_out(a8_wr[159]));
			radix2 #(.width(width)) rd_st7_160  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[160]), .rdlo_in(a7_wr[168]),  .coef_in(coef[0]), .rdup_out(a8_wr[160]), .rdlo_out(a8_wr[168]));
			radix2 #(.width(width)) rd_st7_161  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[161]), .rdlo_in(a7_wr[169]),  .coef_in(coef[128]), .rdup_out(a8_wr[161]), .rdlo_out(a8_wr[169]));
			radix2 #(.width(width)) rd_st7_162  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[162]), .rdlo_in(a7_wr[170]),  .coef_in(coef[256]), .rdup_out(a8_wr[162]), .rdlo_out(a8_wr[170]));
			radix2 #(.width(width)) rd_st7_163  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[163]), .rdlo_in(a7_wr[171]),  .coef_in(coef[384]), .rdup_out(a8_wr[163]), .rdlo_out(a8_wr[171]));
			radix2 #(.width(width)) rd_st7_164  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[164]), .rdlo_in(a7_wr[172]),  .coef_in(coef[512]), .rdup_out(a8_wr[164]), .rdlo_out(a8_wr[172]));
			radix2 #(.width(width)) rd_st7_165  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[165]), .rdlo_in(a7_wr[173]),  .coef_in(coef[640]), .rdup_out(a8_wr[165]), .rdlo_out(a8_wr[173]));
			radix2 #(.width(width)) rd_st7_166  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[166]), .rdlo_in(a7_wr[174]),  .coef_in(coef[768]), .rdup_out(a8_wr[166]), .rdlo_out(a8_wr[174]));
			radix2 #(.width(width)) rd_st7_167  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[167]), .rdlo_in(a7_wr[175]),  .coef_in(coef[896]), .rdup_out(a8_wr[167]), .rdlo_out(a8_wr[175]));
			radix2 #(.width(width)) rd_st7_176  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[176]), .rdlo_in(a7_wr[184]),  .coef_in(coef[0]), .rdup_out(a8_wr[176]), .rdlo_out(a8_wr[184]));
			radix2 #(.width(width)) rd_st7_177  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[177]), .rdlo_in(a7_wr[185]),  .coef_in(coef[128]), .rdup_out(a8_wr[177]), .rdlo_out(a8_wr[185]));
			radix2 #(.width(width)) rd_st7_178  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[178]), .rdlo_in(a7_wr[186]),  .coef_in(coef[256]), .rdup_out(a8_wr[178]), .rdlo_out(a8_wr[186]));
			radix2 #(.width(width)) rd_st7_179  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[179]), .rdlo_in(a7_wr[187]),  .coef_in(coef[384]), .rdup_out(a8_wr[179]), .rdlo_out(a8_wr[187]));
			radix2 #(.width(width)) rd_st7_180  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[180]), .rdlo_in(a7_wr[188]),  .coef_in(coef[512]), .rdup_out(a8_wr[180]), .rdlo_out(a8_wr[188]));
			radix2 #(.width(width)) rd_st7_181  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[181]), .rdlo_in(a7_wr[189]),  .coef_in(coef[640]), .rdup_out(a8_wr[181]), .rdlo_out(a8_wr[189]));
			radix2 #(.width(width)) rd_st7_182  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[182]), .rdlo_in(a7_wr[190]),  .coef_in(coef[768]), .rdup_out(a8_wr[182]), .rdlo_out(a8_wr[190]));
			radix2 #(.width(width)) rd_st7_183  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[183]), .rdlo_in(a7_wr[191]),  .coef_in(coef[896]), .rdup_out(a8_wr[183]), .rdlo_out(a8_wr[191]));
			radix2 #(.width(width)) rd_st7_192  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[192]), .rdlo_in(a7_wr[200]),  .coef_in(coef[0]), .rdup_out(a8_wr[192]), .rdlo_out(a8_wr[200]));
			radix2 #(.width(width)) rd_st7_193  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[193]), .rdlo_in(a7_wr[201]),  .coef_in(coef[128]), .rdup_out(a8_wr[193]), .rdlo_out(a8_wr[201]));
			radix2 #(.width(width)) rd_st7_194  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[194]), .rdlo_in(a7_wr[202]),  .coef_in(coef[256]), .rdup_out(a8_wr[194]), .rdlo_out(a8_wr[202]));
			radix2 #(.width(width)) rd_st7_195  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[195]), .rdlo_in(a7_wr[203]),  .coef_in(coef[384]), .rdup_out(a8_wr[195]), .rdlo_out(a8_wr[203]));
			radix2 #(.width(width)) rd_st7_196  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[196]), .rdlo_in(a7_wr[204]),  .coef_in(coef[512]), .rdup_out(a8_wr[196]), .rdlo_out(a8_wr[204]));
			radix2 #(.width(width)) rd_st7_197  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[197]), .rdlo_in(a7_wr[205]),  .coef_in(coef[640]), .rdup_out(a8_wr[197]), .rdlo_out(a8_wr[205]));
			radix2 #(.width(width)) rd_st7_198  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[198]), .rdlo_in(a7_wr[206]),  .coef_in(coef[768]), .rdup_out(a8_wr[198]), .rdlo_out(a8_wr[206]));
			radix2 #(.width(width)) rd_st7_199  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[199]), .rdlo_in(a7_wr[207]),  .coef_in(coef[896]), .rdup_out(a8_wr[199]), .rdlo_out(a8_wr[207]));
			radix2 #(.width(width)) rd_st7_208  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[208]), .rdlo_in(a7_wr[216]),  .coef_in(coef[0]), .rdup_out(a8_wr[208]), .rdlo_out(a8_wr[216]));
			radix2 #(.width(width)) rd_st7_209  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[209]), .rdlo_in(a7_wr[217]),  .coef_in(coef[128]), .rdup_out(a8_wr[209]), .rdlo_out(a8_wr[217]));
			radix2 #(.width(width)) rd_st7_210  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[210]), .rdlo_in(a7_wr[218]),  .coef_in(coef[256]), .rdup_out(a8_wr[210]), .rdlo_out(a8_wr[218]));
			radix2 #(.width(width)) rd_st7_211  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[211]), .rdlo_in(a7_wr[219]),  .coef_in(coef[384]), .rdup_out(a8_wr[211]), .rdlo_out(a8_wr[219]));
			radix2 #(.width(width)) rd_st7_212  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[212]), .rdlo_in(a7_wr[220]),  .coef_in(coef[512]), .rdup_out(a8_wr[212]), .rdlo_out(a8_wr[220]));
			radix2 #(.width(width)) rd_st7_213  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[213]), .rdlo_in(a7_wr[221]),  .coef_in(coef[640]), .rdup_out(a8_wr[213]), .rdlo_out(a8_wr[221]));
			radix2 #(.width(width)) rd_st7_214  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[214]), .rdlo_in(a7_wr[222]),  .coef_in(coef[768]), .rdup_out(a8_wr[214]), .rdlo_out(a8_wr[222]));
			radix2 #(.width(width)) rd_st7_215  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[215]), .rdlo_in(a7_wr[223]),  .coef_in(coef[896]), .rdup_out(a8_wr[215]), .rdlo_out(a8_wr[223]));
			radix2 #(.width(width)) rd_st7_224  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[224]), .rdlo_in(a7_wr[232]),  .coef_in(coef[0]), .rdup_out(a8_wr[224]), .rdlo_out(a8_wr[232]));
			radix2 #(.width(width)) rd_st7_225  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[225]), .rdlo_in(a7_wr[233]),  .coef_in(coef[128]), .rdup_out(a8_wr[225]), .rdlo_out(a8_wr[233]));
			radix2 #(.width(width)) rd_st7_226  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[226]), .rdlo_in(a7_wr[234]),  .coef_in(coef[256]), .rdup_out(a8_wr[226]), .rdlo_out(a8_wr[234]));
			radix2 #(.width(width)) rd_st7_227  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[227]), .rdlo_in(a7_wr[235]),  .coef_in(coef[384]), .rdup_out(a8_wr[227]), .rdlo_out(a8_wr[235]));
			radix2 #(.width(width)) rd_st7_228  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[228]), .rdlo_in(a7_wr[236]),  .coef_in(coef[512]), .rdup_out(a8_wr[228]), .rdlo_out(a8_wr[236]));
			radix2 #(.width(width)) rd_st7_229  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[229]), .rdlo_in(a7_wr[237]),  .coef_in(coef[640]), .rdup_out(a8_wr[229]), .rdlo_out(a8_wr[237]));
			radix2 #(.width(width)) rd_st7_230  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[230]), .rdlo_in(a7_wr[238]),  .coef_in(coef[768]), .rdup_out(a8_wr[230]), .rdlo_out(a8_wr[238]));
			radix2 #(.width(width)) rd_st7_231  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[231]), .rdlo_in(a7_wr[239]),  .coef_in(coef[896]), .rdup_out(a8_wr[231]), .rdlo_out(a8_wr[239]));
			radix2 #(.width(width)) rd_st7_240  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[240]), .rdlo_in(a7_wr[248]),  .coef_in(coef[0]), .rdup_out(a8_wr[240]), .rdlo_out(a8_wr[248]));
			radix2 #(.width(width)) rd_st7_241  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[241]), .rdlo_in(a7_wr[249]),  .coef_in(coef[128]), .rdup_out(a8_wr[241]), .rdlo_out(a8_wr[249]));
			radix2 #(.width(width)) rd_st7_242  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[242]), .rdlo_in(a7_wr[250]),  .coef_in(coef[256]), .rdup_out(a8_wr[242]), .rdlo_out(a8_wr[250]));
			radix2 #(.width(width)) rd_st7_243  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[243]), .rdlo_in(a7_wr[251]),  .coef_in(coef[384]), .rdup_out(a8_wr[243]), .rdlo_out(a8_wr[251]));
			radix2 #(.width(width)) rd_st7_244  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[244]), .rdlo_in(a7_wr[252]),  .coef_in(coef[512]), .rdup_out(a8_wr[244]), .rdlo_out(a8_wr[252]));
			radix2 #(.width(width)) rd_st7_245  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[245]), .rdlo_in(a7_wr[253]),  .coef_in(coef[640]), .rdup_out(a8_wr[245]), .rdlo_out(a8_wr[253]));
			radix2 #(.width(width)) rd_st7_246  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[246]), .rdlo_in(a7_wr[254]),  .coef_in(coef[768]), .rdup_out(a8_wr[246]), .rdlo_out(a8_wr[254]));
			radix2 #(.width(width)) rd_st7_247  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[247]), .rdlo_in(a7_wr[255]),  .coef_in(coef[896]), .rdup_out(a8_wr[247]), .rdlo_out(a8_wr[255]));
			radix2 #(.width(width)) rd_st7_256  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[256]), .rdlo_in(a7_wr[264]),  .coef_in(coef[0]), .rdup_out(a8_wr[256]), .rdlo_out(a8_wr[264]));
			radix2 #(.width(width)) rd_st7_257  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[257]), .rdlo_in(a7_wr[265]),  .coef_in(coef[128]), .rdup_out(a8_wr[257]), .rdlo_out(a8_wr[265]));
			radix2 #(.width(width)) rd_st7_258  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[258]), .rdlo_in(a7_wr[266]),  .coef_in(coef[256]), .rdup_out(a8_wr[258]), .rdlo_out(a8_wr[266]));
			radix2 #(.width(width)) rd_st7_259  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[259]), .rdlo_in(a7_wr[267]),  .coef_in(coef[384]), .rdup_out(a8_wr[259]), .rdlo_out(a8_wr[267]));
			radix2 #(.width(width)) rd_st7_260  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[260]), .rdlo_in(a7_wr[268]),  .coef_in(coef[512]), .rdup_out(a8_wr[260]), .rdlo_out(a8_wr[268]));
			radix2 #(.width(width)) rd_st7_261  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[261]), .rdlo_in(a7_wr[269]),  .coef_in(coef[640]), .rdup_out(a8_wr[261]), .rdlo_out(a8_wr[269]));
			radix2 #(.width(width)) rd_st7_262  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[262]), .rdlo_in(a7_wr[270]),  .coef_in(coef[768]), .rdup_out(a8_wr[262]), .rdlo_out(a8_wr[270]));
			radix2 #(.width(width)) rd_st7_263  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[263]), .rdlo_in(a7_wr[271]),  .coef_in(coef[896]), .rdup_out(a8_wr[263]), .rdlo_out(a8_wr[271]));
			radix2 #(.width(width)) rd_st7_272  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[272]), .rdlo_in(a7_wr[280]),  .coef_in(coef[0]), .rdup_out(a8_wr[272]), .rdlo_out(a8_wr[280]));
			radix2 #(.width(width)) rd_st7_273  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[273]), .rdlo_in(a7_wr[281]),  .coef_in(coef[128]), .rdup_out(a8_wr[273]), .rdlo_out(a8_wr[281]));
			radix2 #(.width(width)) rd_st7_274  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[274]), .rdlo_in(a7_wr[282]),  .coef_in(coef[256]), .rdup_out(a8_wr[274]), .rdlo_out(a8_wr[282]));
			radix2 #(.width(width)) rd_st7_275  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[275]), .rdlo_in(a7_wr[283]),  .coef_in(coef[384]), .rdup_out(a8_wr[275]), .rdlo_out(a8_wr[283]));
			radix2 #(.width(width)) rd_st7_276  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[276]), .rdlo_in(a7_wr[284]),  .coef_in(coef[512]), .rdup_out(a8_wr[276]), .rdlo_out(a8_wr[284]));
			radix2 #(.width(width)) rd_st7_277  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[277]), .rdlo_in(a7_wr[285]),  .coef_in(coef[640]), .rdup_out(a8_wr[277]), .rdlo_out(a8_wr[285]));
			radix2 #(.width(width)) rd_st7_278  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[278]), .rdlo_in(a7_wr[286]),  .coef_in(coef[768]), .rdup_out(a8_wr[278]), .rdlo_out(a8_wr[286]));
			radix2 #(.width(width)) rd_st7_279  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[279]), .rdlo_in(a7_wr[287]),  .coef_in(coef[896]), .rdup_out(a8_wr[279]), .rdlo_out(a8_wr[287]));
			radix2 #(.width(width)) rd_st7_288  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[288]), .rdlo_in(a7_wr[296]),  .coef_in(coef[0]), .rdup_out(a8_wr[288]), .rdlo_out(a8_wr[296]));
			radix2 #(.width(width)) rd_st7_289  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[289]), .rdlo_in(a7_wr[297]),  .coef_in(coef[128]), .rdup_out(a8_wr[289]), .rdlo_out(a8_wr[297]));
			radix2 #(.width(width)) rd_st7_290  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[290]), .rdlo_in(a7_wr[298]),  .coef_in(coef[256]), .rdup_out(a8_wr[290]), .rdlo_out(a8_wr[298]));
			radix2 #(.width(width)) rd_st7_291  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[291]), .rdlo_in(a7_wr[299]),  .coef_in(coef[384]), .rdup_out(a8_wr[291]), .rdlo_out(a8_wr[299]));
			radix2 #(.width(width)) rd_st7_292  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[292]), .rdlo_in(a7_wr[300]),  .coef_in(coef[512]), .rdup_out(a8_wr[292]), .rdlo_out(a8_wr[300]));
			radix2 #(.width(width)) rd_st7_293  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[293]), .rdlo_in(a7_wr[301]),  .coef_in(coef[640]), .rdup_out(a8_wr[293]), .rdlo_out(a8_wr[301]));
			radix2 #(.width(width)) rd_st7_294  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[294]), .rdlo_in(a7_wr[302]),  .coef_in(coef[768]), .rdup_out(a8_wr[294]), .rdlo_out(a8_wr[302]));
			radix2 #(.width(width)) rd_st7_295  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[295]), .rdlo_in(a7_wr[303]),  .coef_in(coef[896]), .rdup_out(a8_wr[295]), .rdlo_out(a8_wr[303]));
			radix2 #(.width(width)) rd_st7_304  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[304]), .rdlo_in(a7_wr[312]),  .coef_in(coef[0]), .rdup_out(a8_wr[304]), .rdlo_out(a8_wr[312]));
			radix2 #(.width(width)) rd_st7_305  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[305]), .rdlo_in(a7_wr[313]),  .coef_in(coef[128]), .rdup_out(a8_wr[305]), .rdlo_out(a8_wr[313]));
			radix2 #(.width(width)) rd_st7_306  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[306]), .rdlo_in(a7_wr[314]),  .coef_in(coef[256]), .rdup_out(a8_wr[306]), .rdlo_out(a8_wr[314]));
			radix2 #(.width(width)) rd_st7_307  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[307]), .rdlo_in(a7_wr[315]),  .coef_in(coef[384]), .rdup_out(a8_wr[307]), .rdlo_out(a8_wr[315]));
			radix2 #(.width(width)) rd_st7_308  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[308]), .rdlo_in(a7_wr[316]),  .coef_in(coef[512]), .rdup_out(a8_wr[308]), .rdlo_out(a8_wr[316]));
			radix2 #(.width(width)) rd_st7_309  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[309]), .rdlo_in(a7_wr[317]),  .coef_in(coef[640]), .rdup_out(a8_wr[309]), .rdlo_out(a8_wr[317]));
			radix2 #(.width(width)) rd_st7_310  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[310]), .rdlo_in(a7_wr[318]),  .coef_in(coef[768]), .rdup_out(a8_wr[310]), .rdlo_out(a8_wr[318]));
			radix2 #(.width(width)) rd_st7_311  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[311]), .rdlo_in(a7_wr[319]),  .coef_in(coef[896]), .rdup_out(a8_wr[311]), .rdlo_out(a8_wr[319]));
			radix2 #(.width(width)) rd_st7_320  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[320]), .rdlo_in(a7_wr[328]),  .coef_in(coef[0]), .rdup_out(a8_wr[320]), .rdlo_out(a8_wr[328]));
			radix2 #(.width(width)) rd_st7_321  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[321]), .rdlo_in(a7_wr[329]),  .coef_in(coef[128]), .rdup_out(a8_wr[321]), .rdlo_out(a8_wr[329]));
			radix2 #(.width(width)) rd_st7_322  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[322]), .rdlo_in(a7_wr[330]),  .coef_in(coef[256]), .rdup_out(a8_wr[322]), .rdlo_out(a8_wr[330]));
			radix2 #(.width(width)) rd_st7_323  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[323]), .rdlo_in(a7_wr[331]),  .coef_in(coef[384]), .rdup_out(a8_wr[323]), .rdlo_out(a8_wr[331]));
			radix2 #(.width(width)) rd_st7_324  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[324]), .rdlo_in(a7_wr[332]),  .coef_in(coef[512]), .rdup_out(a8_wr[324]), .rdlo_out(a8_wr[332]));
			radix2 #(.width(width)) rd_st7_325  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[325]), .rdlo_in(a7_wr[333]),  .coef_in(coef[640]), .rdup_out(a8_wr[325]), .rdlo_out(a8_wr[333]));
			radix2 #(.width(width)) rd_st7_326  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[326]), .rdlo_in(a7_wr[334]),  .coef_in(coef[768]), .rdup_out(a8_wr[326]), .rdlo_out(a8_wr[334]));
			radix2 #(.width(width)) rd_st7_327  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[327]), .rdlo_in(a7_wr[335]),  .coef_in(coef[896]), .rdup_out(a8_wr[327]), .rdlo_out(a8_wr[335]));
			radix2 #(.width(width)) rd_st7_336  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[336]), .rdlo_in(a7_wr[344]),  .coef_in(coef[0]), .rdup_out(a8_wr[336]), .rdlo_out(a8_wr[344]));
			radix2 #(.width(width)) rd_st7_337  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[337]), .rdlo_in(a7_wr[345]),  .coef_in(coef[128]), .rdup_out(a8_wr[337]), .rdlo_out(a8_wr[345]));
			radix2 #(.width(width)) rd_st7_338  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[338]), .rdlo_in(a7_wr[346]),  .coef_in(coef[256]), .rdup_out(a8_wr[338]), .rdlo_out(a8_wr[346]));
			radix2 #(.width(width)) rd_st7_339  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[339]), .rdlo_in(a7_wr[347]),  .coef_in(coef[384]), .rdup_out(a8_wr[339]), .rdlo_out(a8_wr[347]));
			radix2 #(.width(width)) rd_st7_340  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[340]), .rdlo_in(a7_wr[348]),  .coef_in(coef[512]), .rdup_out(a8_wr[340]), .rdlo_out(a8_wr[348]));
			radix2 #(.width(width)) rd_st7_341  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[341]), .rdlo_in(a7_wr[349]),  .coef_in(coef[640]), .rdup_out(a8_wr[341]), .rdlo_out(a8_wr[349]));
			radix2 #(.width(width)) rd_st7_342  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[342]), .rdlo_in(a7_wr[350]),  .coef_in(coef[768]), .rdup_out(a8_wr[342]), .rdlo_out(a8_wr[350]));
			radix2 #(.width(width)) rd_st7_343  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[343]), .rdlo_in(a7_wr[351]),  .coef_in(coef[896]), .rdup_out(a8_wr[343]), .rdlo_out(a8_wr[351]));
			radix2 #(.width(width)) rd_st7_352  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[352]), .rdlo_in(a7_wr[360]),  .coef_in(coef[0]), .rdup_out(a8_wr[352]), .rdlo_out(a8_wr[360]));
			radix2 #(.width(width)) rd_st7_353  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[353]), .rdlo_in(a7_wr[361]),  .coef_in(coef[128]), .rdup_out(a8_wr[353]), .rdlo_out(a8_wr[361]));
			radix2 #(.width(width)) rd_st7_354  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[354]), .rdlo_in(a7_wr[362]),  .coef_in(coef[256]), .rdup_out(a8_wr[354]), .rdlo_out(a8_wr[362]));
			radix2 #(.width(width)) rd_st7_355  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[355]), .rdlo_in(a7_wr[363]),  .coef_in(coef[384]), .rdup_out(a8_wr[355]), .rdlo_out(a8_wr[363]));
			radix2 #(.width(width)) rd_st7_356  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[356]), .rdlo_in(a7_wr[364]),  .coef_in(coef[512]), .rdup_out(a8_wr[356]), .rdlo_out(a8_wr[364]));
			radix2 #(.width(width)) rd_st7_357  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[357]), .rdlo_in(a7_wr[365]),  .coef_in(coef[640]), .rdup_out(a8_wr[357]), .rdlo_out(a8_wr[365]));
			radix2 #(.width(width)) rd_st7_358  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[358]), .rdlo_in(a7_wr[366]),  .coef_in(coef[768]), .rdup_out(a8_wr[358]), .rdlo_out(a8_wr[366]));
			radix2 #(.width(width)) rd_st7_359  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[359]), .rdlo_in(a7_wr[367]),  .coef_in(coef[896]), .rdup_out(a8_wr[359]), .rdlo_out(a8_wr[367]));
			radix2 #(.width(width)) rd_st7_368  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[368]), .rdlo_in(a7_wr[376]),  .coef_in(coef[0]), .rdup_out(a8_wr[368]), .rdlo_out(a8_wr[376]));
			radix2 #(.width(width)) rd_st7_369  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[369]), .rdlo_in(a7_wr[377]),  .coef_in(coef[128]), .rdup_out(a8_wr[369]), .rdlo_out(a8_wr[377]));
			radix2 #(.width(width)) rd_st7_370  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[370]), .rdlo_in(a7_wr[378]),  .coef_in(coef[256]), .rdup_out(a8_wr[370]), .rdlo_out(a8_wr[378]));
			radix2 #(.width(width)) rd_st7_371  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[371]), .rdlo_in(a7_wr[379]),  .coef_in(coef[384]), .rdup_out(a8_wr[371]), .rdlo_out(a8_wr[379]));
			radix2 #(.width(width)) rd_st7_372  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[372]), .rdlo_in(a7_wr[380]),  .coef_in(coef[512]), .rdup_out(a8_wr[372]), .rdlo_out(a8_wr[380]));
			radix2 #(.width(width)) rd_st7_373  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[373]), .rdlo_in(a7_wr[381]),  .coef_in(coef[640]), .rdup_out(a8_wr[373]), .rdlo_out(a8_wr[381]));
			radix2 #(.width(width)) rd_st7_374  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[374]), .rdlo_in(a7_wr[382]),  .coef_in(coef[768]), .rdup_out(a8_wr[374]), .rdlo_out(a8_wr[382]));
			radix2 #(.width(width)) rd_st7_375  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[375]), .rdlo_in(a7_wr[383]),  .coef_in(coef[896]), .rdup_out(a8_wr[375]), .rdlo_out(a8_wr[383]));
			radix2 #(.width(width)) rd_st7_384  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[384]), .rdlo_in(a7_wr[392]),  .coef_in(coef[0]), .rdup_out(a8_wr[384]), .rdlo_out(a8_wr[392]));
			radix2 #(.width(width)) rd_st7_385  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[385]), .rdlo_in(a7_wr[393]),  .coef_in(coef[128]), .rdup_out(a8_wr[385]), .rdlo_out(a8_wr[393]));
			radix2 #(.width(width)) rd_st7_386  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[386]), .rdlo_in(a7_wr[394]),  .coef_in(coef[256]), .rdup_out(a8_wr[386]), .rdlo_out(a8_wr[394]));
			radix2 #(.width(width)) rd_st7_387  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[387]), .rdlo_in(a7_wr[395]),  .coef_in(coef[384]), .rdup_out(a8_wr[387]), .rdlo_out(a8_wr[395]));
			radix2 #(.width(width)) rd_st7_388  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[388]), .rdlo_in(a7_wr[396]),  .coef_in(coef[512]), .rdup_out(a8_wr[388]), .rdlo_out(a8_wr[396]));
			radix2 #(.width(width)) rd_st7_389  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[389]), .rdlo_in(a7_wr[397]),  .coef_in(coef[640]), .rdup_out(a8_wr[389]), .rdlo_out(a8_wr[397]));
			radix2 #(.width(width)) rd_st7_390  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[390]), .rdlo_in(a7_wr[398]),  .coef_in(coef[768]), .rdup_out(a8_wr[390]), .rdlo_out(a8_wr[398]));
			radix2 #(.width(width)) rd_st7_391  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[391]), .rdlo_in(a7_wr[399]),  .coef_in(coef[896]), .rdup_out(a8_wr[391]), .rdlo_out(a8_wr[399]));
			radix2 #(.width(width)) rd_st7_400  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[400]), .rdlo_in(a7_wr[408]),  .coef_in(coef[0]), .rdup_out(a8_wr[400]), .rdlo_out(a8_wr[408]));
			radix2 #(.width(width)) rd_st7_401  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[401]), .rdlo_in(a7_wr[409]),  .coef_in(coef[128]), .rdup_out(a8_wr[401]), .rdlo_out(a8_wr[409]));
			radix2 #(.width(width)) rd_st7_402  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[402]), .rdlo_in(a7_wr[410]),  .coef_in(coef[256]), .rdup_out(a8_wr[402]), .rdlo_out(a8_wr[410]));
			radix2 #(.width(width)) rd_st7_403  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[403]), .rdlo_in(a7_wr[411]),  .coef_in(coef[384]), .rdup_out(a8_wr[403]), .rdlo_out(a8_wr[411]));
			radix2 #(.width(width)) rd_st7_404  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[404]), .rdlo_in(a7_wr[412]),  .coef_in(coef[512]), .rdup_out(a8_wr[404]), .rdlo_out(a8_wr[412]));
			radix2 #(.width(width)) rd_st7_405  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[405]), .rdlo_in(a7_wr[413]),  .coef_in(coef[640]), .rdup_out(a8_wr[405]), .rdlo_out(a8_wr[413]));
			radix2 #(.width(width)) rd_st7_406  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[406]), .rdlo_in(a7_wr[414]),  .coef_in(coef[768]), .rdup_out(a8_wr[406]), .rdlo_out(a8_wr[414]));
			radix2 #(.width(width)) rd_st7_407  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[407]), .rdlo_in(a7_wr[415]),  .coef_in(coef[896]), .rdup_out(a8_wr[407]), .rdlo_out(a8_wr[415]));
			radix2 #(.width(width)) rd_st7_416  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[416]), .rdlo_in(a7_wr[424]),  .coef_in(coef[0]), .rdup_out(a8_wr[416]), .rdlo_out(a8_wr[424]));
			radix2 #(.width(width)) rd_st7_417  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[417]), .rdlo_in(a7_wr[425]),  .coef_in(coef[128]), .rdup_out(a8_wr[417]), .rdlo_out(a8_wr[425]));
			radix2 #(.width(width)) rd_st7_418  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[418]), .rdlo_in(a7_wr[426]),  .coef_in(coef[256]), .rdup_out(a8_wr[418]), .rdlo_out(a8_wr[426]));
			radix2 #(.width(width)) rd_st7_419  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[419]), .rdlo_in(a7_wr[427]),  .coef_in(coef[384]), .rdup_out(a8_wr[419]), .rdlo_out(a8_wr[427]));
			radix2 #(.width(width)) rd_st7_420  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[420]), .rdlo_in(a7_wr[428]),  .coef_in(coef[512]), .rdup_out(a8_wr[420]), .rdlo_out(a8_wr[428]));
			radix2 #(.width(width)) rd_st7_421  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[421]), .rdlo_in(a7_wr[429]),  .coef_in(coef[640]), .rdup_out(a8_wr[421]), .rdlo_out(a8_wr[429]));
			radix2 #(.width(width)) rd_st7_422  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[422]), .rdlo_in(a7_wr[430]),  .coef_in(coef[768]), .rdup_out(a8_wr[422]), .rdlo_out(a8_wr[430]));
			radix2 #(.width(width)) rd_st7_423  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[423]), .rdlo_in(a7_wr[431]),  .coef_in(coef[896]), .rdup_out(a8_wr[423]), .rdlo_out(a8_wr[431]));
			radix2 #(.width(width)) rd_st7_432  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[432]), .rdlo_in(a7_wr[440]),  .coef_in(coef[0]), .rdup_out(a8_wr[432]), .rdlo_out(a8_wr[440]));
			radix2 #(.width(width)) rd_st7_433  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[433]), .rdlo_in(a7_wr[441]),  .coef_in(coef[128]), .rdup_out(a8_wr[433]), .rdlo_out(a8_wr[441]));
			radix2 #(.width(width)) rd_st7_434  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[434]), .rdlo_in(a7_wr[442]),  .coef_in(coef[256]), .rdup_out(a8_wr[434]), .rdlo_out(a8_wr[442]));
			radix2 #(.width(width)) rd_st7_435  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[435]), .rdlo_in(a7_wr[443]),  .coef_in(coef[384]), .rdup_out(a8_wr[435]), .rdlo_out(a8_wr[443]));
			radix2 #(.width(width)) rd_st7_436  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[436]), .rdlo_in(a7_wr[444]),  .coef_in(coef[512]), .rdup_out(a8_wr[436]), .rdlo_out(a8_wr[444]));
			radix2 #(.width(width)) rd_st7_437  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[437]), .rdlo_in(a7_wr[445]),  .coef_in(coef[640]), .rdup_out(a8_wr[437]), .rdlo_out(a8_wr[445]));
			radix2 #(.width(width)) rd_st7_438  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[438]), .rdlo_in(a7_wr[446]),  .coef_in(coef[768]), .rdup_out(a8_wr[438]), .rdlo_out(a8_wr[446]));
			radix2 #(.width(width)) rd_st7_439  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[439]), .rdlo_in(a7_wr[447]),  .coef_in(coef[896]), .rdup_out(a8_wr[439]), .rdlo_out(a8_wr[447]));
			radix2 #(.width(width)) rd_st7_448  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[448]), .rdlo_in(a7_wr[456]),  .coef_in(coef[0]), .rdup_out(a8_wr[448]), .rdlo_out(a8_wr[456]));
			radix2 #(.width(width)) rd_st7_449  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[449]), .rdlo_in(a7_wr[457]),  .coef_in(coef[128]), .rdup_out(a8_wr[449]), .rdlo_out(a8_wr[457]));
			radix2 #(.width(width)) rd_st7_450  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[450]), .rdlo_in(a7_wr[458]),  .coef_in(coef[256]), .rdup_out(a8_wr[450]), .rdlo_out(a8_wr[458]));
			radix2 #(.width(width)) rd_st7_451  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[451]), .rdlo_in(a7_wr[459]),  .coef_in(coef[384]), .rdup_out(a8_wr[451]), .rdlo_out(a8_wr[459]));
			radix2 #(.width(width)) rd_st7_452  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[452]), .rdlo_in(a7_wr[460]),  .coef_in(coef[512]), .rdup_out(a8_wr[452]), .rdlo_out(a8_wr[460]));
			radix2 #(.width(width)) rd_st7_453  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[453]), .rdlo_in(a7_wr[461]),  .coef_in(coef[640]), .rdup_out(a8_wr[453]), .rdlo_out(a8_wr[461]));
			radix2 #(.width(width)) rd_st7_454  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[454]), .rdlo_in(a7_wr[462]),  .coef_in(coef[768]), .rdup_out(a8_wr[454]), .rdlo_out(a8_wr[462]));
			radix2 #(.width(width)) rd_st7_455  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[455]), .rdlo_in(a7_wr[463]),  .coef_in(coef[896]), .rdup_out(a8_wr[455]), .rdlo_out(a8_wr[463]));
			radix2 #(.width(width)) rd_st7_464  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[464]), .rdlo_in(a7_wr[472]),  .coef_in(coef[0]), .rdup_out(a8_wr[464]), .rdlo_out(a8_wr[472]));
			radix2 #(.width(width)) rd_st7_465  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[465]), .rdlo_in(a7_wr[473]),  .coef_in(coef[128]), .rdup_out(a8_wr[465]), .rdlo_out(a8_wr[473]));
			radix2 #(.width(width)) rd_st7_466  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[466]), .rdlo_in(a7_wr[474]),  .coef_in(coef[256]), .rdup_out(a8_wr[466]), .rdlo_out(a8_wr[474]));
			radix2 #(.width(width)) rd_st7_467  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[467]), .rdlo_in(a7_wr[475]),  .coef_in(coef[384]), .rdup_out(a8_wr[467]), .rdlo_out(a8_wr[475]));
			radix2 #(.width(width)) rd_st7_468  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[468]), .rdlo_in(a7_wr[476]),  .coef_in(coef[512]), .rdup_out(a8_wr[468]), .rdlo_out(a8_wr[476]));
			radix2 #(.width(width)) rd_st7_469  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[469]), .rdlo_in(a7_wr[477]),  .coef_in(coef[640]), .rdup_out(a8_wr[469]), .rdlo_out(a8_wr[477]));
			radix2 #(.width(width)) rd_st7_470  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[470]), .rdlo_in(a7_wr[478]),  .coef_in(coef[768]), .rdup_out(a8_wr[470]), .rdlo_out(a8_wr[478]));
			radix2 #(.width(width)) rd_st7_471  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[471]), .rdlo_in(a7_wr[479]),  .coef_in(coef[896]), .rdup_out(a8_wr[471]), .rdlo_out(a8_wr[479]));
			radix2 #(.width(width)) rd_st7_480  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[480]), .rdlo_in(a7_wr[488]),  .coef_in(coef[0]), .rdup_out(a8_wr[480]), .rdlo_out(a8_wr[488]));
			radix2 #(.width(width)) rd_st7_481  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[481]), .rdlo_in(a7_wr[489]),  .coef_in(coef[128]), .rdup_out(a8_wr[481]), .rdlo_out(a8_wr[489]));
			radix2 #(.width(width)) rd_st7_482  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[482]), .rdlo_in(a7_wr[490]),  .coef_in(coef[256]), .rdup_out(a8_wr[482]), .rdlo_out(a8_wr[490]));
			radix2 #(.width(width)) rd_st7_483  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[483]), .rdlo_in(a7_wr[491]),  .coef_in(coef[384]), .rdup_out(a8_wr[483]), .rdlo_out(a8_wr[491]));
			radix2 #(.width(width)) rd_st7_484  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[484]), .rdlo_in(a7_wr[492]),  .coef_in(coef[512]), .rdup_out(a8_wr[484]), .rdlo_out(a8_wr[492]));
			radix2 #(.width(width)) rd_st7_485  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[485]), .rdlo_in(a7_wr[493]),  .coef_in(coef[640]), .rdup_out(a8_wr[485]), .rdlo_out(a8_wr[493]));
			radix2 #(.width(width)) rd_st7_486  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[486]), .rdlo_in(a7_wr[494]),  .coef_in(coef[768]), .rdup_out(a8_wr[486]), .rdlo_out(a8_wr[494]));
			radix2 #(.width(width)) rd_st7_487  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[487]), .rdlo_in(a7_wr[495]),  .coef_in(coef[896]), .rdup_out(a8_wr[487]), .rdlo_out(a8_wr[495]));
			radix2 #(.width(width)) rd_st7_496  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[496]), .rdlo_in(a7_wr[504]),  .coef_in(coef[0]), .rdup_out(a8_wr[496]), .rdlo_out(a8_wr[504]));
			radix2 #(.width(width)) rd_st7_497  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[497]), .rdlo_in(a7_wr[505]),  .coef_in(coef[128]), .rdup_out(a8_wr[497]), .rdlo_out(a8_wr[505]));
			radix2 #(.width(width)) rd_st7_498  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[498]), .rdlo_in(a7_wr[506]),  .coef_in(coef[256]), .rdup_out(a8_wr[498]), .rdlo_out(a8_wr[506]));
			radix2 #(.width(width)) rd_st7_499  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[499]), .rdlo_in(a7_wr[507]),  .coef_in(coef[384]), .rdup_out(a8_wr[499]), .rdlo_out(a8_wr[507]));
			radix2 #(.width(width)) rd_st7_500  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[500]), .rdlo_in(a7_wr[508]),  .coef_in(coef[512]), .rdup_out(a8_wr[500]), .rdlo_out(a8_wr[508]));
			radix2 #(.width(width)) rd_st7_501  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[501]), .rdlo_in(a7_wr[509]),  .coef_in(coef[640]), .rdup_out(a8_wr[501]), .rdlo_out(a8_wr[509]));
			radix2 #(.width(width)) rd_st7_502  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[502]), .rdlo_in(a7_wr[510]),  .coef_in(coef[768]), .rdup_out(a8_wr[502]), .rdlo_out(a8_wr[510]));
			radix2 #(.width(width)) rd_st7_503  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[503]), .rdlo_in(a7_wr[511]),  .coef_in(coef[896]), .rdup_out(a8_wr[503]), .rdlo_out(a8_wr[511]));
			radix2 #(.width(width)) rd_st7_512  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[512]), .rdlo_in(a7_wr[520]),  .coef_in(coef[0]), .rdup_out(a8_wr[512]), .rdlo_out(a8_wr[520]));
			radix2 #(.width(width)) rd_st7_513  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[513]), .rdlo_in(a7_wr[521]),  .coef_in(coef[128]), .rdup_out(a8_wr[513]), .rdlo_out(a8_wr[521]));
			radix2 #(.width(width)) rd_st7_514  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[514]), .rdlo_in(a7_wr[522]),  .coef_in(coef[256]), .rdup_out(a8_wr[514]), .rdlo_out(a8_wr[522]));
			radix2 #(.width(width)) rd_st7_515  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[515]), .rdlo_in(a7_wr[523]),  .coef_in(coef[384]), .rdup_out(a8_wr[515]), .rdlo_out(a8_wr[523]));
			radix2 #(.width(width)) rd_st7_516  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[516]), .rdlo_in(a7_wr[524]),  .coef_in(coef[512]), .rdup_out(a8_wr[516]), .rdlo_out(a8_wr[524]));
			radix2 #(.width(width)) rd_st7_517  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[517]), .rdlo_in(a7_wr[525]),  .coef_in(coef[640]), .rdup_out(a8_wr[517]), .rdlo_out(a8_wr[525]));
			radix2 #(.width(width)) rd_st7_518  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[518]), .rdlo_in(a7_wr[526]),  .coef_in(coef[768]), .rdup_out(a8_wr[518]), .rdlo_out(a8_wr[526]));
			radix2 #(.width(width)) rd_st7_519  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[519]), .rdlo_in(a7_wr[527]),  .coef_in(coef[896]), .rdup_out(a8_wr[519]), .rdlo_out(a8_wr[527]));
			radix2 #(.width(width)) rd_st7_528  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[528]), .rdlo_in(a7_wr[536]),  .coef_in(coef[0]), .rdup_out(a8_wr[528]), .rdlo_out(a8_wr[536]));
			radix2 #(.width(width)) rd_st7_529  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[529]), .rdlo_in(a7_wr[537]),  .coef_in(coef[128]), .rdup_out(a8_wr[529]), .rdlo_out(a8_wr[537]));
			radix2 #(.width(width)) rd_st7_530  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[530]), .rdlo_in(a7_wr[538]),  .coef_in(coef[256]), .rdup_out(a8_wr[530]), .rdlo_out(a8_wr[538]));
			radix2 #(.width(width)) rd_st7_531  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[531]), .rdlo_in(a7_wr[539]),  .coef_in(coef[384]), .rdup_out(a8_wr[531]), .rdlo_out(a8_wr[539]));
			radix2 #(.width(width)) rd_st7_532  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[532]), .rdlo_in(a7_wr[540]),  .coef_in(coef[512]), .rdup_out(a8_wr[532]), .rdlo_out(a8_wr[540]));
			radix2 #(.width(width)) rd_st7_533  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[533]), .rdlo_in(a7_wr[541]),  .coef_in(coef[640]), .rdup_out(a8_wr[533]), .rdlo_out(a8_wr[541]));
			radix2 #(.width(width)) rd_st7_534  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[534]), .rdlo_in(a7_wr[542]),  .coef_in(coef[768]), .rdup_out(a8_wr[534]), .rdlo_out(a8_wr[542]));
			radix2 #(.width(width)) rd_st7_535  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[535]), .rdlo_in(a7_wr[543]),  .coef_in(coef[896]), .rdup_out(a8_wr[535]), .rdlo_out(a8_wr[543]));
			radix2 #(.width(width)) rd_st7_544  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[544]), .rdlo_in(a7_wr[552]),  .coef_in(coef[0]), .rdup_out(a8_wr[544]), .rdlo_out(a8_wr[552]));
			radix2 #(.width(width)) rd_st7_545  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[545]), .rdlo_in(a7_wr[553]),  .coef_in(coef[128]), .rdup_out(a8_wr[545]), .rdlo_out(a8_wr[553]));
			radix2 #(.width(width)) rd_st7_546  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[546]), .rdlo_in(a7_wr[554]),  .coef_in(coef[256]), .rdup_out(a8_wr[546]), .rdlo_out(a8_wr[554]));
			radix2 #(.width(width)) rd_st7_547  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[547]), .rdlo_in(a7_wr[555]),  .coef_in(coef[384]), .rdup_out(a8_wr[547]), .rdlo_out(a8_wr[555]));
			radix2 #(.width(width)) rd_st7_548  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[548]), .rdlo_in(a7_wr[556]),  .coef_in(coef[512]), .rdup_out(a8_wr[548]), .rdlo_out(a8_wr[556]));
			radix2 #(.width(width)) rd_st7_549  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[549]), .rdlo_in(a7_wr[557]),  .coef_in(coef[640]), .rdup_out(a8_wr[549]), .rdlo_out(a8_wr[557]));
			radix2 #(.width(width)) rd_st7_550  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[550]), .rdlo_in(a7_wr[558]),  .coef_in(coef[768]), .rdup_out(a8_wr[550]), .rdlo_out(a8_wr[558]));
			radix2 #(.width(width)) rd_st7_551  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[551]), .rdlo_in(a7_wr[559]),  .coef_in(coef[896]), .rdup_out(a8_wr[551]), .rdlo_out(a8_wr[559]));
			radix2 #(.width(width)) rd_st7_560  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[560]), .rdlo_in(a7_wr[568]),  .coef_in(coef[0]), .rdup_out(a8_wr[560]), .rdlo_out(a8_wr[568]));
			radix2 #(.width(width)) rd_st7_561  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[561]), .rdlo_in(a7_wr[569]),  .coef_in(coef[128]), .rdup_out(a8_wr[561]), .rdlo_out(a8_wr[569]));
			radix2 #(.width(width)) rd_st7_562  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[562]), .rdlo_in(a7_wr[570]),  .coef_in(coef[256]), .rdup_out(a8_wr[562]), .rdlo_out(a8_wr[570]));
			radix2 #(.width(width)) rd_st7_563  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[563]), .rdlo_in(a7_wr[571]),  .coef_in(coef[384]), .rdup_out(a8_wr[563]), .rdlo_out(a8_wr[571]));
			radix2 #(.width(width)) rd_st7_564  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[564]), .rdlo_in(a7_wr[572]),  .coef_in(coef[512]), .rdup_out(a8_wr[564]), .rdlo_out(a8_wr[572]));
			radix2 #(.width(width)) rd_st7_565  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[565]), .rdlo_in(a7_wr[573]),  .coef_in(coef[640]), .rdup_out(a8_wr[565]), .rdlo_out(a8_wr[573]));
			radix2 #(.width(width)) rd_st7_566  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[566]), .rdlo_in(a7_wr[574]),  .coef_in(coef[768]), .rdup_out(a8_wr[566]), .rdlo_out(a8_wr[574]));
			radix2 #(.width(width)) rd_st7_567  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[567]), .rdlo_in(a7_wr[575]),  .coef_in(coef[896]), .rdup_out(a8_wr[567]), .rdlo_out(a8_wr[575]));
			radix2 #(.width(width)) rd_st7_576  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[576]), .rdlo_in(a7_wr[584]),  .coef_in(coef[0]), .rdup_out(a8_wr[576]), .rdlo_out(a8_wr[584]));
			radix2 #(.width(width)) rd_st7_577  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[577]), .rdlo_in(a7_wr[585]),  .coef_in(coef[128]), .rdup_out(a8_wr[577]), .rdlo_out(a8_wr[585]));
			radix2 #(.width(width)) rd_st7_578  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[578]), .rdlo_in(a7_wr[586]),  .coef_in(coef[256]), .rdup_out(a8_wr[578]), .rdlo_out(a8_wr[586]));
			radix2 #(.width(width)) rd_st7_579  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[579]), .rdlo_in(a7_wr[587]),  .coef_in(coef[384]), .rdup_out(a8_wr[579]), .rdlo_out(a8_wr[587]));
			radix2 #(.width(width)) rd_st7_580  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[580]), .rdlo_in(a7_wr[588]),  .coef_in(coef[512]), .rdup_out(a8_wr[580]), .rdlo_out(a8_wr[588]));
			radix2 #(.width(width)) rd_st7_581  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[581]), .rdlo_in(a7_wr[589]),  .coef_in(coef[640]), .rdup_out(a8_wr[581]), .rdlo_out(a8_wr[589]));
			radix2 #(.width(width)) rd_st7_582  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[582]), .rdlo_in(a7_wr[590]),  .coef_in(coef[768]), .rdup_out(a8_wr[582]), .rdlo_out(a8_wr[590]));
			radix2 #(.width(width)) rd_st7_583  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[583]), .rdlo_in(a7_wr[591]),  .coef_in(coef[896]), .rdup_out(a8_wr[583]), .rdlo_out(a8_wr[591]));
			radix2 #(.width(width)) rd_st7_592  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[592]), .rdlo_in(a7_wr[600]),  .coef_in(coef[0]), .rdup_out(a8_wr[592]), .rdlo_out(a8_wr[600]));
			radix2 #(.width(width)) rd_st7_593  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[593]), .rdlo_in(a7_wr[601]),  .coef_in(coef[128]), .rdup_out(a8_wr[593]), .rdlo_out(a8_wr[601]));
			radix2 #(.width(width)) rd_st7_594  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[594]), .rdlo_in(a7_wr[602]),  .coef_in(coef[256]), .rdup_out(a8_wr[594]), .rdlo_out(a8_wr[602]));
			radix2 #(.width(width)) rd_st7_595  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[595]), .rdlo_in(a7_wr[603]),  .coef_in(coef[384]), .rdup_out(a8_wr[595]), .rdlo_out(a8_wr[603]));
			radix2 #(.width(width)) rd_st7_596  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[596]), .rdlo_in(a7_wr[604]),  .coef_in(coef[512]), .rdup_out(a8_wr[596]), .rdlo_out(a8_wr[604]));
			radix2 #(.width(width)) rd_st7_597  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[597]), .rdlo_in(a7_wr[605]),  .coef_in(coef[640]), .rdup_out(a8_wr[597]), .rdlo_out(a8_wr[605]));
			radix2 #(.width(width)) rd_st7_598  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[598]), .rdlo_in(a7_wr[606]),  .coef_in(coef[768]), .rdup_out(a8_wr[598]), .rdlo_out(a8_wr[606]));
			radix2 #(.width(width)) rd_st7_599  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[599]), .rdlo_in(a7_wr[607]),  .coef_in(coef[896]), .rdup_out(a8_wr[599]), .rdlo_out(a8_wr[607]));
			radix2 #(.width(width)) rd_st7_608  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[608]), .rdlo_in(a7_wr[616]),  .coef_in(coef[0]), .rdup_out(a8_wr[608]), .rdlo_out(a8_wr[616]));
			radix2 #(.width(width)) rd_st7_609  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[609]), .rdlo_in(a7_wr[617]),  .coef_in(coef[128]), .rdup_out(a8_wr[609]), .rdlo_out(a8_wr[617]));
			radix2 #(.width(width)) rd_st7_610  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[610]), .rdlo_in(a7_wr[618]),  .coef_in(coef[256]), .rdup_out(a8_wr[610]), .rdlo_out(a8_wr[618]));
			radix2 #(.width(width)) rd_st7_611  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[611]), .rdlo_in(a7_wr[619]),  .coef_in(coef[384]), .rdup_out(a8_wr[611]), .rdlo_out(a8_wr[619]));
			radix2 #(.width(width)) rd_st7_612  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[612]), .rdlo_in(a7_wr[620]),  .coef_in(coef[512]), .rdup_out(a8_wr[612]), .rdlo_out(a8_wr[620]));
			radix2 #(.width(width)) rd_st7_613  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[613]), .rdlo_in(a7_wr[621]),  .coef_in(coef[640]), .rdup_out(a8_wr[613]), .rdlo_out(a8_wr[621]));
			radix2 #(.width(width)) rd_st7_614  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[614]), .rdlo_in(a7_wr[622]),  .coef_in(coef[768]), .rdup_out(a8_wr[614]), .rdlo_out(a8_wr[622]));
			radix2 #(.width(width)) rd_st7_615  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[615]), .rdlo_in(a7_wr[623]),  .coef_in(coef[896]), .rdup_out(a8_wr[615]), .rdlo_out(a8_wr[623]));
			radix2 #(.width(width)) rd_st7_624  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[624]), .rdlo_in(a7_wr[632]),  .coef_in(coef[0]), .rdup_out(a8_wr[624]), .rdlo_out(a8_wr[632]));
			radix2 #(.width(width)) rd_st7_625  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[625]), .rdlo_in(a7_wr[633]),  .coef_in(coef[128]), .rdup_out(a8_wr[625]), .rdlo_out(a8_wr[633]));
			radix2 #(.width(width)) rd_st7_626  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[626]), .rdlo_in(a7_wr[634]),  .coef_in(coef[256]), .rdup_out(a8_wr[626]), .rdlo_out(a8_wr[634]));
			radix2 #(.width(width)) rd_st7_627  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[627]), .rdlo_in(a7_wr[635]),  .coef_in(coef[384]), .rdup_out(a8_wr[627]), .rdlo_out(a8_wr[635]));
			radix2 #(.width(width)) rd_st7_628  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[628]), .rdlo_in(a7_wr[636]),  .coef_in(coef[512]), .rdup_out(a8_wr[628]), .rdlo_out(a8_wr[636]));
			radix2 #(.width(width)) rd_st7_629  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[629]), .rdlo_in(a7_wr[637]),  .coef_in(coef[640]), .rdup_out(a8_wr[629]), .rdlo_out(a8_wr[637]));
			radix2 #(.width(width)) rd_st7_630  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[630]), .rdlo_in(a7_wr[638]),  .coef_in(coef[768]), .rdup_out(a8_wr[630]), .rdlo_out(a8_wr[638]));
			radix2 #(.width(width)) rd_st7_631  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[631]), .rdlo_in(a7_wr[639]),  .coef_in(coef[896]), .rdup_out(a8_wr[631]), .rdlo_out(a8_wr[639]));
			radix2 #(.width(width)) rd_st7_640  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[640]), .rdlo_in(a7_wr[648]),  .coef_in(coef[0]), .rdup_out(a8_wr[640]), .rdlo_out(a8_wr[648]));
			radix2 #(.width(width)) rd_st7_641  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[641]), .rdlo_in(a7_wr[649]),  .coef_in(coef[128]), .rdup_out(a8_wr[641]), .rdlo_out(a8_wr[649]));
			radix2 #(.width(width)) rd_st7_642  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[642]), .rdlo_in(a7_wr[650]),  .coef_in(coef[256]), .rdup_out(a8_wr[642]), .rdlo_out(a8_wr[650]));
			radix2 #(.width(width)) rd_st7_643  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[643]), .rdlo_in(a7_wr[651]),  .coef_in(coef[384]), .rdup_out(a8_wr[643]), .rdlo_out(a8_wr[651]));
			radix2 #(.width(width)) rd_st7_644  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[644]), .rdlo_in(a7_wr[652]),  .coef_in(coef[512]), .rdup_out(a8_wr[644]), .rdlo_out(a8_wr[652]));
			radix2 #(.width(width)) rd_st7_645  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[645]), .rdlo_in(a7_wr[653]),  .coef_in(coef[640]), .rdup_out(a8_wr[645]), .rdlo_out(a8_wr[653]));
			radix2 #(.width(width)) rd_st7_646  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[646]), .rdlo_in(a7_wr[654]),  .coef_in(coef[768]), .rdup_out(a8_wr[646]), .rdlo_out(a8_wr[654]));
			radix2 #(.width(width)) rd_st7_647  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[647]), .rdlo_in(a7_wr[655]),  .coef_in(coef[896]), .rdup_out(a8_wr[647]), .rdlo_out(a8_wr[655]));
			radix2 #(.width(width)) rd_st7_656  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[656]), .rdlo_in(a7_wr[664]),  .coef_in(coef[0]), .rdup_out(a8_wr[656]), .rdlo_out(a8_wr[664]));
			radix2 #(.width(width)) rd_st7_657  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[657]), .rdlo_in(a7_wr[665]),  .coef_in(coef[128]), .rdup_out(a8_wr[657]), .rdlo_out(a8_wr[665]));
			radix2 #(.width(width)) rd_st7_658  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[658]), .rdlo_in(a7_wr[666]),  .coef_in(coef[256]), .rdup_out(a8_wr[658]), .rdlo_out(a8_wr[666]));
			radix2 #(.width(width)) rd_st7_659  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[659]), .rdlo_in(a7_wr[667]),  .coef_in(coef[384]), .rdup_out(a8_wr[659]), .rdlo_out(a8_wr[667]));
			radix2 #(.width(width)) rd_st7_660  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[660]), .rdlo_in(a7_wr[668]),  .coef_in(coef[512]), .rdup_out(a8_wr[660]), .rdlo_out(a8_wr[668]));
			radix2 #(.width(width)) rd_st7_661  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[661]), .rdlo_in(a7_wr[669]),  .coef_in(coef[640]), .rdup_out(a8_wr[661]), .rdlo_out(a8_wr[669]));
			radix2 #(.width(width)) rd_st7_662  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[662]), .rdlo_in(a7_wr[670]),  .coef_in(coef[768]), .rdup_out(a8_wr[662]), .rdlo_out(a8_wr[670]));
			radix2 #(.width(width)) rd_st7_663  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[663]), .rdlo_in(a7_wr[671]),  .coef_in(coef[896]), .rdup_out(a8_wr[663]), .rdlo_out(a8_wr[671]));
			radix2 #(.width(width)) rd_st7_672  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[672]), .rdlo_in(a7_wr[680]),  .coef_in(coef[0]), .rdup_out(a8_wr[672]), .rdlo_out(a8_wr[680]));
			radix2 #(.width(width)) rd_st7_673  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[673]), .rdlo_in(a7_wr[681]),  .coef_in(coef[128]), .rdup_out(a8_wr[673]), .rdlo_out(a8_wr[681]));
			radix2 #(.width(width)) rd_st7_674  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[674]), .rdlo_in(a7_wr[682]),  .coef_in(coef[256]), .rdup_out(a8_wr[674]), .rdlo_out(a8_wr[682]));
			radix2 #(.width(width)) rd_st7_675  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[675]), .rdlo_in(a7_wr[683]),  .coef_in(coef[384]), .rdup_out(a8_wr[675]), .rdlo_out(a8_wr[683]));
			radix2 #(.width(width)) rd_st7_676  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[676]), .rdlo_in(a7_wr[684]),  .coef_in(coef[512]), .rdup_out(a8_wr[676]), .rdlo_out(a8_wr[684]));
			radix2 #(.width(width)) rd_st7_677  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[677]), .rdlo_in(a7_wr[685]),  .coef_in(coef[640]), .rdup_out(a8_wr[677]), .rdlo_out(a8_wr[685]));
			radix2 #(.width(width)) rd_st7_678  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[678]), .rdlo_in(a7_wr[686]),  .coef_in(coef[768]), .rdup_out(a8_wr[678]), .rdlo_out(a8_wr[686]));
			radix2 #(.width(width)) rd_st7_679  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[679]), .rdlo_in(a7_wr[687]),  .coef_in(coef[896]), .rdup_out(a8_wr[679]), .rdlo_out(a8_wr[687]));
			radix2 #(.width(width)) rd_st7_688  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[688]), .rdlo_in(a7_wr[696]),  .coef_in(coef[0]), .rdup_out(a8_wr[688]), .rdlo_out(a8_wr[696]));
			radix2 #(.width(width)) rd_st7_689  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[689]), .rdlo_in(a7_wr[697]),  .coef_in(coef[128]), .rdup_out(a8_wr[689]), .rdlo_out(a8_wr[697]));
			radix2 #(.width(width)) rd_st7_690  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[690]), .rdlo_in(a7_wr[698]),  .coef_in(coef[256]), .rdup_out(a8_wr[690]), .rdlo_out(a8_wr[698]));
			radix2 #(.width(width)) rd_st7_691  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[691]), .rdlo_in(a7_wr[699]),  .coef_in(coef[384]), .rdup_out(a8_wr[691]), .rdlo_out(a8_wr[699]));
			radix2 #(.width(width)) rd_st7_692  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[692]), .rdlo_in(a7_wr[700]),  .coef_in(coef[512]), .rdup_out(a8_wr[692]), .rdlo_out(a8_wr[700]));
			radix2 #(.width(width)) rd_st7_693  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[693]), .rdlo_in(a7_wr[701]),  .coef_in(coef[640]), .rdup_out(a8_wr[693]), .rdlo_out(a8_wr[701]));
			radix2 #(.width(width)) rd_st7_694  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[694]), .rdlo_in(a7_wr[702]),  .coef_in(coef[768]), .rdup_out(a8_wr[694]), .rdlo_out(a8_wr[702]));
			radix2 #(.width(width)) rd_st7_695  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[695]), .rdlo_in(a7_wr[703]),  .coef_in(coef[896]), .rdup_out(a8_wr[695]), .rdlo_out(a8_wr[703]));
			radix2 #(.width(width)) rd_st7_704  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[704]), .rdlo_in(a7_wr[712]),  .coef_in(coef[0]), .rdup_out(a8_wr[704]), .rdlo_out(a8_wr[712]));
			radix2 #(.width(width)) rd_st7_705  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[705]), .rdlo_in(a7_wr[713]),  .coef_in(coef[128]), .rdup_out(a8_wr[705]), .rdlo_out(a8_wr[713]));
			radix2 #(.width(width)) rd_st7_706  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[706]), .rdlo_in(a7_wr[714]),  .coef_in(coef[256]), .rdup_out(a8_wr[706]), .rdlo_out(a8_wr[714]));
			radix2 #(.width(width)) rd_st7_707  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[707]), .rdlo_in(a7_wr[715]),  .coef_in(coef[384]), .rdup_out(a8_wr[707]), .rdlo_out(a8_wr[715]));
			radix2 #(.width(width)) rd_st7_708  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[708]), .rdlo_in(a7_wr[716]),  .coef_in(coef[512]), .rdup_out(a8_wr[708]), .rdlo_out(a8_wr[716]));
			radix2 #(.width(width)) rd_st7_709  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[709]), .rdlo_in(a7_wr[717]),  .coef_in(coef[640]), .rdup_out(a8_wr[709]), .rdlo_out(a8_wr[717]));
			radix2 #(.width(width)) rd_st7_710  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[710]), .rdlo_in(a7_wr[718]),  .coef_in(coef[768]), .rdup_out(a8_wr[710]), .rdlo_out(a8_wr[718]));
			radix2 #(.width(width)) rd_st7_711  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[711]), .rdlo_in(a7_wr[719]),  .coef_in(coef[896]), .rdup_out(a8_wr[711]), .rdlo_out(a8_wr[719]));
			radix2 #(.width(width)) rd_st7_720  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[720]), .rdlo_in(a7_wr[728]),  .coef_in(coef[0]), .rdup_out(a8_wr[720]), .rdlo_out(a8_wr[728]));
			radix2 #(.width(width)) rd_st7_721  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[721]), .rdlo_in(a7_wr[729]),  .coef_in(coef[128]), .rdup_out(a8_wr[721]), .rdlo_out(a8_wr[729]));
			radix2 #(.width(width)) rd_st7_722  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[722]), .rdlo_in(a7_wr[730]),  .coef_in(coef[256]), .rdup_out(a8_wr[722]), .rdlo_out(a8_wr[730]));
			radix2 #(.width(width)) rd_st7_723  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[723]), .rdlo_in(a7_wr[731]),  .coef_in(coef[384]), .rdup_out(a8_wr[723]), .rdlo_out(a8_wr[731]));
			radix2 #(.width(width)) rd_st7_724  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[724]), .rdlo_in(a7_wr[732]),  .coef_in(coef[512]), .rdup_out(a8_wr[724]), .rdlo_out(a8_wr[732]));
			radix2 #(.width(width)) rd_st7_725  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[725]), .rdlo_in(a7_wr[733]),  .coef_in(coef[640]), .rdup_out(a8_wr[725]), .rdlo_out(a8_wr[733]));
			radix2 #(.width(width)) rd_st7_726  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[726]), .rdlo_in(a7_wr[734]),  .coef_in(coef[768]), .rdup_out(a8_wr[726]), .rdlo_out(a8_wr[734]));
			radix2 #(.width(width)) rd_st7_727  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[727]), .rdlo_in(a7_wr[735]),  .coef_in(coef[896]), .rdup_out(a8_wr[727]), .rdlo_out(a8_wr[735]));
			radix2 #(.width(width)) rd_st7_736  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[736]), .rdlo_in(a7_wr[744]),  .coef_in(coef[0]), .rdup_out(a8_wr[736]), .rdlo_out(a8_wr[744]));
			radix2 #(.width(width)) rd_st7_737  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[737]), .rdlo_in(a7_wr[745]),  .coef_in(coef[128]), .rdup_out(a8_wr[737]), .rdlo_out(a8_wr[745]));
			radix2 #(.width(width)) rd_st7_738  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[738]), .rdlo_in(a7_wr[746]),  .coef_in(coef[256]), .rdup_out(a8_wr[738]), .rdlo_out(a8_wr[746]));
			radix2 #(.width(width)) rd_st7_739  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[739]), .rdlo_in(a7_wr[747]),  .coef_in(coef[384]), .rdup_out(a8_wr[739]), .rdlo_out(a8_wr[747]));
			radix2 #(.width(width)) rd_st7_740  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[740]), .rdlo_in(a7_wr[748]),  .coef_in(coef[512]), .rdup_out(a8_wr[740]), .rdlo_out(a8_wr[748]));
			radix2 #(.width(width)) rd_st7_741  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[741]), .rdlo_in(a7_wr[749]),  .coef_in(coef[640]), .rdup_out(a8_wr[741]), .rdlo_out(a8_wr[749]));
			radix2 #(.width(width)) rd_st7_742  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[742]), .rdlo_in(a7_wr[750]),  .coef_in(coef[768]), .rdup_out(a8_wr[742]), .rdlo_out(a8_wr[750]));
			radix2 #(.width(width)) rd_st7_743  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[743]), .rdlo_in(a7_wr[751]),  .coef_in(coef[896]), .rdup_out(a8_wr[743]), .rdlo_out(a8_wr[751]));
			radix2 #(.width(width)) rd_st7_752  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[752]), .rdlo_in(a7_wr[760]),  .coef_in(coef[0]), .rdup_out(a8_wr[752]), .rdlo_out(a8_wr[760]));
			radix2 #(.width(width)) rd_st7_753  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[753]), .rdlo_in(a7_wr[761]),  .coef_in(coef[128]), .rdup_out(a8_wr[753]), .rdlo_out(a8_wr[761]));
			radix2 #(.width(width)) rd_st7_754  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[754]), .rdlo_in(a7_wr[762]),  .coef_in(coef[256]), .rdup_out(a8_wr[754]), .rdlo_out(a8_wr[762]));
			radix2 #(.width(width)) rd_st7_755  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[755]), .rdlo_in(a7_wr[763]),  .coef_in(coef[384]), .rdup_out(a8_wr[755]), .rdlo_out(a8_wr[763]));
			radix2 #(.width(width)) rd_st7_756  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[756]), .rdlo_in(a7_wr[764]),  .coef_in(coef[512]), .rdup_out(a8_wr[756]), .rdlo_out(a8_wr[764]));
			radix2 #(.width(width)) rd_st7_757  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[757]), .rdlo_in(a7_wr[765]),  .coef_in(coef[640]), .rdup_out(a8_wr[757]), .rdlo_out(a8_wr[765]));
			radix2 #(.width(width)) rd_st7_758  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[758]), .rdlo_in(a7_wr[766]),  .coef_in(coef[768]), .rdup_out(a8_wr[758]), .rdlo_out(a8_wr[766]));
			radix2 #(.width(width)) rd_st7_759  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[759]), .rdlo_in(a7_wr[767]),  .coef_in(coef[896]), .rdup_out(a8_wr[759]), .rdlo_out(a8_wr[767]));
			radix2 #(.width(width)) rd_st7_768  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[768]), .rdlo_in(a7_wr[776]),  .coef_in(coef[0]), .rdup_out(a8_wr[768]), .rdlo_out(a8_wr[776]));
			radix2 #(.width(width)) rd_st7_769  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[769]), .rdlo_in(a7_wr[777]),  .coef_in(coef[128]), .rdup_out(a8_wr[769]), .rdlo_out(a8_wr[777]));
			radix2 #(.width(width)) rd_st7_770  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[770]), .rdlo_in(a7_wr[778]),  .coef_in(coef[256]), .rdup_out(a8_wr[770]), .rdlo_out(a8_wr[778]));
			radix2 #(.width(width)) rd_st7_771  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[771]), .rdlo_in(a7_wr[779]),  .coef_in(coef[384]), .rdup_out(a8_wr[771]), .rdlo_out(a8_wr[779]));
			radix2 #(.width(width)) rd_st7_772  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[772]), .rdlo_in(a7_wr[780]),  .coef_in(coef[512]), .rdup_out(a8_wr[772]), .rdlo_out(a8_wr[780]));
			radix2 #(.width(width)) rd_st7_773  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[773]), .rdlo_in(a7_wr[781]),  .coef_in(coef[640]), .rdup_out(a8_wr[773]), .rdlo_out(a8_wr[781]));
			radix2 #(.width(width)) rd_st7_774  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[774]), .rdlo_in(a7_wr[782]),  .coef_in(coef[768]), .rdup_out(a8_wr[774]), .rdlo_out(a8_wr[782]));
			radix2 #(.width(width)) rd_st7_775  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[775]), .rdlo_in(a7_wr[783]),  .coef_in(coef[896]), .rdup_out(a8_wr[775]), .rdlo_out(a8_wr[783]));
			radix2 #(.width(width)) rd_st7_784  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[784]), .rdlo_in(a7_wr[792]),  .coef_in(coef[0]), .rdup_out(a8_wr[784]), .rdlo_out(a8_wr[792]));
			radix2 #(.width(width)) rd_st7_785  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[785]), .rdlo_in(a7_wr[793]),  .coef_in(coef[128]), .rdup_out(a8_wr[785]), .rdlo_out(a8_wr[793]));
			radix2 #(.width(width)) rd_st7_786  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[786]), .rdlo_in(a7_wr[794]),  .coef_in(coef[256]), .rdup_out(a8_wr[786]), .rdlo_out(a8_wr[794]));
			radix2 #(.width(width)) rd_st7_787  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[787]), .rdlo_in(a7_wr[795]),  .coef_in(coef[384]), .rdup_out(a8_wr[787]), .rdlo_out(a8_wr[795]));
			radix2 #(.width(width)) rd_st7_788  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[788]), .rdlo_in(a7_wr[796]),  .coef_in(coef[512]), .rdup_out(a8_wr[788]), .rdlo_out(a8_wr[796]));
			radix2 #(.width(width)) rd_st7_789  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[789]), .rdlo_in(a7_wr[797]),  .coef_in(coef[640]), .rdup_out(a8_wr[789]), .rdlo_out(a8_wr[797]));
			radix2 #(.width(width)) rd_st7_790  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[790]), .rdlo_in(a7_wr[798]),  .coef_in(coef[768]), .rdup_out(a8_wr[790]), .rdlo_out(a8_wr[798]));
			radix2 #(.width(width)) rd_st7_791  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[791]), .rdlo_in(a7_wr[799]),  .coef_in(coef[896]), .rdup_out(a8_wr[791]), .rdlo_out(a8_wr[799]));
			radix2 #(.width(width)) rd_st7_800  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[800]), .rdlo_in(a7_wr[808]),  .coef_in(coef[0]), .rdup_out(a8_wr[800]), .rdlo_out(a8_wr[808]));
			radix2 #(.width(width)) rd_st7_801  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[801]), .rdlo_in(a7_wr[809]),  .coef_in(coef[128]), .rdup_out(a8_wr[801]), .rdlo_out(a8_wr[809]));
			radix2 #(.width(width)) rd_st7_802  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[802]), .rdlo_in(a7_wr[810]),  .coef_in(coef[256]), .rdup_out(a8_wr[802]), .rdlo_out(a8_wr[810]));
			radix2 #(.width(width)) rd_st7_803  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[803]), .rdlo_in(a7_wr[811]),  .coef_in(coef[384]), .rdup_out(a8_wr[803]), .rdlo_out(a8_wr[811]));
			radix2 #(.width(width)) rd_st7_804  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[804]), .rdlo_in(a7_wr[812]),  .coef_in(coef[512]), .rdup_out(a8_wr[804]), .rdlo_out(a8_wr[812]));
			radix2 #(.width(width)) rd_st7_805  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[805]), .rdlo_in(a7_wr[813]),  .coef_in(coef[640]), .rdup_out(a8_wr[805]), .rdlo_out(a8_wr[813]));
			radix2 #(.width(width)) rd_st7_806  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[806]), .rdlo_in(a7_wr[814]),  .coef_in(coef[768]), .rdup_out(a8_wr[806]), .rdlo_out(a8_wr[814]));
			radix2 #(.width(width)) rd_st7_807  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[807]), .rdlo_in(a7_wr[815]),  .coef_in(coef[896]), .rdup_out(a8_wr[807]), .rdlo_out(a8_wr[815]));
			radix2 #(.width(width)) rd_st7_816  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[816]), .rdlo_in(a7_wr[824]),  .coef_in(coef[0]), .rdup_out(a8_wr[816]), .rdlo_out(a8_wr[824]));
			radix2 #(.width(width)) rd_st7_817  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[817]), .rdlo_in(a7_wr[825]),  .coef_in(coef[128]), .rdup_out(a8_wr[817]), .rdlo_out(a8_wr[825]));
			radix2 #(.width(width)) rd_st7_818  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[818]), .rdlo_in(a7_wr[826]),  .coef_in(coef[256]), .rdup_out(a8_wr[818]), .rdlo_out(a8_wr[826]));
			radix2 #(.width(width)) rd_st7_819  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[819]), .rdlo_in(a7_wr[827]),  .coef_in(coef[384]), .rdup_out(a8_wr[819]), .rdlo_out(a8_wr[827]));
			radix2 #(.width(width)) rd_st7_820  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[820]), .rdlo_in(a7_wr[828]),  .coef_in(coef[512]), .rdup_out(a8_wr[820]), .rdlo_out(a8_wr[828]));
			radix2 #(.width(width)) rd_st7_821  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[821]), .rdlo_in(a7_wr[829]),  .coef_in(coef[640]), .rdup_out(a8_wr[821]), .rdlo_out(a8_wr[829]));
			radix2 #(.width(width)) rd_st7_822  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[822]), .rdlo_in(a7_wr[830]),  .coef_in(coef[768]), .rdup_out(a8_wr[822]), .rdlo_out(a8_wr[830]));
			radix2 #(.width(width)) rd_st7_823  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[823]), .rdlo_in(a7_wr[831]),  .coef_in(coef[896]), .rdup_out(a8_wr[823]), .rdlo_out(a8_wr[831]));
			radix2 #(.width(width)) rd_st7_832  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[832]), .rdlo_in(a7_wr[840]),  .coef_in(coef[0]), .rdup_out(a8_wr[832]), .rdlo_out(a8_wr[840]));
			radix2 #(.width(width)) rd_st7_833  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[833]), .rdlo_in(a7_wr[841]),  .coef_in(coef[128]), .rdup_out(a8_wr[833]), .rdlo_out(a8_wr[841]));
			radix2 #(.width(width)) rd_st7_834  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[834]), .rdlo_in(a7_wr[842]),  .coef_in(coef[256]), .rdup_out(a8_wr[834]), .rdlo_out(a8_wr[842]));
			radix2 #(.width(width)) rd_st7_835  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[835]), .rdlo_in(a7_wr[843]),  .coef_in(coef[384]), .rdup_out(a8_wr[835]), .rdlo_out(a8_wr[843]));
			radix2 #(.width(width)) rd_st7_836  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[836]), .rdlo_in(a7_wr[844]),  .coef_in(coef[512]), .rdup_out(a8_wr[836]), .rdlo_out(a8_wr[844]));
			radix2 #(.width(width)) rd_st7_837  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[837]), .rdlo_in(a7_wr[845]),  .coef_in(coef[640]), .rdup_out(a8_wr[837]), .rdlo_out(a8_wr[845]));
			radix2 #(.width(width)) rd_st7_838  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[838]), .rdlo_in(a7_wr[846]),  .coef_in(coef[768]), .rdup_out(a8_wr[838]), .rdlo_out(a8_wr[846]));
			radix2 #(.width(width)) rd_st7_839  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[839]), .rdlo_in(a7_wr[847]),  .coef_in(coef[896]), .rdup_out(a8_wr[839]), .rdlo_out(a8_wr[847]));
			radix2 #(.width(width)) rd_st7_848  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[848]), .rdlo_in(a7_wr[856]),  .coef_in(coef[0]), .rdup_out(a8_wr[848]), .rdlo_out(a8_wr[856]));
			radix2 #(.width(width)) rd_st7_849  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[849]), .rdlo_in(a7_wr[857]),  .coef_in(coef[128]), .rdup_out(a8_wr[849]), .rdlo_out(a8_wr[857]));
			radix2 #(.width(width)) rd_st7_850  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[850]), .rdlo_in(a7_wr[858]),  .coef_in(coef[256]), .rdup_out(a8_wr[850]), .rdlo_out(a8_wr[858]));
			radix2 #(.width(width)) rd_st7_851  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[851]), .rdlo_in(a7_wr[859]),  .coef_in(coef[384]), .rdup_out(a8_wr[851]), .rdlo_out(a8_wr[859]));
			radix2 #(.width(width)) rd_st7_852  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[852]), .rdlo_in(a7_wr[860]),  .coef_in(coef[512]), .rdup_out(a8_wr[852]), .rdlo_out(a8_wr[860]));
			radix2 #(.width(width)) rd_st7_853  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[853]), .rdlo_in(a7_wr[861]),  .coef_in(coef[640]), .rdup_out(a8_wr[853]), .rdlo_out(a8_wr[861]));
			radix2 #(.width(width)) rd_st7_854  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[854]), .rdlo_in(a7_wr[862]),  .coef_in(coef[768]), .rdup_out(a8_wr[854]), .rdlo_out(a8_wr[862]));
			radix2 #(.width(width)) rd_st7_855  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[855]), .rdlo_in(a7_wr[863]),  .coef_in(coef[896]), .rdup_out(a8_wr[855]), .rdlo_out(a8_wr[863]));
			radix2 #(.width(width)) rd_st7_864  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[864]), .rdlo_in(a7_wr[872]),  .coef_in(coef[0]), .rdup_out(a8_wr[864]), .rdlo_out(a8_wr[872]));
			radix2 #(.width(width)) rd_st7_865  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[865]), .rdlo_in(a7_wr[873]),  .coef_in(coef[128]), .rdup_out(a8_wr[865]), .rdlo_out(a8_wr[873]));
			radix2 #(.width(width)) rd_st7_866  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[866]), .rdlo_in(a7_wr[874]),  .coef_in(coef[256]), .rdup_out(a8_wr[866]), .rdlo_out(a8_wr[874]));
			radix2 #(.width(width)) rd_st7_867  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[867]), .rdlo_in(a7_wr[875]),  .coef_in(coef[384]), .rdup_out(a8_wr[867]), .rdlo_out(a8_wr[875]));
			radix2 #(.width(width)) rd_st7_868  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[868]), .rdlo_in(a7_wr[876]),  .coef_in(coef[512]), .rdup_out(a8_wr[868]), .rdlo_out(a8_wr[876]));
			radix2 #(.width(width)) rd_st7_869  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[869]), .rdlo_in(a7_wr[877]),  .coef_in(coef[640]), .rdup_out(a8_wr[869]), .rdlo_out(a8_wr[877]));
			radix2 #(.width(width)) rd_st7_870  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[870]), .rdlo_in(a7_wr[878]),  .coef_in(coef[768]), .rdup_out(a8_wr[870]), .rdlo_out(a8_wr[878]));
			radix2 #(.width(width)) rd_st7_871  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[871]), .rdlo_in(a7_wr[879]),  .coef_in(coef[896]), .rdup_out(a8_wr[871]), .rdlo_out(a8_wr[879]));
			radix2 #(.width(width)) rd_st7_880  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[880]), .rdlo_in(a7_wr[888]),  .coef_in(coef[0]), .rdup_out(a8_wr[880]), .rdlo_out(a8_wr[888]));
			radix2 #(.width(width)) rd_st7_881  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[881]), .rdlo_in(a7_wr[889]),  .coef_in(coef[128]), .rdup_out(a8_wr[881]), .rdlo_out(a8_wr[889]));
			radix2 #(.width(width)) rd_st7_882  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[882]), .rdlo_in(a7_wr[890]),  .coef_in(coef[256]), .rdup_out(a8_wr[882]), .rdlo_out(a8_wr[890]));
			radix2 #(.width(width)) rd_st7_883  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[883]), .rdlo_in(a7_wr[891]),  .coef_in(coef[384]), .rdup_out(a8_wr[883]), .rdlo_out(a8_wr[891]));
			radix2 #(.width(width)) rd_st7_884  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[884]), .rdlo_in(a7_wr[892]),  .coef_in(coef[512]), .rdup_out(a8_wr[884]), .rdlo_out(a8_wr[892]));
			radix2 #(.width(width)) rd_st7_885  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[885]), .rdlo_in(a7_wr[893]),  .coef_in(coef[640]), .rdup_out(a8_wr[885]), .rdlo_out(a8_wr[893]));
			radix2 #(.width(width)) rd_st7_886  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[886]), .rdlo_in(a7_wr[894]),  .coef_in(coef[768]), .rdup_out(a8_wr[886]), .rdlo_out(a8_wr[894]));
			radix2 #(.width(width)) rd_st7_887  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[887]), .rdlo_in(a7_wr[895]),  .coef_in(coef[896]), .rdup_out(a8_wr[887]), .rdlo_out(a8_wr[895]));
			radix2 #(.width(width)) rd_st7_896  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[896]), .rdlo_in(a7_wr[904]),  .coef_in(coef[0]), .rdup_out(a8_wr[896]), .rdlo_out(a8_wr[904]));
			radix2 #(.width(width)) rd_st7_897  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[897]), .rdlo_in(a7_wr[905]),  .coef_in(coef[128]), .rdup_out(a8_wr[897]), .rdlo_out(a8_wr[905]));
			radix2 #(.width(width)) rd_st7_898  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[898]), .rdlo_in(a7_wr[906]),  .coef_in(coef[256]), .rdup_out(a8_wr[898]), .rdlo_out(a8_wr[906]));
			radix2 #(.width(width)) rd_st7_899  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[899]), .rdlo_in(a7_wr[907]),  .coef_in(coef[384]), .rdup_out(a8_wr[899]), .rdlo_out(a8_wr[907]));
			radix2 #(.width(width)) rd_st7_900  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[900]), .rdlo_in(a7_wr[908]),  .coef_in(coef[512]), .rdup_out(a8_wr[900]), .rdlo_out(a8_wr[908]));
			radix2 #(.width(width)) rd_st7_901  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[901]), .rdlo_in(a7_wr[909]),  .coef_in(coef[640]), .rdup_out(a8_wr[901]), .rdlo_out(a8_wr[909]));
			radix2 #(.width(width)) rd_st7_902  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[902]), .rdlo_in(a7_wr[910]),  .coef_in(coef[768]), .rdup_out(a8_wr[902]), .rdlo_out(a8_wr[910]));
			radix2 #(.width(width)) rd_st7_903  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[903]), .rdlo_in(a7_wr[911]),  .coef_in(coef[896]), .rdup_out(a8_wr[903]), .rdlo_out(a8_wr[911]));
			radix2 #(.width(width)) rd_st7_912  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[912]), .rdlo_in(a7_wr[920]),  .coef_in(coef[0]), .rdup_out(a8_wr[912]), .rdlo_out(a8_wr[920]));
			radix2 #(.width(width)) rd_st7_913  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[913]), .rdlo_in(a7_wr[921]),  .coef_in(coef[128]), .rdup_out(a8_wr[913]), .rdlo_out(a8_wr[921]));
			radix2 #(.width(width)) rd_st7_914  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[914]), .rdlo_in(a7_wr[922]),  .coef_in(coef[256]), .rdup_out(a8_wr[914]), .rdlo_out(a8_wr[922]));
			radix2 #(.width(width)) rd_st7_915  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[915]), .rdlo_in(a7_wr[923]),  .coef_in(coef[384]), .rdup_out(a8_wr[915]), .rdlo_out(a8_wr[923]));
			radix2 #(.width(width)) rd_st7_916  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[916]), .rdlo_in(a7_wr[924]),  .coef_in(coef[512]), .rdup_out(a8_wr[916]), .rdlo_out(a8_wr[924]));
			radix2 #(.width(width)) rd_st7_917  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[917]), .rdlo_in(a7_wr[925]),  .coef_in(coef[640]), .rdup_out(a8_wr[917]), .rdlo_out(a8_wr[925]));
			radix2 #(.width(width)) rd_st7_918  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[918]), .rdlo_in(a7_wr[926]),  .coef_in(coef[768]), .rdup_out(a8_wr[918]), .rdlo_out(a8_wr[926]));
			radix2 #(.width(width)) rd_st7_919  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[919]), .rdlo_in(a7_wr[927]),  .coef_in(coef[896]), .rdup_out(a8_wr[919]), .rdlo_out(a8_wr[927]));
			radix2 #(.width(width)) rd_st7_928  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[928]), .rdlo_in(a7_wr[936]),  .coef_in(coef[0]), .rdup_out(a8_wr[928]), .rdlo_out(a8_wr[936]));
			radix2 #(.width(width)) rd_st7_929  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[929]), .rdlo_in(a7_wr[937]),  .coef_in(coef[128]), .rdup_out(a8_wr[929]), .rdlo_out(a8_wr[937]));
			radix2 #(.width(width)) rd_st7_930  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[930]), .rdlo_in(a7_wr[938]),  .coef_in(coef[256]), .rdup_out(a8_wr[930]), .rdlo_out(a8_wr[938]));
			radix2 #(.width(width)) rd_st7_931  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[931]), .rdlo_in(a7_wr[939]),  .coef_in(coef[384]), .rdup_out(a8_wr[931]), .rdlo_out(a8_wr[939]));
			radix2 #(.width(width)) rd_st7_932  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[932]), .rdlo_in(a7_wr[940]),  .coef_in(coef[512]), .rdup_out(a8_wr[932]), .rdlo_out(a8_wr[940]));
			radix2 #(.width(width)) rd_st7_933  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[933]), .rdlo_in(a7_wr[941]),  .coef_in(coef[640]), .rdup_out(a8_wr[933]), .rdlo_out(a8_wr[941]));
			radix2 #(.width(width)) rd_st7_934  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[934]), .rdlo_in(a7_wr[942]),  .coef_in(coef[768]), .rdup_out(a8_wr[934]), .rdlo_out(a8_wr[942]));
			radix2 #(.width(width)) rd_st7_935  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[935]), .rdlo_in(a7_wr[943]),  .coef_in(coef[896]), .rdup_out(a8_wr[935]), .rdlo_out(a8_wr[943]));
			radix2 #(.width(width)) rd_st7_944  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[944]), .rdlo_in(a7_wr[952]),  .coef_in(coef[0]), .rdup_out(a8_wr[944]), .rdlo_out(a8_wr[952]));
			radix2 #(.width(width)) rd_st7_945  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[945]), .rdlo_in(a7_wr[953]),  .coef_in(coef[128]), .rdup_out(a8_wr[945]), .rdlo_out(a8_wr[953]));
			radix2 #(.width(width)) rd_st7_946  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[946]), .rdlo_in(a7_wr[954]),  .coef_in(coef[256]), .rdup_out(a8_wr[946]), .rdlo_out(a8_wr[954]));
			radix2 #(.width(width)) rd_st7_947  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[947]), .rdlo_in(a7_wr[955]),  .coef_in(coef[384]), .rdup_out(a8_wr[947]), .rdlo_out(a8_wr[955]));
			radix2 #(.width(width)) rd_st7_948  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[948]), .rdlo_in(a7_wr[956]),  .coef_in(coef[512]), .rdup_out(a8_wr[948]), .rdlo_out(a8_wr[956]));
			radix2 #(.width(width)) rd_st7_949  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[949]), .rdlo_in(a7_wr[957]),  .coef_in(coef[640]), .rdup_out(a8_wr[949]), .rdlo_out(a8_wr[957]));
			radix2 #(.width(width)) rd_st7_950  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[950]), .rdlo_in(a7_wr[958]),  .coef_in(coef[768]), .rdup_out(a8_wr[950]), .rdlo_out(a8_wr[958]));
			radix2 #(.width(width)) rd_st7_951  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[951]), .rdlo_in(a7_wr[959]),  .coef_in(coef[896]), .rdup_out(a8_wr[951]), .rdlo_out(a8_wr[959]));
			radix2 #(.width(width)) rd_st7_960  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[960]), .rdlo_in(a7_wr[968]),  .coef_in(coef[0]), .rdup_out(a8_wr[960]), .rdlo_out(a8_wr[968]));
			radix2 #(.width(width)) rd_st7_961  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[961]), .rdlo_in(a7_wr[969]),  .coef_in(coef[128]), .rdup_out(a8_wr[961]), .rdlo_out(a8_wr[969]));
			radix2 #(.width(width)) rd_st7_962  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[962]), .rdlo_in(a7_wr[970]),  .coef_in(coef[256]), .rdup_out(a8_wr[962]), .rdlo_out(a8_wr[970]));
			radix2 #(.width(width)) rd_st7_963  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[963]), .rdlo_in(a7_wr[971]),  .coef_in(coef[384]), .rdup_out(a8_wr[963]), .rdlo_out(a8_wr[971]));
			radix2 #(.width(width)) rd_st7_964  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[964]), .rdlo_in(a7_wr[972]),  .coef_in(coef[512]), .rdup_out(a8_wr[964]), .rdlo_out(a8_wr[972]));
			radix2 #(.width(width)) rd_st7_965  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[965]), .rdlo_in(a7_wr[973]),  .coef_in(coef[640]), .rdup_out(a8_wr[965]), .rdlo_out(a8_wr[973]));
			radix2 #(.width(width)) rd_st7_966  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[966]), .rdlo_in(a7_wr[974]),  .coef_in(coef[768]), .rdup_out(a8_wr[966]), .rdlo_out(a8_wr[974]));
			radix2 #(.width(width)) rd_st7_967  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[967]), .rdlo_in(a7_wr[975]),  .coef_in(coef[896]), .rdup_out(a8_wr[967]), .rdlo_out(a8_wr[975]));
			radix2 #(.width(width)) rd_st7_976  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[976]), .rdlo_in(a7_wr[984]),  .coef_in(coef[0]), .rdup_out(a8_wr[976]), .rdlo_out(a8_wr[984]));
			radix2 #(.width(width)) rd_st7_977  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[977]), .rdlo_in(a7_wr[985]),  .coef_in(coef[128]), .rdup_out(a8_wr[977]), .rdlo_out(a8_wr[985]));
			radix2 #(.width(width)) rd_st7_978  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[978]), .rdlo_in(a7_wr[986]),  .coef_in(coef[256]), .rdup_out(a8_wr[978]), .rdlo_out(a8_wr[986]));
			radix2 #(.width(width)) rd_st7_979  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[979]), .rdlo_in(a7_wr[987]),  .coef_in(coef[384]), .rdup_out(a8_wr[979]), .rdlo_out(a8_wr[987]));
			radix2 #(.width(width)) rd_st7_980  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[980]), .rdlo_in(a7_wr[988]),  .coef_in(coef[512]), .rdup_out(a8_wr[980]), .rdlo_out(a8_wr[988]));
			radix2 #(.width(width)) rd_st7_981  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[981]), .rdlo_in(a7_wr[989]),  .coef_in(coef[640]), .rdup_out(a8_wr[981]), .rdlo_out(a8_wr[989]));
			radix2 #(.width(width)) rd_st7_982  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[982]), .rdlo_in(a7_wr[990]),  .coef_in(coef[768]), .rdup_out(a8_wr[982]), .rdlo_out(a8_wr[990]));
			radix2 #(.width(width)) rd_st7_983  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[983]), .rdlo_in(a7_wr[991]),  .coef_in(coef[896]), .rdup_out(a8_wr[983]), .rdlo_out(a8_wr[991]));
			radix2 #(.width(width)) rd_st7_992  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[992]), .rdlo_in(a7_wr[1000]),  .coef_in(coef[0]), .rdup_out(a8_wr[992]), .rdlo_out(a8_wr[1000]));
			radix2 #(.width(width)) rd_st7_993  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[993]), .rdlo_in(a7_wr[1001]),  .coef_in(coef[128]), .rdup_out(a8_wr[993]), .rdlo_out(a8_wr[1001]));
			radix2 #(.width(width)) rd_st7_994  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[994]), .rdlo_in(a7_wr[1002]),  .coef_in(coef[256]), .rdup_out(a8_wr[994]), .rdlo_out(a8_wr[1002]));
			radix2 #(.width(width)) rd_st7_995  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[995]), .rdlo_in(a7_wr[1003]),  .coef_in(coef[384]), .rdup_out(a8_wr[995]), .rdlo_out(a8_wr[1003]));
			radix2 #(.width(width)) rd_st7_996  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[996]), .rdlo_in(a7_wr[1004]),  .coef_in(coef[512]), .rdup_out(a8_wr[996]), .rdlo_out(a8_wr[1004]));
			radix2 #(.width(width)) rd_st7_997  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[997]), .rdlo_in(a7_wr[1005]),  .coef_in(coef[640]), .rdup_out(a8_wr[997]), .rdlo_out(a8_wr[1005]));
			radix2 #(.width(width)) rd_st7_998  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[998]), .rdlo_in(a7_wr[1006]),  .coef_in(coef[768]), .rdup_out(a8_wr[998]), .rdlo_out(a8_wr[1006]));
			radix2 #(.width(width)) rd_st7_999  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[999]), .rdlo_in(a7_wr[1007]),  .coef_in(coef[896]), .rdup_out(a8_wr[999]), .rdlo_out(a8_wr[1007]));
			radix2 #(.width(width)) rd_st7_1008  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1008]), .rdlo_in(a7_wr[1016]),  .coef_in(coef[0]), .rdup_out(a8_wr[1008]), .rdlo_out(a8_wr[1016]));
			radix2 #(.width(width)) rd_st7_1009  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1009]), .rdlo_in(a7_wr[1017]),  .coef_in(coef[128]), .rdup_out(a8_wr[1009]), .rdlo_out(a8_wr[1017]));
			radix2 #(.width(width)) rd_st7_1010  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1010]), .rdlo_in(a7_wr[1018]),  .coef_in(coef[256]), .rdup_out(a8_wr[1010]), .rdlo_out(a8_wr[1018]));
			radix2 #(.width(width)) rd_st7_1011  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1011]), .rdlo_in(a7_wr[1019]),  .coef_in(coef[384]), .rdup_out(a8_wr[1011]), .rdlo_out(a8_wr[1019]));
			radix2 #(.width(width)) rd_st7_1012  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1012]), .rdlo_in(a7_wr[1020]),  .coef_in(coef[512]), .rdup_out(a8_wr[1012]), .rdlo_out(a8_wr[1020]));
			radix2 #(.width(width)) rd_st7_1013  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1013]), .rdlo_in(a7_wr[1021]),  .coef_in(coef[640]), .rdup_out(a8_wr[1013]), .rdlo_out(a8_wr[1021]));
			radix2 #(.width(width)) rd_st7_1014  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1014]), .rdlo_in(a7_wr[1022]),  .coef_in(coef[768]), .rdup_out(a8_wr[1014]), .rdlo_out(a8_wr[1022]));
			radix2 #(.width(width)) rd_st7_1015  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1015]), .rdlo_in(a7_wr[1023]),  .coef_in(coef[896]), .rdup_out(a8_wr[1015]), .rdlo_out(a8_wr[1023]));
			radix2 #(.width(width)) rd_st7_1024  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1024]), .rdlo_in(a7_wr[1032]),  .coef_in(coef[0]), .rdup_out(a8_wr[1024]), .rdlo_out(a8_wr[1032]));
			radix2 #(.width(width)) rd_st7_1025  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1025]), .rdlo_in(a7_wr[1033]),  .coef_in(coef[128]), .rdup_out(a8_wr[1025]), .rdlo_out(a8_wr[1033]));
			radix2 #(.width(width)) rd_st7_1026  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1026]), .rdlo_in(a7_wr[1034]),  .coef_in(coef[256]), .rdup_out(a8_wr[1026]), .rdlo_out(a8_wr[1034]));
			radix2 #(.width(width)) rd_st7_1027  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1027]), .rdlo_in(a7_wr[1035]),  .coef_in(coef[384]), .rdup_out(a8_wr[1027]), .rdlo_out(a8_wr[1035]));
			radix2 #(.width(width)) rd_st7_1028  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1028]), .rdlo_in(a7_wr[1036]),  .coef_in(coef[512]), .rdup_out(a8_wr[1028]), .rdlo_out(a8_wr[1036]));
			radix2 #(.width(width)) rd_st7_1029  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1029]), .rdlo_in(a7_wr[1037]),  .coef_in(coef[640]), .rdup_out(a8_wr[1029]), .rdlo_out(a8_wr[1037]));
			radix2 #(.width(width)) rd_st7_1030  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1030]), .rdlo_in(a7_wr[1038]),  .coef_in(coef[768]), .rdup_out(a8_wr[1030]), .rdlo_out(a8_wr[1038]));
			radix2 #(.width(width)) rd_st7_1031  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1031]), .rdlo_in(a7_wr[1039]),  .coef_in(coef[896]), .rdup_out(a8_wr[1031]), .rdlo_out(a8_wr[1039]));
			radix2 #(.width(width)) rd_st7_1040  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1040]), .rdlo_in(a7_wr[1048]),  .coef_in(coef[0]), .rdup_out(a8_wr[1040]), .rdlo_out(a8_wr[1048]));
			radix2 #(.width(width)) rd_st7_1041  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1041]), .rdlo_in(a7_wr[1049]),  .coef_in(coef[128]), .rdup_out(a8_wr[1041]), .rdlo_out(a8_wr[1049]));
			radix2 #(.width(width)) rd_st7_1042  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1042]), .rdlo_in(a7_wr[1050]),  .coef_in(coef[256]), .rdup_out(a8_wr[1042]), .rdlo_out(a8_wr[1050]));
			radix2 #(.width(width)) rd_st7_1043  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1043]), .rdlo_in(a7_wr[1051]),  .coef_in(coef[384]), .rdup_out(a8_wr[1043]), .rdlo_out(a8_wr[1051]));
			radix2 #(.width(width)) rd_st7_1044  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1044]), .rdlo_in(a7_wr[1052]),  .coef_in(coef[512]), .rdup_out(a8_wr[1044]), .rdlo_out(a8_wr[1052]));
			radix2 #(.width(width)) rd_st7_1045  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1045]), .rdlo_in(a7_wr[1053]),  .coef_in(coef[640]), .rdup_out(a8_wr[1045]), .rdlo_out(a8_wr[1053]));
			radix2 #(.width(width)) rd_st7_1046  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1046]), .rdlo_in(a7_wr[1054]),  .coef_in(coef[768]), .rdup_out(a8_wr[1046]), .rdlo_out(a8_wr[1054]));
			radix2 #(.width(width)) rd_st7_1047  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1047]), .rdlo_in(a7_wr[1055]),  .coef_in(coef[896]), .rdup_out(a8_wr[1047]), .rdlo_out(a8_wr[1055]));
			radix2 #(.width(width)) rd_st7_1056  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1056]), .rdlo_in(a7_wr[1064]),  .coef_in(coef[0]), .rdup_out(a8_wr[1056]), .rdlo_out(a8_wr[1064]));
			radix2 #(.width(width)) rd_st7_1057  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1057]), .rdlo_in(a7_wr[1065]),  .coef_in(coef[128]), .rdup_out(a8_wr[1057]), .rdlo_out(a8_wr[1065]));
			radix2 #(.width(width)) rd_st7_1058  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1058]), .rdlo_in(a7_wr[1066]),  .coef_in(coef[256]), .rdup_out(a8_wr[1058]), .rdlo_out(a8_wr[1066]));
			radix2 #(.width(width)) rd_st7_1059  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1059]), .rdlo_in(a7_wr[1067]),  .coef_in(coef[384]), .rdup_out(a8_wr[1059]), .rdlo_out(a8_wr[1067]));
			radix2 #(.width(width)) rd_st7_1060  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1060]), .rdlo_in(a7_wr[1068]),  .coef_in(coef[512]), .rdup_out(a8_wr[1060]), .rdlo_out(a8_wr[1068]));
			radix2 #(.width(width)) rd_st7_1061  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1061]), .rdlo_in(a7_wr[1069]),  .coef_in(coef[640]), .rdup_out(a8_wr[1061]), .rdlo_out(a8_wr[1069]));
			radix2 #(.width(width)) rd_st7_1062  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1062]), .rdlo_in(a7_wr[1070]),  .coef_in(coef[768]), .rdup_out(a8_wr[1062]), .rdlo_out(a8_wr[1070]));
			radix2 #(.width(width)) rd_st7_1063  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1063]), .rdlo_in(a7_wr[1071]),  .coef_in(coef[896]), .rdup_out(a8_wr[1063]), .rdlo_out(a8_wr[1071]));
			radix2 #(.width(width)) rd_st7_1072  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1072]), .rdlo_in(a7_wr[1080]),  .coef_in(coef[0]), .rdup_out(a8_wr[1072]), .rdlo_out(a8_wr[1080]));
			radix2 #(.width(width)) rd_st7_1073  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1073]), .rdlo_in(a7_wr[1081]),  .coef_in(coef[128]), .rdup_out(a8_wr[1073]), .rdlo_out(a8_wr[1081]));
			radix2 #(.width(width)) rd_st7_1074  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1074]), .rdlo_in(a7_wr[1082]),  .coef_in(coef[256]), .rdup_out(a8_wr[1074]), .rdlo_out(a8_wr[1082]));
			radix2 #(.width(width)) rd_st7_1075  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1075]), .rdlo_in(a7_wr[1083]),  .coef_in(coef[384]), .rdup_out(a8_wr[1075]), .rdlo_out(a8_wr[1083]));
			radix2 #(.width(width)) rd_st7_1076  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1076]), .rdlo_in(a7_wr[1084]),  .coef_in(coef[512]), .rdup_out(a8_wr[1076]), .rdlo_out(a8_wr[1084]));
			radix2 #(.width(width)) rd_st7_1077  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1077]), .rdlo_in(a7_wr[1085]),  .coef_in(coef[640]), .rdup_out(a8_wr[1077]), .rdlo_out(a8_wr[1085]));
			radix2 #(.width(width)) rd_st7_1078  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1078]), .rdlo_in(a7_wr[1086]),  .coef_in(coef[768]), .rdup_out(a8_wr[1078]), .rdlo_out(a8_wr[1086]));
			radix2 #(.width(width)) rd_st7_1079  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1079]), .rdlo_in(a7_wr[1087]),  .coef_in(coef[896]), .rdup_out(a8_wr[1079]), .rdlo_out(a8_wr[1087]));
			radix2 #(.width(width)) rd_st7_1088  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1088]), .rdlo_in(a7_wr[1096]),  .coef_in(coef[0]), .rdup_out(a8_wr[1088]), .rdlo_out(a8_wr[1096]));
			radix2 #(.width(width)) rd_st7_1089  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1089]), .rdlo_in(a7_wr[1097]),  .coef_in(coef[128]), .rdup_out(a8_wr[1089]), .rdlo_out(a8_wr[1097]));
			radix2 #(.width(width)) rd_st7_1090  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1090]), .rdlo_in(a7_wr[1098]),  .coef_in(coef[256]), .rdup_out(a8_wr[1090]), .rdlo_out(a8_wr[1098]));
			radix2 #(.width(width)) rd_st7_1091  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1091]), .rdlo_in(a7_wr[1099]),  .coef_in(coef[384]), .rdup_out(a8_wr[1091]), .rdlo_out(a8_wr[1099]));
			radix2 #(.width(width)) rd_st7_1092  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1092]), .rdlo_in(a7_wr[1100]),  .coef_in(coef[512]), .rdup_out(a8_wr[1092]), .rdlo_out(a8_wr[1100]));
			radix2 #(.width(width)) rd_st7_1093  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1093]), .rdlo_in(a7_wr[1101]),  .coef_in(coef[640]), .rdup_out(a8_wr[1093]), .rdlo_out(a8_wr[1101]));
			radix2 #(.width(width)) rd_st7_1094  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1094]), .rdlo_in(a7_wr[1102]),  .coef_in(coef[768]), .rdup_out(a8_wr[1094]), .rdlo_out(a8_wr[1102]));
			radix2 #(.width(width)) rd_st7_1095  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1095]), .rdlo_in(a7_wr[1103]),  .coef_in(coef[896]), .rdup_out(a8_wr[1095]), .rdlo_out(a8_wr[1103]));
			radix2 #(.width(width)) rd_st7_1104  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1104]), .rdlo_in(a7_wr[1112]),  .coef_in(coef[0]), .rdup_out(a8_wr[1104]), .rdlo_out(a8_wr[1112]));
			radix2 #(.width(width)) rd_st7_1105  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1105]), .rdlo_in(a7_wr[1113]),  .coef_in(coef[128]), .rdup_out(a8_wr[1105]), .rdlo_out(a8_wr[1113]));
			radix2 #(.width(width)) rd_st7_1106  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1106]), .rdlo_in(a7_wr[1114]),  .coef_in(coef[256]), .rdup_out(a8_wr[1106]), .rdlo_out(a8_wr[1114]));
			radix2 #(.width(width)) rd_st7_1107  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1107]), .rdlo_in(a7_wr[1115]),  .coef_in(coef[384]), .rdup_out(a8_wr[1107]), .rdlo_out(a8_wr[1115]));
			radix2 #(.width(width)) rd_st7_1108  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1108]), .rdlo_in(a7_wr[1116]),  .coef_in(coef[512]), .rdup_out(a8_wr[1108]), .rdlo_out(a8_wr[1116]));
			radix2 #(.width(width)) rd_st7_1109  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1109]), .rdlo_in(a7_wr[1117]),  .coef_in(coef[640]), .rdup_out(a8_wr[1109]), .rdlo_out(a8_wr[1117]));
			radix2 #(.width(width)) rd_st7_1110  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1110]), .rdlo_in(a7_wr[1118]),  .coef_in(coef[768]), .rdup_out(a8_wr[1110]), .rdlo_out(a8_wr[1118]));
			radix2 #(.width(width)) rd_st7_1111  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1111]), .rdlo_in(a7_wr[1119]),  .coef_in(coef[896]), .rdup_out(a8_wr[1111]), .rdlo_out(a8_wr[1119]));
			radix2 #(.width(width)) rd_st7_1120  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1120]), .rdlo_in(a7_wr[1128]),  .coef_in(coef[0]), .rdup_out(a8_wr[1120]), .rdlo_out(a8_wr[1128]));
			radix2 #(.width(width)) rd_st7_1121  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1121]), .rdlo_in(a7_wr[1129]),  .coef_in(coef[128]), .rdup_out(a8_wr[1121]), .rdlo_out(a8_wr[1129]));
			radix2 #(.width(width)) rd_st7_1122  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1122]), .rdlo_in(a7_wr[1130]),  .coef_in(coef[256]), .rdup_out(a8_wr[1122]), .rdlo_out(a8_wr[1130]));
			radix2 #(.width(width)) rd_st7_1123  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1123]), .rdlo_in(a7_wr[1131]),  .coef_in(coef[384]), .rdup_out(a8_wr[1123]), .rdlo_out(a8_wr[1131]));
			radix2 #(.width(width)) rd_st7_1124  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1124]), .rdlo_in(a7_wr[1132]),  .coef_in(coef[512]), .rdup_out(a8_wr[1124]), .rdlo_out(a8_wr[1132]));
			radix2 #(.width(width)) rd_st7_1125  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1125]), .rdlo_in(a7_wr[1133]),  .coef_in(coef[640]), .rdup_out(a8_wr[1125]), .rdlo_out(a8_wr[1133]));
			radix2 #(.width(width)) rd_st7_1126  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1126]), .rdlo_in(a7_wr[1134]),  .coef_in(coef[768]), .rdup_out(a8_wr[1126]), .rdlo_out(a8_wr[1134]));
			radix2 #(.width(width)) rd_st7_1127  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1127]), .rdlo_in(a7_wr[1135]),  .coef_in(coef[896]), .rdup_out(a8_wr[1127]), .rdlo_out(a8_wr[1135]));
			radix2 #(.width(width)) rd_st7_1136  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1136]), .rdlo_in(a7_wr[1144]),  .coef_in(coef[0]), .rdup_out(a8_wr[1136]), .rdlo_out(a8_wr[1144]));
			radix2 #(.width(width)) rd_st7_1137  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1137]), .rdlo_in(a7_wr[1145]),  .coef_in(coef[128]), .rdup_out(a8_wr[1137]), .rdlo_out(a8_wr[1145]));
			radix2 #(.width(width)) rd_st7_1138  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1138]), .rdlo_in(a7_wr[1146]),  .coef_in(coef[256]), .rdup_out(a8_wr[1138]), .rdlo_out(a8_wr[1146]));
			radix2 #(.width(width)) rd_st7_1139  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1139]), .rdlo_in(a7_wr[1147]),  .coef_in(coef[384]), .rdup_out(a8_wr[1139]), .rdlo_out(a8_wr[1147]));
			radix2 #(.width(width)) rd_st7_1140  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1140]), .rdlo_in(a7_wr[1148]),  .coef_in(coef[512]), .rdup_out(a8_wr[1140]), .rdlo_out(a8_wr[1148]));
			radix2 #(.width(width)) rd_st7_1141  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1141]), .rdlo_in(a7_wr[1149]),  .coef_in(coef[640]), .rdup_out(a8_wr[1141]), .rdlo_out(a8_wr[1149]));
			radix2 #(.width(width)) rd_st7_1142  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1142]), .rdlo_in(a7_wr[1150]),  .coef_in(coef[768]), .rdup_out(a8_wr[1142]), .rdlo_out(a8_wr[1150]));
			radix2 #(.width(width)) rd_st7_1143  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1143]), .rdlo_in(a7_wr[1151]),  .coef_in(coef[896]), .rdup_out(a8_wr[1143]), .rdlo_out(a8_wr[1151]));
			radix2 #(.width(width)) rd_st7_1152  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1152]), .rdlo_in(a7_wr[1160]),  .coef_in(coef[0]), .rdup_out(a8_wr[1152]), .rdlo_out(a8_wr[1160]));
			radix2 #(.width(width)) rd_st7_1153  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1153]), .rdlo_in(a7_wr[1161]),  .coef_in(coef[128]), .rdup_out(a8_wr[1153]), .rdlo_out(a8_wr[1161]));
			radix2 #(.width(width)) rd_st7_1154  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1154]), .rdlo_in(a7_wr[1162]),  .coef_in(coef[256]), .rdup_out(a8_wr[1154]), .rdlo_out(a8_wr[1162]));
			radix2 #(.width(width)) rd_st7_1155  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1155]), .rdlo_in(a7_wr[1163]),  .coef_in(coef[384]), .rdup_out(a8_wr[1155]), .rdlo_out(a8_wr[1163]));
			radix2 #(.width(width)) rd_st7_1156  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1156]), .rdlo_in(a7_wr[1164]),  .coef_in(coef[512]), .rdup_out(a8_wr[1156]), .rdlo_out(a8_wr[1164]));
			radix2 #(.width(width)) rd_st7_1157  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1157]), .rdlo_in(a7_wr[1165]),  .coef_in(coef[640]), .rdup_out(a8_wr[1157]), .rdlo_out(a8_wr[1165]));
			radix2 #(.width(width)) rd_st7_1158  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1158]), .rdlo_in(a7_wr[1166]),  .coef_in(coef[768]), .rdup_out(a8_wr[1158]), .rdlo_out(a8_wr[1166]));
			radix2 #(.width(width)) rd_st7_1159  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1159]), .rdlo_in(a7_wr[1167]),  .coef_in(coef[896]), .rdup_out(a8_wr[1159]), .rdlo_out(a8_wr[1167]));
			radix2 #(.width(width)) rd_st7_1168  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1168]), .rdlo_in(a7_wr[1176]),  .coef_in(coef[0]), .rdup_out(a8_wr[1168]), .rdlo_out(a8_wr[1176]));
			radix2 #(.width(width)) rd_st7_1169  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1169]), .rdlo_in(a7_wr[1177]),  .coef_in(coef[128]), .rdup_out(a8_wr[1169]), .rdlo_out(a8_wr[1177]));
			radix2 #(.width(width)) rd_st7_1170  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1170]), .rdlo_in(a7_wr[1178]),  .coef_in(coef[256]), .rdup_out(a8_wr[1170]), .rdlo_out(a8_wr[1178]));
			radix2 #(.width(width)) rd_st7_1171  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1171]), .rdlo_in(a7_wr[1179]),  .coef_in(coef[384]), .rdup_out(a8_wr[1171]), .rdlo_out(a8_wr[1179]));
			radix2 #(.width(width)) rd_st7_1172  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1172]), .rdlo_in(a7_wr[1180]),  .coef_in(coef[512]), .rdup_out(a8_wr[1172]), .rdlo_out(a8_wr[1180]));
			radix2 #(.width(width)) rd_st7_1173  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1173]), .rdlo_in(a7_wr[1181]),  .coef_in(coef[640]), .rdup_out(a8_wr[1173]), .rdlo_out(a8_wr[1181]));
			radix2 #(.width(width)) rd_st7_1174  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1174]), .rdlo_in(a7_wr[1182]),  .coef_in(coef[768]), .rdup_out(a8_wr[1174]), .rdlo_out(a8_wr[1182]));
			radix2 #(.width(width)) rd_st7_1175  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1175]), .rdlo_in(a7_wr[1183]),  .coef_in(coef[896]), .rdup_out(a8_wr[1175]), .rdlo_out(a8_wr[1183]));
			radix2 #(.width(width)) rd_st7_1184  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1184]), .rdlo_in(a7_wr[1192]),  .coef_in(coef[0]), .rdup_out(a8_wr[1184]), .rdlo_out(a8_wr[1192]));
			radix2 #(.width(width)) rd_st7_1185  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1185]), .rdlo_in(a7_wr[1193]),  .coef_in(coef[128]), .rdup_out(a8_wr[1185]), .rdlo_out(a8_wr[1193]));
			radix2 #(.width(width)) rd_st7_1186  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1186]), .rdlo_in(a7_wr[1194]),  .coef_in(coef[256]), .rdup_out(a8_wr[1186]), .rdlo_out(a8_wr[1194]));
			radix2 #(.width(width)) rd_st7_1187  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1187]), .rdlo_in(a7_wr[1195]),  .coef_in(coef[384]), .rdup_out(a8_wr[1187]), .rdlo_out(a8_wr[1195]));
			radix2 #(.width(width)) rd_st7_1188  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1188]), .rdlo_in(a7_wr[1196]),  .coef_in(coef[512]), .rdup_out(a8_wr[1188]), .rdlo_out(a8_wr[1196]));
			radix2 #(.width(width)) rd_st7_1189  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1189]), .rdlo_in(a7_wr[1197]),  .coef_in(coef[640]), .rdup_out(a8_wr[1189]), .rdlo_out(a8_wr[1197]));
			radix2 #(.width(width)) rd_st7_1190  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1190]), .rdlo_in(a7_wr[1198]),  .coef_in(coef[768]), .rdup_out(a8_wr[1190]), .rdlo_out(a8_wr[1198]));
			radix2 #(.width(width)) rd_st7_1191  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1191]), .rdlo_in(a7_wr[1199]),  .coef_in(coef[896]), .rdup_out(a8_wr[1191]), .rdlo_out(a8_wr[1199]));
			radix2 #(.width(width)) rd_st7_1200  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1200]), .rdlo_in(a7_wr[1208]),  .coef_in(coef[0]), .rdup_out(a8_wr[1200]), .rdlo_out(a8_wr[1208]));
			radix2 #(.width(width)) rd_st7_1201  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1201]), .rdlo_in(a7_wr[1209]),  .coef_in(coef[128]), .rdup_out(a8_wr[1201]), .rdlo_out(a8_wr[1209]));
			radix2 #(.width(width)) rd_st7_1202  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1202]), .rdlo_in(a7_wr[1210]),  .coef_in(coef[256]), .rdup_out(a8_wr[1202]), .rdlo_out(a8_wr[1210]));
			radix2 #(.width(width)) rd_st7_1203  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1203]), .rdlo_in(a7_wr[1211]),  .coef_in(coef[384]), .rdup_out(a8_wr[1203]), .rdlo_out(a8_wr[1211]));
			radix2 #(.width(width)) rd_st7_1204  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1204]), .rdlo_in(a7_wr[1212]),  .coef_in(coef[512]), .rdup_out(a8_wr[1204]), .rdlo_out(a8_wr[1212]));
			radix2 #(.width(width)) rd_st7_1205  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1205]), .rdlo_in(a7_wr[1213]),  .coef_in(coef[640]), .rdup_out(a8_wr[1205]), .rdlo_out(a8_wr[1213]));
			radix2 #(.width(width)) rd_st7_1206  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1206]), .rdlo_in(a7_wr[1214]),  .coef_in(coef[768]), .rdup_out(a8_wr[1206]), .rdlo_out(a8_wr[1214]));
			radix2 #(.width(width)) rd_st7_1207  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1207]), .rdlo_in(a7_wr[1215]),  .coef_in(coef[896]), .rdup_out(a8_wr[1207]), .rdlo_out(a8_wr[1215]));
			radix2 #(.width(width)) rd_st7_1216  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1216]), .rdlo_in(a7_wr[1224]),  .coef_in(coef[0]), .rdup_out(a8_wr[1216]), .rdlo_out(a8_wr[1224]));
			radix2 #(.width(width)) rd_st7_1217  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1217]), .rdlo_in(a7_wr[1225]),  .coef_in(coef[128]), .rdup_out(a8_wr[1217]), .rdlo_out(a8_wr[1225]));
			radix2 #(.width(width)) rd_st7_1218  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1218]), .rdlo_in(a7_wr[1226]),  .coef_in(coef[256]), .rdup_out(a8_wr[1218]), .rdlo_out(a8_wr[1226]));
			radix2 #(.width(width)) rd_st7_1219  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1219]), .rdlo_in(a7_wr[1227]),  .coef_in(coef[384]), .rdup_out(a8_wr[1219]), .rdlo_out(a8_wr[1227]));
			radix2 #(.width(width)) rd_st7_1220  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1220]), .rdlo_in(a7_wr[1228]),  .coef_in(coef[512]), .rdup_out(a8_wr[1220]), .rdlo_out(a8_wr[1228]));
			radix2 #(.width(width)) rd_st7_1221  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1221]), .rdlo_in(a7_wr[1229]),  .coef_in(coef[640]), .rdup_out(a8_wr[1221]), .rdlo_out(a8_wr[1229]));
			radix2 #(.width(width)) rd_st7_1222  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1222]), .rdlo_in(a7_wr[1230]),  .coef_in(coef[768]), .rdup_out(a8_wr[1222]), .rdlo_out(a8_wr[1230]));
			radix2 #(.width(width)) rd_st7_1223  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1223]), .rdlo_in(a7_wr[1231]),  .coef_in(coef[896]), .rdup_out(a8_wr[1223]), .rdlo_out(a8_wr[1231]));
			radix2 #(.width(width)) rd_st7_1232  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1232]), .rdlo_in(a7_wr[1240]),  .coef_in(coef[0]), .rdup_out(a8_wr[1232]), .rdlo_out(a8_wr[1240]));
			radix2 #(.width(width)) rd_st7_1233  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1233]), .rdlo_in(a7_wr[1241]),  .coef_in(coef[128]), .rdup_out(a8_wr[1233]), .rdlo_out(a8_wr[1241]));
			radix2 #(.width(width)) rd_st7_1234  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1234]), .rdlo_in(a7_wr[1242]),  .coef_in(coef[256]), .rdup_out(a8_wr[1234]), .rdlo_out(a8_wr[1242]));
			radix2 #(.width(width)) rd_st7_1235  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1235]), .rdlo_in(a7_wr[1243]),  .coef_in(coef[384]), .rdup_out(a8_wr[1235]), .rdlo_out(a8_wr[1243]));
			radix2 #(.width(width)) rd_st7_1236  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1236]), .rdlo_in(a7_wr[1244]),  .coef_in(coef[512]), .rdup_out(a8_wr[1236]), .rdlo_out(a8_wr[1244]));
			radix2 #(.width(width)) rd_st7_1237  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1237]), .rdlo_in(a7_wr[1245]),  .coef_in(coef[640]), .rdup_out(a8_wr[1237]), .rdlo_out(a8_wr[1245]));
			radix2 #(.width(width)) rd_st7_1238  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1238]), .rdlo_in(a7_wr[1246]),  .coef_in(coef[768]), .rdup_out(a8_wr[1238]), .rdlo_out(a8_wr[1246]));
			radix2 #(.width(width)) rd_st7_1239  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1239]), .rdlo_in(a7_wr[1247]),  .coef_in(coef[896]), .rdup_out(a8_wr[1239]), .rdlo_out(a8_wr[1247]));
			radix2 #(.width(width)) rd_st7_1248  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1248]), .rdlo_in(a7_wr[1256]),  .coef_in(coef[0]), .rdup_out(a8_wr[1248]), .rdlo_out(a8_wr[1256]));
			radix2 #(.width(width)) rd_st7_1249  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1249]), .rdlo_in(a7_wr[1257]),  .coef_in(coef[128]), .rdup_out(a8_wr[1249]), .rdlo_out(a8_wr[1257]));
			radix2 #(.width(width)) rd_st7_1250  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1250]), .rdlo_in(a7_wr[1258]),  .coef_in(coef[256]), .rdup_out(a8_wr[1250]), .rdlo_out(a8_wr[1258]));
			radix2 #(.width(width)) rd_st7_1251  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1251]), .rdlo_in(a7_wr[1259]),  .coef_in(coef[384]), .rdup_out(a8_wr[1251]), .rdlo_out(a8_wr[1259]));
			radix2 #(.width(width)) rd_st7_1252  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1252]), .rdlo_in(a7_wr[1260]),  .coef_in(coef[512]), .rdup_out(a8_wr[1252]), .rdlo_out(a8_wr[1260]));
			radix2 #(.width(width)) rd_st7_1253  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1253]), .rdlo_in(a7_wr[1261]),  .coef_in(coef[640]), .rdup_out(a8_wr[1253]), .rdlo_out(a8_wr[1261]));
			radix2 #(.width(width)) rd_st7_1254  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1254]), .rdlo_in(a7_wr[1262]),  .coef_in(coef[768]), .rdup_out(a8_wr[1254]), .rdlo_out(a8_wr[1262]));
			radix2 #(.width(width)) rd_st7_1255  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1255]), .rdlo_in(a7_wr[1263]),  .coef_in(coef[896]), .rdup_out(a8_wr[1255]), .rdlo_out(a8_wr[1263]));
			radix2 #(.width(width)) rd_st7_1264  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1264]), .rdlo_in(a7_wr[1272]),  .coef_in(coef[0]), .rdup_out(a8_wr[1264]), .rdlo_out(a8_wr[1272]));
			radix2 #(.width(width)) rd_st7_1265  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1265]), .rdlo_in(a7_wr[1273]),  .coef_in(coef[128]), .rdup_out(a8_wr[1265]), .rdlo_out(a8_wr[1273]));
			radix2 #(.width(width)) rd_st7_1266  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1266]), .rdlo_in(a7_wr[1274]),  .coef_in(coef[256]), .rdup_out(a8_wr[1266]), .rdlo_out(a8_wr[1274]));
			radix2 #(.width(width)) rd_st7_1267  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1267]), .rdlo_in(a7_wr[1275]),  .coef_in(coef[384]), .rdup_out(a8_wr[1267]), .rdlo_out(a8_wr[1275]));
			radix2 #(.width(width)) rd_st7_1268  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1268]), .rdlo_in(a7_wr[1276]),  .coef_in(coef[512]), .rdup_out(a8_wr[1268]), .rdlo_out(a8_wr[1276]));
			radix2 #(.width(width)) rd_st7_1269  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1269]), .rdlo_in(a7_wr[1277]),  .coef_in(coef[640]), .rdup_out(a8_wr[1269]), .rdlo_out(a8_wr[1277]));
			radix2 #(.width(width)) rd_st7_1270  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1270]), .rdlo_in(a7_wr[1278]),  .coef_in(coef[768]), .rdup_out(a8_wr[1270]), .rdlo_out(a8_wr[1278]));
			radix2 #(.width(width)) rd_st7_1271  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1271]), .rdlo_in(a7_wr[1279]),  .coef_in(coef[896]), .rdup_out(a8_wr[1271]), .rdlo_out(a8_wr[1279]));
			radix2 #(.width(width)) rd_st7_1280  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1280]), .rdlo_in(a7_wr[1288]),  .coef_in(coef[0]), .rdup_out(a8_wr[1280]), .rdlo_out(a8_wr[1288]));
			radix2 #(.width(width)) rd_st7_1281  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1281]), .rdlo_in(a7_wr[1289]),  .coef_in(coef[128]), .rdup_out(a8_wr[1281]), .rdlo_out(a8_wr[1289]));
			radix2 #(.width(width)) rd_st7_1282  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1282]), .rdlo_in(a7_wr[1290]),  .coef_in(coef[256]), .rdup_out(a8_wr[1282]), .rdlo_out(a8_wr[1290]));
			radix2 #(.width(width)) rd_st7_1283  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1283]), .rdlo_in(a7_wr[1291]),  .coef_in(coef[384]), .rdup_out(a8_wr[1283]), .rdlo_out(a8_wr[1291]));
			radix2 #(.width(width)) rd_st7_1284  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1284]), .rdlo_in(a7_wr[1292]),  .coef_in(coef[512]), .rdup_out(a8_wr[1284]), .rdlo_out(a8_wr[1292]));
			radix2 #(.width(width)) rd_st7_1285  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1285]), .rdlo_in(a7_wr[1293]),  .coef_in(coef[640]), .rdup_out(a8_wr[1285]), .rdlo_out(a8_wr[1293]));
			radix2 #(.width(width)) rd_st7_1286  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1286]), .rdlo_in(a7_wr[1294]),  .coef_in(coef[768]), .rdup_out(a8_wr[1286]), .rdlo_out(a8_wr[1294]));
			radix2 #(.width(width)) rd_st7_1287  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1287]), .rdlo_in(a7_wr[1295]),  .coef_in(coef[896]), .rdup_out(a8_wr[1287]), .rdlo_out(a8_wr[1295]));
			radix2 #(.width(width)) rd_st7_1296  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1296]), .rdlo_in(a7_wr[1304]),  .coef_in(coef[0]), .rdup_out(a8_wr[1296]), .rdlo_out(a8_wr[1304]));
			radix2 #(.width(width)) rd_st7_1297  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1297]), .rdlo_in(a7_wr[1305]),  .coef_in(coef[128]), .rdup_out(a8_wr[1297]), .rdlo_out(a8_wr[1305]));
			radix2 #(.width(width)) rd_st7_1298  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1298]), .rdlo_in(a7_wr[1306]),  .coef_in(coef[256]), .rdup_out(a8_wr[1298]), .rdlo_out(a8_wr[1306]));
			radix2 #(.width(width)) rd_st7_1299  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1299]), .rdlo_in(a7_wr[1307]),  .coef_in(coef[384]), .rdup_out(a8_wr[1299]), .rdlo_out(a8_wr[1307]));
			radix2 #(.width(width)) rd_st7_1300  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1300]), .rdlo_in(a7_wr[1308]),  .coef_in(coef[512]), .rdup_out(a8_wr[1300]), .rdlo_out(a8_wr[1308]));
			radix2 #(.width(width)) rd_st7_1301  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1301]), .rdlo_in(a7_wr[1309]),  .coef_in(coef[640]), .rdup_out(a8_wr[1301]), .rdlo_out(a8_wr[1309]));
			radix2 #(.width(width)) rd_st7_1302  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1302]), .rdlo_in(a7_wr[1310]),  .coef_in(coef[768]), .rdup_out(a8_wr[1302]), .rdlo_out(a8_wr[1310]));
			radix2 #(.width(width)) rd_st7_1303  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1303]), .rdlo_in(a7_wr[1311]),  .coef_in(coef[896]), .rdup_out(a8_wr[1303]), .rdlo_out(a8_wr[1311]));
			radix2 #(.width(width)) rd_st7_1312  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1312]), .rdlo_in(a7_wr[1320]),  .coef_in(coef[0]), .rdup_out(a8_wr[1312]), .rdlo_out(a8_wr[1320]));
			radix2 #(.width(width)) rd_st7_1313  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1313]), .rdlo_in(a7_wr[1321]),  .coef_in(coef[128]), .rdup_out(a8_wr[1313]), .rdlo_out(a8_wr[1321]));
			radix2 #(.width(width)) rd_st7_1314  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1314]), .rdlo_in(a7_wr[1322]),  .coef_in(coef[256]), .rdup_out(a8_wr[1314]), .rdlo_out(a8_wr[1322]));
			radix2 #(.width(width)) rd_st7_1315  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1315]), .rdlo_in(a7_wr[1323]),  .coef_in(coef[384]), .rdup_out(a8_wr[1315]), .rdlo_out(a8_wr[1323]));
			radix2 #(.width(width)) rd_st7_1316  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1316]), .rdlo_in(a7_wr[1324]),  .coef_in(coef[512]), .rdup_out(a8_wr[1316]), .rdlo_out(a8_wr[1324]));
			radix2 #(.width(width)) rd_st7_1317  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1317]), .rdlo_in(a7_wr[1325]),  .coef_in(coef[640]), .rdup_out(a8_wr[1317]), .rdlo_out(a8_wr[1325]));
			radix2 #(.width(width)) rd_st7_1318  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1318]), .rdlo_in(a7_wr[1326]),  .coef_in(coef[768]), .rdup_out(a8_wr[1318]), .rdlo_out(a8_wr[1326]));
			radix2 #(.width(width)) rd_st7_1319  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1319]), .rdlo_in(a7_wr[1327]),  .coef_in(coef[896]), .rdup_out(a8_wr[1319]), .rdlo_out(a8_wr[1327]));
			radix2 #(.width(width)) rd_st7_1328  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1328]), .rdlo_in(a7_wr[1336]),  .coef_in(coef[0]), .rdup_out(a8_wr[1328]), .rdlo_out(a8_wr[1336]));
			radix2 #(.width(width)) rd_st7_1329  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1329]), .rdlo_in(a7_wr[1337]),  .coef_in(coef[128]), .rdup_out(a8_wr[1329]), .rdlo_out(a8_wr[1337]));
			radix2 #(.width(width)) rd_st7_1330  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1330]), .rdlo_in(a7_wr[1338]),  .coef_in(coef[256]), .rdup_out(a8_wr[1330]), .rdlo_out(a8_wr[1338]));
			radix2 #(.width(width)) rd_st7_1331  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1331]), .rdlo_in(a7_wr[1339]),  .coef_in(coef[384]), .rdup_out(a8_wr[1331]), .rdlo_out(a8_wr[1339]));
			radix2 #(.width(width)) rd_st7_1332  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1332]), .rdlo_in(a7_wr[1340]),  .coef_in(coef[512]), .rdup_out(a8_wr[1332]), .rdlo_out(a8_wr[1340]));
			radix2 #(.width(width)) rd_st7_1333  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1333]), .rdlo_in(a7_wr[1341]),  .coef_in(coef[640]), .rdup_out(a8_wr[1333]), .rdlo_out(a8_wr[1341]));
			radix2 #(.width(width)) rd_st7_1334  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1334]), .rdlo_in(a7_wr[1342]),  .coef_in(coef[768]), .rdup_out(a8_wr[1334]), .rdlo_out(a8_wr[1342]));
			radix2 #(.width(width)) rd_st7_1335  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1335]), .rdlo_in(a7_wr[1343]),  .coef_in(coef[896]), .rdup_out(a8_wr[1335]), .rdlo_out(a8_wr[1343]));
			radix2 #(.width(width)) rd_st7_1344  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1344]), .rdlo_in(a7_wr[1352]),  .coef_in(coef[0]), .rdup_out(a8_wr[1344]), .rdlo_out(a8_wr[1352]));
			radix2 #(.width(width)) rd_st7_1345  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1345]), .rdlo_in(a7_wr[1353]),  .coef_in(coef[128]), .rdup_out(a8_wr[1345]), .rdlo_out(a8_wr[1353]));
			radix2 #(.width(width)) rd_st7_1346  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1346]), .rdlo_in(a7_wr[1354]),  .coef_in(coef[256]), .rdup_out(a8_wr[1346]), .rdlo_out(a8_wr[1354]));
			radix2 #(.width(width)) rd_st7_1347  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1347]), .rdlo_in(a7_wr[1355]),  .coef_in(coef[384]), .rdup_out(a8_wr[1347]), .rdlo_out(a8_wr[1355]));
			radix2 #(.width(width)) rd_st7_1348  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1348]), .rdlo_in(a7_wr[1356]),  .coef_in(coef[512]), .rdup_out(a8_wr[1348]), .rdlo_out(a8_wr[1356]));
			radix2 #(.width(width)) rd_st7_1349  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1349]), .rdlo_in(a7_wr[1357]),  .coef_in(coef[640]), .rdup_out(a8_wr[1349]), .rdlo_out(a8_wr[1357]));
			radix2 #(.width(width)) rd_st7_1350  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1350]), .rdlo_in(a7_wr[1358]),  .coef_in(coef[768]), .rdup_out(a8_wr[1350]), .rdlo_out(a8_wr[1358]));
			radix2 #(.width(width)) rd_st7_1351  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1351]), .rdlo_in(a7_wr[1359]),  .coef_in(coef[896]), .rdup_out(a8_wr[1351]), .rdlo_out(a8_wr[1359]));
			radix2 #(.width(width)) rd_st7_1360  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1360]), .rdlo_in(a7_wr[1368]),  .coef_in(coef[0]), .rdup_out(a8_wr[1360]), .rdlo_out(a8_wr[1368]));
			radix2 #(.width(width)) rd_st7_1361  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1361]), .rdlo_in(a7_wr[1369]),  .coef_in(coef[128]), .rdup_out(a8_wr[1361]), .rdlo_out(a8_wr[1369]));
			radix2 #(.width(width)) rd_st7_1362  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1362]), .rdlo_in(a7_wr[1370]),  .coef_in(coef[256]), .rdup_out(a8_wr[1362]), .rdlo_out(a8_wr[1370]));
			radix2 #(.width(width)) rd_st7_1363  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1363]), .rdlo_in(a7_wr[1371]),  .coef_in(coef[384]), .rdup_out(a8_wr[1363]), .rdlo_out(a8_wr[1371]));
			radix2 #(.width(width)) rd_st7_1364  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1364]), .rdlo_in(a7_wr[1372]),  .coef_in(coef[512]), .rdup_out(a8_wr[1364]), .rdlo_out(a8_wr[1372]));
			radix2 #(.width(width)) rd_st7_1365  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1365]), .rdlo_in(a7_wr[1373]),  .coef_in(coef[640]), .rdup_out(a8_wr[1365]), .rdlo_out(a8_wr[1373]));
			radix2 #(.width(width)) rd_st7_1366  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1366]), .rdlo_in(a7_wr[1374]),  .coef_in(coef[768]), .rdup_out(a8_wr[1366]), .rdlo_out(a8_wr[1374]));
			radix2 #(.width(width)) rd_st7_1367  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1367]), .rdlo_in(a7_wr[1375]),  .coef_in(coef[896]), .rdup_out(a8_wr[1367]), .rdlo_out(a8_wr[1375]));
			radix2 #(.width(width)) rd_st7_1376  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1376]), .rdlo_in(a7_wr[1384]),  .coef_in(coef[0]), .rdup_out(a8_wr[1376]), .rdlo_out(a8_wr[1384]));
			radix2 #(.width(width)) rd_st7_1377  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1377]), .rdlo_in(a7_wr[1385]),  .coef_in(coef[128]), .rdup_out(a8_wr[1377]), .rdlo_out(a8_wr[1385]));
			radix2 #(.width(width)) rd_st7_1378  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1378]), .rdlo_in(a7_wr[1386]),  .coef_in(coef[256]), .rdup_out(a8_wr[1378]), .rdlo_out(a8_wr[1386]));
			radix2 #(.width(width)) rd_st7_1379  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1379]), .rdlo_in(a7_wr[1387]),  .coef_in(coef[384]), .rdup_out(a8_wr[1379]), .rdlo_out(a8_wr[1387]));
			radix2 #(.width(width)) rd_st7_1380  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1380]), .rdlo_in(a7_wr[1388]),  .coef_in(coef[512]), .rdup_out(a8_wr[1380]), .rdlo_out(a8_wr[1388]));
			radix2 #(.width(width)) rd_st7_1381  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1381]), .rdlo_in(a7_wr[1389]),  .coef_in(coef[640]), .rdup_out(a8_wr[1381]), .rdlo_out(a8_wr[1389]));
			radix2 #(.width(width)) rd_st7_1382  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1382]), .rdlo_in(a7_wr[1390]),  .coef_in(coef[768]), .rdup_out(a8_wr[1382]), .rdlo_out(a8_wr[1390]));
			radix2 #(.width(width)) rd_st7_1383  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1383]), .rdlo_in(a7_wr[1391]),  .coef_in(coef[896]), .rdup_out(a8_wr[1383]), .rdlo_out(a8_wr[1391]));
			radix2 #(.width(width)) rd_st7_1392  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1392]), .rdlo_in(a7_wr[1400]),  .coef_in(coef[0]), .rdup_out(a8_wr[1392]), .rdlo_out(a8_wr[1400]));
			radix2 #(.width(width)) rd_st7_1393  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1393]), .rdlo_in(a7_wr[1401]),  .coef_in(coef[128]), .rdup_out(a8_wr[1393]), .rdlo_out(a8_wr[1401]));
			radix2 #(.width(width)) rd_st7_1394  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1394]), .rdlo_in(a7_wr[1402]),  .coef_in(coef[256]), .rdup_out(a8_wr[1394]), .rdlo_out(a8_wr[1402]));
			radix2 #(.width(width)) rd_st7_1395  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1395]), .rdlo_in(a7_wr[1403]),  .coef_in(coef[384]), .rdup_out(a8_wr[1395]), .rdlo_out(a8_wr[1403]));
			radix2 #(.width(width)) rd_st7_1396  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1396]), .rdlo_in(a7_wr[1404]),  .coef_in(coef[512]), .rdup_out(a8_wr[1396]), .rdlo_out(a8_wr[1404]));
			radix2 #(.width(width)) rd_st7_1397  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1397]), .rdlo_in(a7_wr[1405]),  .coef_in(coef[640]), .rdup_out(a8_wr[1397]), .rdlo_out(a8_wr[1405]));
			radix2 #(.width(width)) rd_st7_1398  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1398]), .rdlo_in(a7_wr[1406]),  .coef_in(coef[768]), .rdup_out(a8_wr[1398]), .rdlo_out(a8_wr[1406]));
			radix2 #(.width(width)) rd_st7_1399  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1399]), .rdlo_in(a7_wr[1407]),  .coef_in(coef[896]), .rdup_out(a8_wr[1399]), .rdlo_out(a8_wr[1407]));
			radix2 #(.width(width)) rd_st7_1408  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1408]), .rdlo_in(a7_wr[1416]),  .coef_in(coef[0]), .rdup_out(a8_wr[1408]), .rdlo_out(a8_wr[1416]));
			radix2 #(.width(width)) rd_st7_1409  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1409]), .rdlo_in(a7_wr[1417]),  .coef_in(coef[128]), .rdup_out(a8_wr[1409]), .rdlo_out(a8_wr[1417]));
			radix2 #(.width(width)) rd_st7_1410  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1410]), .rdlo_in(a7_wr[1418]),  .coef_in(coef[256]), .rdup_out(a8_wr[1410]), .rdlo_out(a8_wr[1418]));
			radix2 #(.width(width)) rd_st7_1411  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1411]), .rdlo_in(a7_wr[1419]),  .coef_in(coef[384]), .rdup_out(a8_wr[1411]), .rdlo_out(a8_wr[1419]));
			radix2 #(.width(width)) rd_st7_1412  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1412]), .rdlo_in(a7_wr[1420]),  .coef_in(coef[512]), .rdup_out(a8_wr[1412]), .rdlo_out(a8_wr[1420]));
			radix2 #(.width(width)) rd_st7_1413  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1413]), .rdlo_in(a7_wr[1421]),  .coef_in(coef[640]), .rdup_out(a8_wr[1413]), .rdlo_out(a8_wr[1421]));
			radix2 #(.width(width)) rd_st7_1414  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1414]), .rdlo_in(a7_wr[1422]),  .coef_in(coef[768]), .rdup_out(a8_wr[1414]), .rdlo_out(a8_wr[1422]));
			radix2 #(.width(width)) rd_st7_1415  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1415]), .rdlo_in(a7_wr[1423]),  .coef_in(coef[896]), .rdup_out(a8_wr[1415]), .rdlo_out(a8_wr[1423]));
			radix2 #(.width(width)) rd_st7_1424  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1424]), .rdlo_in(a7_wr[1432]),  .coef_in(coef[0]), .rdup_out(a8_wr[1424]), .rdlo_out(a8_wr[1432]));
			radix2 #(.width(width)) rd_st7_1425  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1425]), .rdlo_in(a7_wr[1433]),  .coef_in(coef[128]), .rdup_out(a8_wr[1425]), .rdlo_out(a8_wr[1433]));
			radix2 #(.width(width)) rd_st7_1426  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1426]), .rdlo_in(a7_wr[1434]),  .coef_in(coef[256]), .rdup_out(a8_wr[1426]), .rdlo_out(a8_wr[1434]));
			radix2 #(.width(width)) rd_st7_1427  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1427]), .rdlo_in(a7_wr[1435]),  .coef_in(coef[384]), .rdup_out(a8_wr[1427]), .rdlo_out(a8_wr[1435]));
			radix2 #(.width(width)) rd_st7_1428  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1428]), .rdlo_in(a7_wr[1436]),  .coef_in(coef[512]), .rdup_out(a8_wr[1428]), .rdlo_out(a8_wr[1436]));
			radix2 #(.width(width)) rd_st7_1429  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1429]), .rdlo_in(a7_wr[1437]),  .coef_in(coef[640]), .rdup_out(a8_wr[1429]), .rdlo_out(a8_wr[1437]));
			radix2 #(.width(width)) rd_st7_1430  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1430]), .rdlo_in(a7_wr[1438]),  .coef_in(coef[768]), .rdup_out(a8_wr[1430]), .rdlo_out(a8_wr[1438]));
			radix2 #(.width(width)) rd_st7_1431  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1431]), .rdlo_in(a7_wr[1439]),  .coef_in(coef[896]), .rdup_out(a8_wr[1431]), .rdlo_out(a8_wr[1439]));
			radix2 #(.width(width)) rd_st7_1440  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1440]), .rdlo_in(a7_wr[1448]),  .coef_in(coef[0]), .rdup_out(a8_wr[1440]), .rdlo_out(a8_wr[1448]));
			radix2 #(.width(width)) rd_st7_1441  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1441]), .rdlo_in(a7_wr[1449]),  .coef_in(coef[128]), .rdup_out(a8_wr[1441]), .rdlo_out(a8_wr[1449]));
			radix2 #(.width(width)) rd_st7_1442  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1442]), .rdlo_in(a7_wr[1450]),  .coef_in(coef[256]), .rdup_out(a8_wr[1442]), .rdlo_out(a8_wr[1450]));
			radix2 #(.width(width)) rd_st7_1443  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1443]), .rdlo_in(a7_wr[1451]),  .coef_in(coef[384]), .rdup_out(a8_wr[1443]), .rdlo_out(a8_wr[1451]));
			radix2 #(.width(width)) rd_st7_1444  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1444]), .rdlo_in(a7_wr[1452]),  .coef_in(coef[512]), .rdup_out(a8_wr[1444]), .rdlo_out(a8_wr[1452]));
			radix2 #(.width(width)) rd_st7_1445  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1445]), .rdlo_in(a7_wr[1453]),  .coef_in(coef[640]), .rdup_out(a8_wr[1445]), .rdlo_out(a8_wr[1453]));
			radix2 #(.width(width)) rd_st7_1446  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1446]), .rdlo_in(a7_wr[1454]),  .coef_in(coef[768]), .rdup_out(a8_wr[1446]), .rdlo_out(a8_wr[1454]));
			radix2 #(.width(width)) rd_st7_1447  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1447]), .rdlo_in(a7_wr[1455]),  .coef_in(coef[896]), .rdup_out(a8_wr[1447]), .rdlo_out(a8_wr[1455]));
			radix2 #(.width(width)) rd_st7_1456  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1456]), .rdlo_in(a7_wr[1464]),  .coef_in(coef[0]), .rdup_out(a8_wr[1456]), .rdlo_out(a8_wr[1464]));
			radix2 #(.width(width)) rd_st7_1457  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1457]), .rdlo_in(a7_wr[1465]),  .coef_in(coef[128]), .rdup_out(a8_wr[1457]), .rdlo_out(a8_wr[1465]));
			radix2 #(.width(width)) rd_st7_1458  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1458]), .rdlo_in(a7_wr[1466]),  .coef_in(coef[256]), .rdup_out(a8_wr[1458]), .rdlo_out(a8_wr[1466]));
			radix2 #(.width(width)) rd_st7_1459  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1459]), .rdlo_in(a7_wr[1467]),  .coef_in(coef[384]), .rdup_out(a8_wr[1459]), .rdlo_out(a8_wr[1467]));
			radix2 #(.width(width)) rd_st7_1460  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1460]), .rdlo_in(a7_wr[1468]),  .coef_in(coef[512]), .rdup_out(a8_wr[1460]), .rdlo_out(a8_wr[1468]));
			radix2 #(.width(width)) rd_st7_1461  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1461]), .rdlo_in(a7_wr[1469]),  .coef_in(coef[640]), .rdup_out(a8_wr[1461]), .rdlo_out(a8_wr[1469]));
			radix2 #(.width(width)) rd_st7_1462  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1462]), .rdlo_in(a7_wr[1470]),  .coef_in(coef[768]), .rdup_out(a8_wr[1462]), .rdlo_out(a8_wr[1470]));
			radix2 #(.width(width)) rd_st7_1463  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1463]), .rdlo_in(a7_wr[1471]),  .coef_in(coef[896]), .rdup_out(a8_wr[1463]), .rdlo_out(a8_wr[1471]));
			radix2 #(.width(width)) rd_st7_1472  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1472]), .rdlo_in(a7_wr[1480]),  .coef_in(coef[0]), .rdup_out(a8_wr[1472]), .rdlo_out(a8_wr[1480]));
			radix2 #(.width(width)) rd_st7_1473  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1473]), .rdlo_in(a7_wr[1481]),  .coef_in(coef[128]), .rdup_out(a8_wr[1473]), .rdlo_out(a8_wr[1481]));
			radix2 #(.width(width)) rd_st7_1474  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1474]), .rdlo_in(a7_wr[1482]),  .coef_in(coef[256]), .rdup_out(a8_wr[1474]), .rdlo_out(a8_wr[1482]));
			radix2 #(.width(width)) rd_st7_1475  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1475]), .rdlo_in(a7_wr[1483]),  .coef_in(coef[384]), .rdup_out(a8_wr[1475]), .rdlo_out(a8_wr[1483]));
			radix2 #(.width(width)) rd_st7_1476  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1476]), .rdlo_in(a7_wr[1484]),  .coef_in(coef[512]), .rdup_out(a8_wr[1476]), .rdlo_out(a8_wr[1484]));
			radix2 #(.width(width)) rd_st7_1477  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1477]), .rdlo_in(a7_wr[1485]),  .coef_in(coef[640]), .rdup_out(a8_wr[1477]), .rdlo_out(a8_wr[1485]));
			radix2 #(.width(width)) rd_st7_1478  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1478]), .rdlo_in(a7_wr[1486]),  .coef_in(coef[768]), .rdup_out(a8_wr[1478]), .rdlo_out(a8_wr[1486]));
			radix2 #(.width(width)) rd_st7_1479  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1479]), .rdlo_in(a7_wr[1487]),  .coef_in(coef[896]), .rdup_out(a8_wr[1479]), .rdlo_out(a8_wr[1487]));
			radix2 #(.width(width)) rd_st7_1488  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1488]), .rdlo_in(a7_wr[1496]),  .coef_in(coef[0]), .rdup_out(a8_wr[1488]), .rdlo_out(a8_wr[1496]));
			radix2 #(.width(width)) rd_st7_1489  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1489]), .rdlo_in(a7_wr[1497]),  .coef_in(coef[128]), .rdup_out(a8_wr[1489]), .rdlo_out(a8_wr[1497]));
			radix2 #(.width(width)) rd_st7_1490  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1490]), .rdlo_in(a7_wr[1498]),  .coef_in(coef[256]), .rdup_out(a8_wr[1490]), .rdlo_out(a8_wr[1498]));
			radix2 #(.width(width)) rd_st7_1491  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1491]), .rdlo_in(a7_wr[1499]),  .coef_in(coef[384]), .rdup_out(a8_wr[1491]), .rdlo_out(a8_wr[1499]));
			radix2 #(.width(width)) rd_st7_1492  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1492]), .rdlo_in(a7_wr[1500]),  .coef_in(coef[512]), .rdup_out(a8_wr[1492]), .rdlo_out(a8_wr[1500]));
			radix2 #(.width(width)) rd_st7_1493  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1493]), .rdlo_in(a7_wr[1501]),  .coef_in(coef[640]), .rdup_out(a8_wr[1493]), .rdlo_out(a8_wr[1501]));
			radix2 #(.width(width)) rd_st7_1494  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1494]), .rdlo_in(a7_wr[1502]),  .coef_in(coef[768]), .rdup_out(a8_wr[1494]), .rdlo_out(a8_wr[1502]));
			radix2 #(.width(width)) rd_st7_1495  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1495]), .rdlo_in(a7_wr[1503]),  .coef_in(coef[896]), .rdup_out(a8_wr[1495]), .rdlo_out(a8_wr[1503]));
			radix2 #(.width(width)) rd_st7_1504  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1504]), .rdlo_in(a7_wr[1512]),  .coef_in(coef[0]), .rdup_out(a8_wr[1504]), .rdlo_out(a8_wr[1512]));
			radix2 #(.width(width)) rd_st7_1505  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1505]), .rdlo_in(a7_wr[1513]),  .coef_in(coef[128]), .rdup_out(a8_wr[1505]), .rdlo_out(a8_wr[1513]));
			radix2 #(.width(width)) rd_st7_1506  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1506]), .rdlo_in(a7_wr[1514]),  .coef_in(coef[256]), .rdup_out(a8_wr[1506]), .rdlo_out(a8_wr[1514]));
			radix2 #(.width(width)) rd_st7_1507  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1507]), .rdlo_in(a7_wr[1515]),  .coef_in(coef[384]), .rdup_out(a8_wr[1507]), .rdlo_out(a8_wr[1515]));
			radix2 #(.width(width)) rd_st7_1508  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1508]), .rdlo_in(a7_wr[1516]),  .coef_in(coef[512]), .rdup_out(a8_wr[1508]), .rdlo_out(a8_wr[1516]));
			radix2 #(.width(width)) rd_st7_1509  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1509]), .rdlo_in(a7_wr[1517]),  .coef_in(coef[640]), .rdup_out(a8_wr[1509]), .rdlo_out(a8_wr[1517]));
			radix2 #(.width(width)) rd_st7_1510  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1510]), .rdlo_in(a7_wr[1518]),  .coef_in(coef[768]), .rdup_out(a8_wr[1510]), .rdlo_out(a8_wr[1518]));
			radix2 #(.width(width)) rd_st7_1511  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1511]), .rdlo_in(a7_wr[1519]),  .coef_in(coef[896]), .rdup_out(a8_wr[1511]), .rdlo_out(a8_wr[1519]));
			radix2 #(.width(width)) rd_st7_1520  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1520]), .rdlo_in(a7_wr[1528]),  .coef_in(coef[0]), .rdup_out(a8_wr[1520]), .rdlo_out(a8_wr[1528]));
			radix2 #(.width(width)) rd_st7_1521  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1521]), .rdlo_in(a7_wr[1529]),  .coef_in(coef[128]), .rdup_out(a8_wr[1521]), .rdlo_out(a8_wr[1529]));
			radix2 #(.width(width)) rd_st7_1522  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1522]), .rdlo_in(a7_wr[1530]),  .coef_in(coef[256]), .rdup_out(a8_wr[1522]), .rdlo_out(a8_wr[1530]));
			radix2 #(.width(width)) rd_st7_1523  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1523]), .rdlo_in(a7_wr[1531]),  .coef_in(coef[384]), .rdup_out(a8_wr[1523]), .rdlo_out(a8_wr[1531]));
			radix2 #(.width(width)) rd_st7_1524  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1524]), .rdlo_in(a7_wr[1532]),  .coef_in(coef[512]), .rdup_out(a8_wr[1524]), .rdlo_out(a8_wr[1532]));
			radix2 #(.width(width)) rd_st7_1525  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1525]), .rdlo_in(a7_wr[1533]),  .coef_in(coef[640]), .rdup_out(a8_wr[1525]), .rdlo_out(a8_wr[1533]));
			radix2 #(.width(width)) rd_st7_1526  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1526]), .rdlo_in(a7_wr[1534]),  .coef_in(coef[768]), .rdup_out(a8_wr[1526]), .rdlo_out(a8_wr[1534]));
			radix2 #(.width(width)) rd_st7_1527  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1527]), .rdlo_in(a7_wr[1535]),  .coef_in(coef[896]), .rdup_out(a8_wr[1527]), .rdlo_out(a8_wr[1535]));
			radix2 #(.width(width)) rd_st7_1536  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1536]), .rdlo_in(a7_wr[1544]),  .coef_in(coef[0]), .rdup_out(a8_wr[1536]), .rdlo_out(a8_wr[1544]));
			radix2 #(.width(width)) rd_st7_1537  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1537]), .rdlo_in(a7_wr[1545]),  .coef_in(coef[128]), .rdup_out(a8_wr[1537]), .rdlo_out(a8_wr[1545]));
			radix2 #(.width(width)) rd_st7_1538  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1538]), .rdlo_in(a7_wr[1546]),  .coef_in(coef[256]), .rdup_out(a8_wr[1538]), .rdlo_out(a8_wr[1546]));
			radix2 #(.width(width)) rd_st7_1539  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1539]), .rdlo_in(a7_wr[1547]),  .coef_in(coef[384]), .rdup_out(a8_wr[1539]), .rdlo_out(a8_wr[1547]));
			radix2 #(.width(width)) rd_st7_1540  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1540]), .rdlo_in(a7_wr[1548]),  .coef_in(coef[512]), .rdup_out(a8_wr[1540]), .rdlo_out(a8_wr[1548]));
			radix2 #(.width(width)) rd_st7_1541  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1541]), .rdlo_in(a7_wr[1549]),  .coef_in(coef[640]), .rdup_out(a8_wr[1541]), .rdlo_out(a8_wr[1549]));
			radix2 #(.width(width)) rd_st7_1542  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1542]), .rdlo_in(a7_wr[1550]),  .coef_in(coef[768]), .rdup_out(a8_wr[1542]), .rdlo_out(a8_wr[1550]));
			radix2 #(.width(width)) rd_st7_1543  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1543]), .rdlo_in(a7_wr[1551]),  .coef_in(coef[896]), .rdup_out(a8_wr[1543]), .rdlo_out(a8_wr[1551]));
			radix2 #(.width(width)) rd_st7_1552  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1552]), .rdlo_in(a7_wr[1560]),  .coef_in(coef[0]), .rdup_out(a8_wr[1552]), .rdlo_out(a8_wr[1560]));
			radix2 #(.width(width)) rd_st7_1553  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1553]), .rdlo_in(a7_wr[1561]),  .coef_in(coef[128]), .rdup_out(a8_wr[1553]), .rdlo_out(a8_wr[1561]));
			radix2 #(.width(width)) rd_st7_1554  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1554]), .rdlo_in(a7_wr[1562]),  .coef_in(coef[256]), .rdup_out(a8_wr[1554]), .rdlo_out(a8_wr[1562]));
			radix2 #(.width(width)) rd_st7_1555  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1555]), .rdlo_in(a7_wr[1563]),  .coef_in(coef[384]), .rdup_out(a8_wr[1555]), .rdlo_out(a8_wr[1563]));
			radix2 #(.width(width)) rd_st7_1556  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1556]), .rdlo_in(a7_wr[1564]),  .coef_in(coef[512]), .rdup_out(a8_wr[1556]), .rdlo_out(a8_wr[1564]));
			radix2 #(.width(width)) rd_st7_1557  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1557]), .rdlo_in(a7_wr[1565]),  .coef_in(coef[640]), .rdup_out(a8_wr[1557]), .rdlo_out(a8_wr[1565]));
			radix2 #(.width(width)) rd_st7_1558  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1558]), .rdlo_in(a7_wr[1566]),  .coef_in(coef[768]), .rdup_out(a8_wr[1558]), .rdlo_out(a8_wr[1566]));
			radix2 #(.width(width)) rd_st7_1559  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1559]), .rdlo_in(a7_wr[1567]),  .coef_in(coef[896]), .rdup_out(a8_wr[1559]), .rdlo_out(a8_wr[1567]));
			radix2 #(.width(width)) rd_st7_1568  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1568]), .rdlo_in(a7_wr[1576]),  .coef_in(coef[0]), .rdup_out(a8_wr[1568]), .rdlo_out(a8_wr[1576]));
			radix2 #(.width(width)) rd_st7_1569  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1569]), .rdlo_in(a7_wr[1577]),  .coef_in(coef[128]), .rdup_out(a8_wr[1569]), .rdlo_out(a8_wr[1577]));
			radix2 #(.width(width)) rd_st7_1570  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1570]), .rdlo_in(a7_wr[1578]),  .coef_in(coef[256]), .rdup_out(a8_wr[1570]), .rdlo_out(a8_wr[1578]));
			radix2 #(.width(width)) rd_st7_1571  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1571]), .rdlo_in(a7_wr[1579]),  .coef_in(coef[384]), .rdup_out(a8_wr[1571]), .rdlo_out(a8_wr[1579]));
			radix2 #(.width(width)) rd_st7_1572  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1572]), .rdlo_in(a7_wr[1580]),  .coef_in(coef[512]), .rdup_out(a8_wr[1572]), .rdlo_out(a8_wr[1580]));
			radix2 #(.width(width)) rd_st7_1573  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1573]), .rdlo_in(a7_wr[1581]),  .coef_in(coef[640]), .rdup_out(a8_wr[1573]), .rdlo_out(a8_wr[1581]));
			radix2 #(.width(width)) rd_st7_1574  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1574]), .rdlo_in(a7_wr[1582]),  .coef_in(coef[768]), .rdup_out(a8_wr[1574]), .rdlo_out(a8_wr[1582]));
			radix2 #(.width(width)) rd_st7_1575  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1575]), .rdlo_in(a7_wr[1583]),  .coef_in(coef[896]), .rdup_out(a8_wr[1575]), .rdlo_out(a8_wr[1583]));
			radix2 #(.width(width)) rd_st7_1584  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1584]), .rdlo_in(a7_wr[1592]),  .coef_in(coef[0]), .rdup_out(a8_wr[1584]), .rdlo_out(a8_wr[1592]));
			radix2 #(.width(width)) rd_st7_1585  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1585]), .rdlo_in(a7_wr[1593]),  .coef_in(coef[128]), .rdup_out(a8_wr[1585]), .rdlo_out(a8_wr[1593]));
			radix2 #(.width(width)) rd_st7_1586  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1586]), .rdlo_in(a7_wr[1594]),  .coef_in(coef[256]), .rdup_out(a8_wr[1586]), .rdlo_out(a8_wr[1594]));
			radix2 #(.width(width)) rd_st7_1587  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1587]), .rdlo_in(a7_wr[1595]),  .coef_in(coef[384]), .rdup_out(a8_wr[1587]), .rdlo_out(a8_wr[1595]));
			radix2 #(.width(width)) rd_st7_1588  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1588]), .rdlo_in(a7_wr[1596]),  .coef_in(coef[512]), .rdup_out(a8_wr[1588]), .rdlo_out(a8_wr[1596]));
			radix2 #(.width(width)) rd_st7_1589  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1589]), .rdlo_in(a7_wr[1597]),  .coef_in(coef[640]), .rdup_out(a8_wr[1589]), .rdlo_out(a8_wr[1597]));
			radix2 #(.width(width)) rd_st7_1590  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1590]), .rdlo_in(a7_wr[1598]),  .coef_in(coef[768]), .rdup_out(a8_wr[1590]), .rdlo_out(a8_wr[1598]));
			radix2 #(.width(width)) rd_st7_1591  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1591]), .rdlo_in(a7_wr[1599]),  .coef_in(coef[896]), .rdup_out(a8_wr[1591]), .rdlo_out(a8_wr[1599]));
			radix2 #(.width(width)) rd_st7_1600  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1600]), .rdlo_in(a7_wr[1608]),  .coef_in(coef[0]), .rdup_out(a8_wr[1600]), .rdlo_out(a8_wr[1608]));
			radix2 #(.width(width)) rd_st7_1601  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1601]), .rdlo_in(a7_wr[1609]),  .coef_in(coef[128]), .rdup_out(a8_wr[1601]), .rdlo_out(a8_wr[1609]));
			radix2 #(.width(width)) rd_st7_1602  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1602]), .rdlo_in(a7_wr[1610]),  .coef_in(coef[256]), .rdup_out(a8_wr[1602]), .rdlo_out(a8_wr[1610]));
			radix2 #(.width(width)) rd_st7_1603  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1603]), .rdlo_in(a7_wr[1611]),  .coef_in(coef[384]), .rdup_out(a8_wr[1603]), .rdlo_out(a8_wr[1611]));
			radix2 #(.width(width)) rd_st7_1604  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1604]), .rdlo_in(a7_wr[1612]),  .coef_in(coef[512]), .rdup_out(a8_wr[1604]), .rdlo_out(a8_wr[1612]));
			radix2 #(.width(width)) rd_st7_1605  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1605]), .rdlo_in(a7_wr[1613]),  .coef_in(coef[640]), .rdup_out(a8_wr[1605]), .rdlo_out(a8_wr[1613]));
			radix2 #(.width(width)) rd_st7_1606  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1606]), .rdlo_in(a7_wr[1614]),  .coef_in(coef[768]), .rdup_out(a8_wr[1606]), .rdlo_out(a8_wr[1614]));
			radix2 #(.width(width)) rd_st7_1607  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1607]), .rdlo_in(a7_wr[1615]),  .coef_in(coef[896]), .rdup_out(a8_wr[1607]), .rdlo_out(a8_wr[1615]));
			radix2 #(.width(width)) rd_st7_1616  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1616]), .rdlo_in(a7_wr[1624]),  .coef_in(coef[0]), .rdup_out(a8_wr[1616]), .rdlo_out(a8_wr[1624]));
			radix2 #(.width(width)) rd_st7_1617  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1617]), .rdlo_in(a7_wr[1625]),  .coef_in(coef[128]), .rdup_out(a8_wr[1617]), .rdlo_out(a8_wr[1625]));
			radix2 #(.width(width)) rd_st7_1618  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1618]), .rdlo_in(a7_wr[1626]),  .coef_in(coef[256]), .rdup_out(a8_wr[1618]), .rdlo_out(a8_wr[1626]));
			radix2 #(.width(width)) rd_st7_1619  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1619]), .rdlo_in(a7_wr[1627]),  .coef_in(coef[384]), .rdup_out(a8_wr[1619]), .rdlo_out(a8_wr[1627]));
			radix2 #(.width(width)) rd_st7_1620  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1620]), .rdlo_in(a7_wr[1628]),  .coef_in(coef[512]), .rdup_out(a8_wr[1620]), .rdlo_out(a8_wr[1628]));
			radix2 #(.width(width)) rd_st7_1621  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1621]), .rdlo_in(a7_wr[1629]),  .coef_in(coef[640]), .rdup_out(a8_wr[1621]), .rdlo_out(a8_wr[1629]));
			radix2 #(.width(width)) rd_st7_1622  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1622]), .rdlo_in(a7_wr[1630]),  .coef_in(coef[768]), .rdup_out(a8_wr[1622]), .rdlo_out(a8_wr[1630]));
			radix2 #(.width(width)) rd_st7_1623  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1623]), .rdlo_in(a7_wr[1631]),  .coef_in(coef[896]), .rdup_out(a8_wr[1623]), .rdlo_out(a8_wr[1631]));
			radix2 #(.width(width)) rd_st7_1632  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1632]), .rdlo_in(a7_wr[1640]),  .coef_in(coef[0]), .rdup_out(a8_wr[1632]), .rdlo_out(a8_wr[1640]));
			radix2 #(.width(width)) rd_st7_1633  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1633]), .rdlo_in(a7_wr[1641]),  .coef_in(coef[128]), .rdup_out(a8_wr[1633]), .rdlo_out(a8_wr[1641]));
			radix2 #(.width(width)) rd_st7_1634  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1634]), .rdlo_in(a7_wr[1642]),  .coef_in(coef[256]), .rdup_out(a8_wr[1634]), .rdlo_out(a8_wr[1642]));
			radix2 #(.width(width)) rd_st7_1635  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1635]), .rdlo_in(a7_wr[1643]),  .coef_in(coef[384]), .rdup_out(a8_wr[1635]), .rdlo_out(a8_wr[1643]));
			radix2 #(.width(width)) rd_st7_1636  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1636]), .rdlo_in(a7_wr[1644]),  .coef_in(coef[512]), .rdup_out(a8_wr[1636]), .rdlo_out(a8_wr[1644]));
			radix2 #(.width(width)) rd_st7_1637  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1637]), .rdlo_in(a7_wr[1645]),  .coef_in(coef[640]), .rdup_out(a8_wr[1637]), .rdlo_out(a8_wr[1645]));
			radix2 #(.width(width)) rd_st7_1638  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1638]), .rdlo_in(a7_wr[1646]),  .coef_in(coef[768]), .rdup_out(a8_wr[1638]), .rdlo_out(a8_wr[1646]));
			radix2 #(.width(width)) rd_st7_1639  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1639]), .rdlo_in(a7_wr[1647]),  .coef_in(coef[896]), .rdup_out(a8_wr[1639]), .rdlo_out(a8_wr[1647]));
			radix2 #(.width(width)) rd_st7_1648  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1648]), .rdlo_in(a7_wr[1656]),  .coef_in(coef[0]), .rdup_out(a8_wr[1648]), .rdlo_out(a8_wr[1656]));
			radix2 #(.width(width)) rd_st7_1649  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1649]), .rdlo_in(a7_wr[1657]),  .coef_in(coef[128]), .rdup_out(a8_wr[1649]), .rdlo_out(a8_wr[1657]));
			radix2 #(.width(width)) rd_st7_1650  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1650]), .rdlo_in(a7_wr[1658]),  .coef_in(coef[256]), .rdup_out(a8_wr[1650]), .rdlo_out(a8_wr[1658]));
			radix2 #(.width(width)) rd_st7_1651  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1651]), .rdlo_in(a7_wr[1659]),  .coef_in(coef[384]), .rdup_out(a8_wr[1651]), .rdlo_out(a8_wr[1659]));
			radix2 #(.width(width)) rd_st7_1652  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1652]), .rdlo_in(a7_wr[1660]),  .coef_in(coef[512]), .rdup_out(a8_wr[1652]), .rdlo_out(a8_wr[1660]));
			radix2 #(.width(width)) rd_st7_1653  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1653]), .rdlo_in(a7_wr[1661]),  .coef_in(coef[640]), .rdup_out(a8_wr[1653]), .rdlo_out(a8_wr[1661]));
			radix2 #(.width(width)) rd_st7_1654  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1654]), .rdlo_in(a7_wr[1662]),  .coef_in(coef[768]), .rdup_out(a8_wr[1654]), .rdlo_out(a8_wr[1662]));
			radix2 #(.width(width)) rd_st7_1655  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1655]), .rdlo_in(a7_wr[1663]),  .coef_in(coef[896]), .rdup_out(a8_wr[1655]), .rdlo_out(a8_wr[1663]));
			radix2 #(.width(width)) rd_st7_1664  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1664]), .rdlo_in(a7_wr[1672]),  .coef_in(coef[0]), .rdup_out(a8_wr[1664]), .rdlo_out(a8_wr[1672]));
			radix2 #(.width(width)) rd_st7_1665  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1665]), .rdlo_in(a7_wr[1673]),  .coef_in(coef[128]), .rdup_out(a8_wr[1665]), .rdlo_out(a8_wr[1673]));
			radix2 #(.width(width)) rd_st7_1666  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1666]), .rdlo_in(a7_wr[1674]),  .coef_in(coef[256]), .rdup_out(a8_wr[1666]), .rdlo_out(a8_wr[1674]));
			radix2 #(.width(width)) rd_st7_1667  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1667]), .rdlo_in(a7_wr[1675]),  .coef_in(coef[384]), .rdup_out(a8_wr[1667]), .rdlo_out(a8_wr[1675]));
			radix2 #(.width(width)) rd_st7_1668  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1668]), .rdlo_in(a7_wr[1676]),  .coef_in(coef[512]), .rdup_out(a8_wr[1668]), .rdlo_out(a8_wr[1676]));
			radix2 #(.width(width)) rd_st7_1669  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1669]), .rdlo_in(a7_wr[1677]),  .coef_in(coef[640]), .rdup_out(a8_wr[1669]), .rdlo_out(a8_wr[1677]));
			radix2 #(.width(width)) rd_st7_1670  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1670]), .rdlo_in(a7_wr[1678]),  .coef_in(coef[768]), .rdup_out(a8_wr[1670]), .rdlo_out(a8_wr[1678]));
			radix2 #(.width(width)) rd_st7_1671  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1671]), .rdlo_in(a7_wr[1679]),  .coef_in(coef[896]), .rdup_out(a8_wr[1671]), .rdlo_out(a8_wr[1679]));
			radix2 #(.width(width)) rd_st7_1680  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1680]), .rdlo_in(a7_wr[1688]),  .coef_in(coef[0]), .rdup_out(a8_wr[1680]), .rdlo_out(a8_wr[1688]));
			radix2 #(.width(width)) rd_st7_1681  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1681]), .rdlo_in(a7_wr[1689]),  .coef_in(coef[128]), .rdup_out(a8_wr[1681]), .rdlo_out(a8_wr[1689]));
			radix2 #(.width(width)) rd_st7_1682  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1682]), .rdlo_in(a7_wr[1690]),  .coef_in(coef[256]), .rdup_out(a8_wr[1682]), .rdlo_out(a8_wr[1690]));
			radix2 #(.width(width)) rd_st7_1683  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1683]), .rdlo_in(a7_wr[1691]),  .coef_in(coef[384]), .rdup_out(a8_wr[1683]), .rdlo_out(a8_wr[1691]));
			radix2 #(.width(width)) rd_st7_1684  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1684]), .rdlo_in(a7_wr[1692]),  .coef_in(coef[512]), .rdup_out(a8_wr[1684]), .rdlo_out(a8_wr[1692]));
			radix2 #(.width(width)) rd_st7_1685  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1685]), .rdlo_in(a7_wr[1693]),  .coef_in(coef[640]), .rdup_out(a8_wr[1685]), .rdlo_out(a8_wr[1693]));
			radix2 #(.width(width)) rd_st7_1686  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1686]), .rdlo_in(a7_wr[1694]),  .coef_in(coef[768]), .rdup_out(a8_wr[1686]), .rdlo_out(a8_wr[1694]));
			radix2 #(.width(width)) rd_st7_1687  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1687]), .rdlo_in(a7_wr[1695]),  .coef_in(coef[896]), .rdup_out(a8_wr[1687]), .rdlo_out(a8_wr[1695]));
			radix2 #(.width(width)) rd_st7_1696  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1696]), .rdlo_in(a7_wr[1704]),  .coef_in(coef[0]), .rdup_out(a8_wr[1696]), .rdlo_out(a8_wr[1704]));
			radix2 #(.width(width)) rd_st7_1697  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1697]), .rdlo_in(a7_wr[1705]),  .coef_in(coef[128]), .rdup_out(a8_wr[1697]), .rdlo_out(a8_wr[1705]));
			radix2 #(.width(width)) rd_st7_1698  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1698]), .rdlo_in(a7_wr[1706]),  .coef_in(coef[256]), .rdup_out(a8_wr[1698]), .rdlo_out(a8_wr[1706]));
			radix2 #(.width(width)) rd_st7_1699  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1699]), .rdlo_in(a7_wr[1707]),  .coef_in(coef[384]), .rdup_out(a8_wr[1699]), .rdlo_out(a8_wr[1707]));
			radix2 #(.width(width)) rd_st7_1700  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1700]), .rdlo_in(a7_wr[1708]),  .coef_in(coef[512]), .rdup_out(a8_wr[1700]), .rdlo_out(a8_wr[1708]));
			radix2 #(.width(width)) rd_st7_1701  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1701]), .rdlo_in(a7_wr[1709]),  .coef_in(coef[640]), .rdup_out(a8_wr[1701]), .rdlo_out(a8_wr[1709]));
			radix2 #(.width(width)) rd_st7_1702  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1702]), .rdlo_in(a7_wr[1710]),  .coef_in(coef[768]), .rdup_out(a8_wr[1702]), .rdlo_out(a8_wr[1710]));
			radix2 #(.width(width)) rd_st7_1703  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1703]), .rdlo_in(a7_wr[1711]),  .coef_in(coef[896]), .rdup_out(a8_wr[1703]), .rdlo_out(a8_wr[1711]));
			radix2 #(.width(width)) rd_st7_1712  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1712]), .rdlo_in(a7_wr[1720]),  .coef_in(coef[0]), .rdup_out(a8_wr[1712]), .rdlo_out(a8_wr[1720]));
			radix2 #(.width(width)) rd_st7_1713  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1713]), .rdlo_in(a7_wr[1721]),  .coef_in(coef[128]), .rdup_out(a8_wr[1713]), .rdlo_out(a8_wr[1721]));
			radix2 #(.width(width)) rd_st7_1714  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1714]), .rdlo_in(a7_wr[1722]),  .coef_in(coef[256]), .rdup_out(a8_wr[1714]), .rdlo_out(a8_wr[1722]));
			radix2 #(.width(width)) rd_st7_1715  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1715]), .rdlo_in(a7_wr[1723]),  .coef_in(coef[384]), .rdup_out(a8_wr[1715]), .rdlo_out(a8_wr[1723]));
			radix2 #(.width(width)) rd_st7_1716  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1716]), .rdlo_in(a7_wr[1724]),  .coef_in(coef[512]), .rdup_out(a8_wr[1716]), .rdlo_out(a8_wr[1724]));
			radix2 #(.width(width)) rd_st7_1717  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1717]), .rdlo_in(a7_wr[1725]),  .coef_in(coef[640]), .rdup_out(a8_wr[1717]), .rdlo_out(a8_wr[1725]));
			radix2 #(.width(width)) rd_st7_1718  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1718]), .rdlo_in(a7_wr[1726]),  .coef_in(coef[768]), .rdup_out(a8_wr[1718]), .rdlo_out(a8_wr[1726]));
			radix2 #(.width(width)) rd_st7_1719  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1719]), .rdlo_in(a7_wr[1727]),  .coef_in(coef[896]), .rdup_out(a8_wr[1719]), .rdlo_out(a8_wr[1727]));
			radix2 #(.width(width)) rd_st7_1728  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1728]), .rdlo_in(a7_wr[1736]),  .coef_in(coef[0]), .rdup_out(a8_wr[1728]), .rdlo_out(a8_wr[1736]));
			radix2 #(.width(width)) rd_st7_1729  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1729]), .rdlo_in(a7_wr[1737]),  .coef_in(coef[128]), .rdup_out(a8_wr[1729]), .rdlo_out(a8_wr[1737]));
			radix2 #(.width(width)) rd_st7_1730  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1730]), .rdlo_in(a7_wr[1738]),  .coef_in(coef[256]), .rdup_out(a8_wr[1730]), .rdlo_out(a8_wr[1738]));
			radix2 #(.width(width)) rd_st7_1731  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1731]), .rdlo_in(a7_wr[1739]),  .coef_in(coef[384]), .rdup_out(a8_wr[1731]), .rdlo_out(a8_wr[1739]));
			radix2 #(.width(width)) rd_st7_1732  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1732]), .rdlo_in(a7_wr[1740]),  .coef_in(coef[512]), .rdup_out(a8_wr[1732]), .rdlo_out(a8_wr[1740]));
			radix2 #(.width(width)) rd_st7_1733  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1733]), .rdlo_in(a7_wr[1741]),  .coef_in(coef[640]), .rdup_out(a8_wr[1733]), .rdlo_out(a8_wr[1741]));
			radix2 #(.width(width)) rd_st7_1734  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1734]), .rdlo_in(a7_wr[1742]),  .coef_in(coef[768]), .rdup_out(a8_wr[1734]), .rdlo_out(a8_wr[1742]));
			radix2 #(.width(width)) rd_st7_1735  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1735]), .rdlo_in(a7_wr[1743]),  .coef_in(coef[896]), .rdup_out(a8_wr[1735]), .rdlo_out(a8_wr[1743]));
			radix2 #(.width(width)) rd_st7_1744  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1744]), .rdlo_in(a7_wr[1752]),  .coef_in(coef[0]), .rdup_out(a8_wr[1744]), .rdlo_out(a8_wr[1752]));
			radix2 #(.width(width)) rd_st7_1745  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1745]), .rdlo_in(a7_wr[1753]),  .coef_in(coef[128]), .rdup_out(a8_wr[1745]), .rdlo_out(a8_wr[1753]));
			radix2 #(.width(width)) rd_st7_1746  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1746]), .rdlo_in(a7_wr[1754]),  .coef_in(coef[256]), .rdup_out(a8_wr[1746]), .rdlo_out(a8_wr[1754]));
			radix2 #(.width(width)) rd_st7_1747  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1747]), .rdlo_in(a7_wr[1755]),  .coef_in(coef[384]), .rdup_out(a8_wr[1747]), .rdlo_out(a8_wr[1755]));
			radix2 #(.width(width)) rd_st7_1748  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1748]), .rdlo_in(a7_wr[1756]),  .coef_in(coef[512]), .rdup_out(a8_wr[1748]), .rdlo_out(a8_wr[1756]));
			radix2 #(.width(width)) rd_st7_1749  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1749]), .rdlo_in(a7_wr[1757]),  .coef_in(coef[640]), .rdup_out(a8_wr[1749]), .rdlo_out(a8_wr[1757]));
			radix2 #(.width(width)) rd_st7_1750  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1750]), .rdlo_in(a7_wr[1758]),  .coef_in(coef[768]), .rdup_out(a8_wr[1750]), .rdlo_out(a8_wr[1758]));
			radix2 #(.width(width)) rd_st7_1751  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1751]), .rdlo_in(a7_wr[1759]),  .coef_in(coef[896]), .rdup_out(a8_wr[1751]), .rdlo_out(a8_wr[1759]));
			radix2 #(.width(width)) rd_st7_1760  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1760]), .rdlo_in(a7_wr[1768]),  .coef_in(coef[0]), .rdup_out(a8_wr[1760]), .rdlo_out(a8_wr[1768]));
			radix2 #(.width(width)) rd_st7_1761  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1761]), .rdlo_in(a7_wr[1769]),  .coef_in(coef[128]), .rdup_out(a8_wr[1761]), .rdlo_out(a8_wr[1769]));
			radix2 #(.width(width)) rd_st7_1762  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1762]), .rdlo_in(a7_wr[1770]),  .coef_in(coef[256]), .rdup_out(a8_wr[1762]), .rdlo_out(a8_wr[1770]));
			radix2 #(.width(width)) rd_st7_1763  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1763]), .rdlo_in(a7_wr[1771]),  .coef_in(coef[384]), .rdup_out(a8_wr[1763]), .rdlo_out(a8_wr[1771]));
			radix2 #(.width(width)) rd_st7_1764  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1764]), .rdlo_in(a7_wr[1772]),  .coef_in(coef[512]), .rdup_out(a8_wr[1764]), .rdlo_out(a8_wr[1772]));
			radix2 #(.width(width)) rd_st7_1765  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1765]), .rdlo_in(a7_wr[1773]),  .coef_in(coef[640]), .rdup_out(a8_wr[1765]), .rdlo_out(a8_wr[1773]));
			radix2 #(.width(width)) rd_st7_1766  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1766]), .rdlo_in(a7_wr[1774]),  .coef_in(coef[768]), .rdup_out(a8_wr[1766]), .rdlo_out(a8_wr[1774]));
			radix2 #(.width(width)) rd_st7_1767  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1767]), .rdlo_in(a7_wr[1775]),  .coef_in(coef[896]), .rdup_out(a8_wr[1767]), .rdlo_out(a8_wr[1775]));
			radix2 #(.width(width)) rd_st7_1776  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1776]), .rdlo_in(a7_wr[1784]),  .coef_in(coef[0]), .rdup_out(a8_wr[1776]), .rdlo_out(a8_wr[1784]));
			radix2 #(.width(width)) rd_st7_1777  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1777]), .rdlo_in(a7_wr[1785]),  .coef_in(coef[128]), .rdup_out(a8_wr[1777]), .rdlo_out(a8_wr[1785]));
			radix2 #(.width(width)) rd_st7_1778  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1778]), .rdlo_in(a7_wr[1786]),  .coef_in(coef[256]), .rdup_out(a8_wr[1778]), .rdlo_out(a8_wr[1786]));
			radix2 #(.width(width)) rd_st7_1779  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1779]), .rdlo_in(a7_wr[1787]),  .coef_in(coef[384]), .rdup_out(a8_wr[1779]), .rdlo_out(a8_wr[1787]));
			radix2 #(.width(width)) rd_st7_1780  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1780]), .rdlo_in(a7_wr[1788]),  .coef_in(coef[512]), .rdup_out(a8_wr[1780]), .rdlo_out(a8_wr[1788]));
			radix2 #(.width(width)) rd_st7_1781  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1781]), .rdlo_in(a7_wr[1789]),  .coef_in(coef[640]), .rdup_out(a8_wr[1781]), .rdlo_out(a8_wr[1789]));
			radix2 #(.width(width)) rd_st7_1782  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1782]), .rdlo_in(a7_wr[1790]),  .coef_in(coef[768]), .rdup_out(a8_wr[1782]), .rdlo_out(a8_wr[1790]));
			radix2 #(.width(width)) rd_st7_1783  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1783]), .rdlo_in(a7_wr[1791]),  .coef_in(coef[896]), .rdup_out(a8_wr[1783]), .rdlo_out(a8_wr[1791]));
			radix2 #(.width(width)) rd_st7_1792  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1792]), .rdlo_in(a7_wr[1800]),  .coef_in(coef[0]), .rdup_out(a8_wr[1792]), .rdlo_out(a8_wr[1800]));
			radix2 #(.width(width)) rd_st7_1793  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1793]), .rdlo_in(a7_wr[1801]),  .coef_in(coef[128]), .rdup_out(a8_wr[1793]), .rdlo_out(a8_wr[1801]));
			radix2 #(.width(width)) rd_st7_1794  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1794]), .rdlo_in(a7_wr[1802]),  .coef_in(coef[256]), .rdup_out(a8_wr[1794]), .rdlo_out(a8_wr[1802]));
			radix2 #(.width(width)) rd_st7_1795  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1795]), .rdlo_in(a7_wr[1803]),  .coef_in(coef[384]), .rdup_out(a8_wr[1795]), .rdlo_out(a8_wr[1803]));
			radix2 #(.width(width)) rd_st7_1796  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1796]), .rdlo_in(a7_wr[1804]),  .coef_in(coef[512]), .rdup_out(a8_wr[1796]), .rdlo_out(a8_wr[1804]));
			radix2 #(.width(width)) rd_st7_1797  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1797]), .rdlo_in(a7_wr[1805]),  .coef_in(coef[640]), .rdup_out(a8_wr[1797]), .rdlo_out(a8_wr[1805]));
			radix2 #(.width(width)) rd_st7_1798  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1798]), .rdlo_in(a7_wr[1806]),  .coef_in(coef[768]), .rdup_out(a8_wr[1798]), .rdlo_out(a8_wr[1806]));
			radix2 #(.width(width)) rd_st7_1799  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1799]), .rdlo_in(a7_wr[1807]),  .coef_in(coef[896]), .rdup_out(a8_wr[1799]), .rdlo_out(a8_wr[1807]));
			radix2 #(.width(width)) rd_st7_1808  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1808]), .rdlo_in(a7_wr[1816]),  .coef_in(coef[0]), .rdup_out(a8_wr[1808]), .rdlo_out(a8_wr[1816]));
			radix2 #(.width(width)) rd_st7_1809  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1809]), .rdlo_in(a7_wr[1817]),  .coef_in(coef[128]), .rdup_out(a8_wr[1809]), .rdlo_out(a8_wr[1817]));
			radix2 #(.width(width)) rd_st7_1810  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1810]), .rdlo_in(a7_wr[1818]),  .coef_in(coef[256]), .rdup_out(a8_wr[1810]), .rdlo_out(a8_wr[1818]));
			radix2 #(.width(width)) rd_st7_1811  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1811]), .rdlo_in(a7_wr[1819]),  .coef_in(coef[384]), .rdup_out(a8_wr[1811]), .rdlo_out(a8_wr[1819]));
			radix2 #(.width(width)) rd_st7_1812  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1812]), .rdlo_in(a7_wr[1820]),  .coef_in(coef[512]), .rdup_out(a8_wr[1812]), .rdlo_out(a8_wr[1820]));
			radix2 #(.width(width)) rd_st7_1813  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1813]), .rdlo_in(a7_wr[1821]),  .coef_in(coef[640]), .rdup_out(a8_wr[1813]), .rdlo_out(a8_wr[1821]));
			radix2 #(.width(width)) rd_st7_1814  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1814]), .rdlo_in(a7_wr[1822]),  .coef_in(coef[768]), .rdup_out(a8_wr[1814]), .rdlo_out(a8_wr[1822]));
			radix2 #(.width(width)) rd_st7_1815  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1815]), .rdlo_in(a7_wr[1823]),  .coef_in(coef[896]), .rdup_out(a8_wr[1815]), .rdlo_out(a8_wr[1823]));
			radix2 #(.width(width)) rd_st7_1824  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1824]), .rdlo_in(a7_wr[1832]),  .coef_in(coef[0]), .rdup_out(a8_wr[1824]), .rdlo_out(a8_wr[1832]));
			radix2 #(.width(width)) rd_st7_1825  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1825]), .rdlo_in(a7_wr[1833]),  .coef_in(coef[128]), .rdup_out(a8_wr[1825]), .rdlo_out(a8_wr[1833]));
			radix2 #(.width(width)) rd_st7_1826  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1826]), .rdlo_in(a7_wr[1834]),  .coef_in(coef[256]), .rdup_out(a8_wr[1826]), .rdlo_out(a8_wr[1834]));
			radix2 #(.width(width)) rd_st7_1827  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1827]), .rdlo_in(a7_wr[1835]),  .coef_in(coef[384]), .rdup_out(a8_wr[1827]), .rdlo_out(a8_wr[1835]));
			radix2 #(.width(width)) rd_st7_1828  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1828]), .rdlo_in(a7_wr[1836]),  .coef_in(coef[512]), .rdup_out(a8_wr[1828]), .rdlo_out(a8_wr[1836]));
			radix2 #(.width(width)) rd_st7_1829  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1829]), .rdlo_in(a7_wr[1837]),  .coef_in(coef[640]), .rdup_out(a8_wr[1829]), .rdlo_out(a8_wr[1837]));
			radix2 #(.width(width)) rd_st7_1830  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1830]), .rdlo_in(a7_wr[1838]),  .coef_in(coef[768]), .rdup_out(a8_wr[1830]), .rdlo_out(a8_wr[1838]));
			radix2 #(.width(width)) rd_st7_1831  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1831]), .rdlo_in(a7_wr[1839]),  .coef_in(coef[896]), .rdup_out(a8_wr[1831]), .rdlo_out(a8_wr[1839]));
			radix2 #(.width(width)) rd_st7_1840  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1840]), .rdlo_in(a7_wr[1848]),  .coef_in(coef[0]), .rdup_out(a8_wr[1840]), .rdlo_out(a8_wr[1848]));
			radix2 #(.width(width)) rd_st7_1841  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1841]), .rdlo_in(a7_wr[1849]),  .coef_in(coef[128]), .rdup_out(a8_wr[1841]), .rdlo_out(a8_wr[1849]));
			radix2 #(.width(width)) rd_st7_1842  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1842]), .rdlo_in(a7_wr[1850]),  .coef_in(coef[256]), .rdup_out(a8_wr[1842]), .rdlo_out(a8_wr[1850]));
			radix2 #(.width(width)) rd_st7_1843  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1843]), .rdlo_in(a7_wr[1851]),  .coef_in(coef[384]), .rdup_out(a8_wr[1843]), .rdlo_out(a8_wr[1851]));
			radix2 #(.width(width)) rd_st7_1844  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1844]), .rdlo_in(a7_wr[1852]),  .coef_in(coef[512]), .rdup_out(a8_wr[1844]), .rdlo_out(a8_wr[1852]));
			radix2 #(.width(width)) rd_st7_1845  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1845]), .rdlo_in(a7_wr[1853]),  .coef_in(coef[640]), .rdup_out(a8_wr[1845]), .rdlo_out(a8_wr[1853]));
			radix2 #(.width(width)) rd_st7_1846  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1846]), .rdlo_in(a7_wr[1854]),  .coef_in(coef[768]), .rdup_out(a8_wr[1846]), .rdlo_out(a8_wr[1854]));
			radix2 #(.width(width)) rd_st7_1847  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1847]), .rdlo_in(a7_wr[1855]),  .coef_in(coef[896]), .rdup_out(a8_wr[1847]), .rdlo_out(a8_wr[1855]));
			radix2 #(.width(width)) rd_st7_1856  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1856]), .rdlo_in(a7_wr[1864]),  .coef_in(coef[0]), .rdup_out(a8_wr[1856]), .rdlo_out(a8_wr[1864]));
			radix2 #(.width(width)) rd_st7_1857  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1857]), .rdlo_in(a7_wr[1865]),  .coef_in(coef[128]), .rdup_out(a8_wr[1857]), .rdlo_out(a8_wr[1865]));
			radix2 #(.width(width)) rd_st7_1858  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1858]), .rdlo_in(a7_wr[1866]),  .coef_in(coef[256]), .rdup_out(a8_wr[1858]), .rdlo_out(a8_wr[1866]));
			radix2 #(.width(width)) rd_st7_1859  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1859]), .rdlo_in(a7_wr[1867]),  .coef_in(coef[384]), .rdup_out(a8_wr[1859]), .rdlo_out(a8_wr[1867]));
			radix2 #(.width(width)) rd_st7_1860  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1860]), .rdlo_in(a7_wr[1868]),  .coef_in(coef[512]), .rdup_out(a8_wr[1860]), .rdlo_out(a8_wr[1868]));
			radix2 #(.width(width)) rd_st7_1861  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1861]), .rdlo_in(a7_wr[1869]),  .coef_in(coef[640]), .rdup_out(a8_wr[1861]), .rdlo_out(a8_wr[1869]));
			radix2 #(.width(width)) rd_st7_1862  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1862]), .rdlo_in(a7_wr[1870]),  .coef_in(coef[768]), .rdup_out(a8_wr[1862]), .rdlo_out(a8_wr[1870]));
			radix2 #(.width(width)) rd_st7_1863  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1863]), .rdlo_in(a7_wr[1871]),  .coef_in(coef[896]), .rdup_out(a8_wr[1863]), .rdlo_out(a8_wr[1871]));
			radix2 #(.width(width)) rd_st7_1872  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1872]), .rdlo_in(a7_wr[1880]),  .coef_in(coef[0]), .rdup_out(a8_wr[1872]), .rdlo_out(a8_wr[1880]));
			radix2 #(.width(width)) rd_st7_1873  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1873]), .rdlo_in(a7_wr[1881]),  .coef_in(coef[128]), .rdup_out(a8_wr[1873]), .rdlo_out(a8_wr[1881]));
			radix2 #(.width(width)) rd_st7_1874  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1874]), .rdlo_in(a7_wr[1882]),  .coef_in(coef[256]), .rdup_out(a8_wr[1874]), .rdlo_out(a8_wr[1882]));
			radix2 #(.width(width)) rd_st7_1875  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1875]), .rdlo_in(a7_wr[1883]),  .coef_in(coef[384]), .rdup_out(a8_wr[1875]), .rdlo_out(a8_wr[1883]));
			radix2 #(.width(width)) rd_st7_1876  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1876]), .rdlo_in(a7_wr[1884]),  .coef_in(coef[512]), .rdup_out(a8_wr[1876]), .rdlo_out(a8_wr[1884]));
			radix2 #(.width(width)) rd_st7_1877  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1877]), .rdlo_in(a7_wr[1885]),  .coef_in(coef[640]), .rdup_out(a8_wr[1877]), .rdlo_out(a8_wr[1885]));
			radix2 #(.width(width)) rd_st7_1878  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1878]), .rdlo_in(a7_wr[1886]),  .coef_in(coef[768]), .rdup_out(a8_wr[1878]), .rdlo_out(a8_wr[1886]));
			radix2 #(.width(width)) rd_st7_1879  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1879]), .rdlo_in(a7_wr[1887]),  .coef_in(coef[896]), .rdup_out(a8_wr[1879]), .rdlo_out(a8_wr[1887]));
			radix2 #(.width(width)) rd_st7_1888  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1888]), .rdlo_in(a7_wr[1896]),  .coef_in(coef[0]), .rdup_out(a8_wr[1888]), .rdlo_out(a8_wr[1896]));
			radix2 #(.width(width)) rd_st7_1889  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1889]), .rdlo_in(a7_wr[1897]),  .coef_in(coef[128]), .rdup_out(a8_wr[1889]), .rdlo_out(a8_wr[1897]));
			radix2 #(.width(width)) rd_st7_1890  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1890]), .rdlo_in(a7_wr[1898]),  .coef_in(coef[256]), .rdup_out(a8_wr[1890]), .rdlo_out(a8_wr[1898]));
			radix2 #(.width(width)) rd_st7_1891  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1891]), .rdlo_in(a7_wr[1899]),  .coef_in(coef[384]), .rdup_out(a8_wr[1891]), .rdlo_out(a8_wr[1899]));
			radix2 #(.width(width)) rd_st7_1892  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1892]), .rdlo_in(a7_wr[1900]),  .coef_in(coef[512]), .rdup_out(a8_wr[1892]), .rdlo_out(a8_wr[1900]));
			radix2 #(.width(width)) rd_st7_1893  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1893]), .rdlo_in(a7_wr[1901]),  .coef_in(coef[640]), .rdup_out(a8_wr[1893]), .rdlo_out(a8_wr[1901]));
			radix2 #(.width(width)) rd_st7_1894  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1894]), .rdlo_in(a7_wr[1902]),  .coef_in(coef[768]), .rdup_out(a8_wr[1894]), .rdlo_out(a8_wr[1902]));
			radix2 #(.width(width)) rd_st7_1895  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1895]), .rdlo_in(a7_wr[1903]),  .coef_in(coef[896]), .rdup_out(a8_wr[1895]), .rdlo_out(a8_wr[1903]));
			radix2 #(.width(width)) rd_st7_1904  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1904]), .rdlo_in(a7_wr[1912]),  .coef_in(coef[0]), .rdup_out(a8_wr[1904]), .rdlo_out(a8_wr[1912]));
			radix2 #(.width(width)) rd_st7_1905  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1905]), .rdlo_in(a7_wr[1913]),  .coef_in(coef[128]), .rdup_out(a8_wr[1905]), .rdlo_out(a8_wr[1913]));
			radix2 #(.width(width)) rd_st7_1906  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1906]), .rdlo_in(a7_wr[1914]),  .coef_in(coef[256]), .rdup_out(a8_wr[1906]), .rdlo_out(a8_wr[1914]));
			radix2 #(.width(width)) rd_st7_1907  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1907]), .rdlo_in(a7_wr[1915]),  .coef_in(coef[384]), .rdup_out(a8_wr[1907]), .rdlo_out(a8_wr[1915]));
			radix2 #(.width(width)) rd_st7_1908  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1908]), .rdlo_in(a7_wr[1916]),  .coef_in(coef[512]), .rdup_out(a8_wr[1908]), .rdlo_out(a8_wr[1916]));
			radix2 #(.width(width)) rd_st7_1909  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1909]), .rdlo_in(a7_wr[1917]),  .coef_in(coef[640]), .rdup_out(a8_wr[1909]), .rdlo_out(a8_wr[1917]));
			radix2 #(.width(width)) rd_st7_1910  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1910]), .rdlo_in(a7_wr[1918]),  .coef_in(coef[768]), .rdup_out(a8_wr[1910]), .rdlo_out(a8_wr[1918]));
			radix2 #(.width(width)) rd_st7_1911  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1911]), .rdlo_in(a7_wr[1919]),  .coef_in(coef[896]), .rdup_out(a8_wr[1911]), .rdlo_out(a8_wr[1919]));
			radix2 #(.width(width)) rd_st7_1920  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1920]), .rdlo_in(a7_wr[1928]),  .coef_in(coef[0]), .rdup_out(a8_wr[1920]), .rdlo_out(a8_wr[1928]));
			radix2 #(.width(width)) rd_st7_1921  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1921]), .rdlo_in(a7_wr[1929]),  .coef_in(coef[128]), .rdup_out(a8_wr[1921]), .rdlo_out(a8_wr[1929]));
			radix2 #(.width(width)) rd_st7_1922  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1922]), .rdlo_in(a7_wr[1930]),  .coef_in(coef[256]), .rdup_out(a8_wr[1922]), .rdlo_out(a8_wr[1930]));
			radix2 #(.width(width)) rd_st7_1923  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1923]), .rdlo_in(a7_wr[1931]),  .coef_in(coef[384]), .rdup_out(a8_wr[1923]), .rdlo_out(a8_wr[1931]));
			radix2 #(.width(width)) rd_st7_1924  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1924]), .rdlo_in(a7_wr[1932]),  .coef_in(coef[512]), .rdup_out(a8_wr[1924]), .rdlo_out(a8_wr[1932]));
			radix2 #(.width(width)) rd_st7_1925  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1925]), .rdlo_in(a7_wr[1933]),  .coef_in(coef[640]), .rdup_out(a8_wr[1925]), .rdlo_out(a8_wr[1933]));
			radix2 #(.width(width)) rd_st7_1926  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1926]), .rdlo_in(a7_wr[1934]),  .coef_in(coef[768]), .rdup_out(a8_wr[1926]), .rdlo_out(a8_wr[1934]));
			radix2 #(.width(width)) rd_st7_1927  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1927]), .rdlo_in(a7_wr[1935]),  .coef_in(coef[896]), .rdup_out(a8_wr[1927]), .rdlo_out(a8_wr[1935]));
			radix2 #(.width(width)) rd_st7_1936  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1936]), .rdlo_in(a7_wr[1944]),  .coef_in(coef[0]), .rdup_out(a8_wr[1936]), .rdlo_out(a8_wr[1944]));
			radix2 #(.width(width)) rd_st7_1937  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1937]), .rdlo_in(a7_wr[1945]),  .coef_in(coef[128]), .rdup_out(a8_wr[1937]), .rdlo_out(a8_wr[1945]));
			radix2 #(.width(width)) rd_st7_1938  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1938]), .rdlo_in(a7_wr[1946]),  .coef_in(coef[256]), .rdup_out(a8_wr[1938]), .rdlo_out(a8_wr[1946]));
			radix2 #(.width(width)) rd_st7_1939  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1939]), .rdlo_in(a7_wr[1947]),  .coef_in(coef[384]), .rdup_out(a8_wr[1939]), .rdlo_out(a8_wr[1947]));
			radix2 #(.width(width)) rd_st7_1940  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1940]), .rdlo_in(a7_wr[1948]),  .coef_in(coef[512]), .rdup_out(a8_wr[1940]), .rdlo_out(a8_wr[1948]));
			radix2 #(.width(width)) rd_st7_1941  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1941]), .rdlo_in(a7_wr[1949]),  .coef_in(coef[640]), .rdup_out(a8_wr[1941]), .rdlo_out(a8_wr[1949]));
			radix2 #(.width(width)) rd_st7_1942  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1942]), .rdlo_in(a7_wr[1950]),  .coef_in(coef[768]), .rdup_out(a8_wr[1942]), .rdlo_out(a8_wr[1950]));
			radix2 #(.width(width)) rd_st7_1943  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1943]), .rdlo_in(a7_wr[1951]),  .coef_in(coef[896]), .rdup_out(a8_wr[1943]), .rdlo_out(a8_wr[1951]));
			radix2 #(.width(width)) rd_st7_1952  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1952]), .rdlo_in(a7_wr[1960]),  .coef_in(coef[0]), .rdup_out(a8_wr[1952]), .rdlo_out(a8_wr[1960]));
			radix2 #(.width(width)) rd_st7_1953  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1953]), .rdlo_in(a7_wr[1961]),  .coef_in(coef[128]), .rdup_out(a8_wr[1953]), .rdlo_out(a8_wr[1961]));
			radix2 #(.width(width)) rd_st7_1954  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1954]), .rdlo_in(a7_wr[1962]),  .coef_in(coef[256]), .rdup_out(a8_wr[1954]), .rdlo_out(a8_wr[1962]));
			radix2 #(.width(width)) rd_st7_1955  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1955]), .rdlo_in(a7_wr[1963]),  .coef_in(coef[384]), .rdup_out(a8_wr[1955]), .rdlo_out(a8_wr[1963]));
			radix2 #(.width(width)) rd_st7_1956  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1956]), .rdlo_in(a7_wr[1964]),  .coef_in(coef[512]), .rdup_out(a8_wr[1956]), .rdlo_out(a8_wr[1964]));
			radix2 #(.width(width)) rd_st7_1957  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1957]), .rdlo_in(a7_wr[1965]),  .coef_in(coef[640]), .rdup_out(a8_wr[1957]), .rdlo_out(a8_wr[1965]));
			radix2 #(.width(width)) rd_st7_1958  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1958]), .rdlo_in(a7_wr[1966]),  .coef_in(coef[768]), .rdup_out(a8_wr[1958]), .rdlo_out(a8_wr[1966]));
			radix2 #(.width(width)) rd_st7_1959  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1959]), .rdlo_in(a7_wr[1967]),  .coef_in(coef[896]), .rdup_out(a8_wr[1959]), .rdlo_out(a8_wr[1967]));
			radix2 #(.width(width)) rd_st7_1968  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1968]), .rdlo_in(a7_wr[1976]),  .coef_in(coef[0]), .rdup_out(a8_wr[1968]), .rdlo_out(a8_wr[1976]));
			radix2 #(.width(width)) rd_st7_1969  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1969]), .rdlo_in(a7_wr[1977]),  .coef_in(coef[128]), .rdup_out(a8_wr[1969]), .rdlo_out(a8_wr[1977]));
			radix2 #(.width(width)) rd_st7_1970  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1970]), .rdlo_in(a7_wr[1978]),  .coef_in(coef[256]), .rdup_out(a8_wr[1970]), .rdlo_out(a8_wr[1978]));
			radix2 #(.width(width)) rd_st7_1971  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1971]), .rdlo_in(a7_wr[1979]),  .coef_in(coef[384]), .rdup_out(a8_wr[1971]), .rdlo_out(a8_wr[1979]));
			radix2 #(.width(width)) rd_st7_1972  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1972]), .rdlo_in(a7_wr[1980]),  .coef_in(coef[512]), .rdup_out(a8_wr[1972]), .rdlo_out(a8_wr[1980]));
			radix2 #(.width(width)) rd_st7_1973  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1973]), .rdlo_in(a7_wr[1981]),  .coef_in(coef[640]), .rdup_out(a8_wr[1973]), .rdlo_out(a8_wr[1981]));
			radix2 #(.width(width)) rd_st7_1974  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1974]), .rdlo_in(a7_wr[1982]),  .coef_in(coef[768]), .rdup_out(a8_wr[1974]), .rdlo_out(a8_wr[1982]));
			radix2 #(.width(width)) rd_st7_1975  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1975]), .rdlo_in(a7_wr[1983]),  .coef_in(coef[896]), .rdup_out(a8_wr[1975]), .rdlo_out(a8_wr[1983]));
			radix2 #(.width(width)) rd_st7_1984  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1984]), .rdlo_in(a7_wr[1992]),  .coef_in(coef[0]), .rdup_out(a8_wr[1984]), .rdlo_out(a8_wr[1992]));
			radix2 #(.width(width)) rd_st7_1985  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1985]), .rdlo_in(a7_wr[1993]),  .coef_in(coef[128]), .rdup_out(a8_wr[1985]), .rdlo_out(a8_wr[1993]));
			radix2 #(.width(width)) rd_st7_1986  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1986]), .rdlo_in(a7_wr[1994]),  .coef_in(coef[256]), .rdup_out(a8_wr[1986]), .rdlo_out(a8_wr[1994]));
			radix2 #(.width(width)) rd_st7_1987  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1987]), .rdlo_in(a7_wr[1995]),  .coef_in(coef[384]), .rdup_out(a8_wr[1987]), .rdlo_out(a8_wr[1995]));
			radix2 #(.width(width)) rd_st7_1988  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1988]), .rdlo_in(a7_wr[1996]),  .coef_in(coef[512]), .rdup_out(a8_wr[1988]), .rdlo_out(a8_wr[1996]));
			radix2 #(.width(width)) rd_st7_1989  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1989]), .rdlo_in(a7_wr[1997]),  .coef_in(coef[640]), .rdup_out(a8_wr[1989]), .rdlo_out(a8_wr[1997]));
			radix2 #(.width(width)) rd_st7_1990  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1990]), .rdlo_in(a7_wr[1998]),  .coef_in(coef[768]), .rdup_out(a8_wr[1990]), .rdlo_out(a8_wr[1998]));
			radix2 #(.width(width)) rd_st7_1991  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[1991]), .rdlo_in(a7_wr[1999]),  .coef_in(coef[896]), .rdup_out(a8_wr[1991]), .rdlo_out(a8_wr[1999]));
			radix2 #(.width(width)) rd_st7_2000  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[2000]), .rdlo_in(a7_wr[2008]),  .coef_in(coef[0]), .rdup_out(a8_wr[2000]), .rdlo_out(a8_wr[2008]));
			radix2 #(.width(width)) rd_st7_2001  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[2001]), .rdlo_in(a7_wr[2009]),  .coef_in(coef[128]), .rdup_out(a8_wr[2001]), .rdlo_out(a8_wr[2009]));
			radix2 #(.width(width)) rd_st7_2002  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[2002]), .rdlo_in(a7_wr[2010]),  .coef_in(coef[256]), .rdup_out(a8_wr[2002]), .rdlo_out(a8_wr[2010]));
			radix2 #(.width(width)) rd_st7_2003  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[2003]), .rdlo_in(a7_wr[2011]),  .coef_in(coef[384]), .rdup_out(a8_wr[2003]), .rdlo_out(a8_wr[2011]));
			radix2 #(.width(width)) rd_st7_2004  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[2004]), .rdlo_in(a7_wr[2012]),  .coef_in(coef[512]), .rdup_out(a8_wr[2004]), .rdlo_out(a8_wr[2012]));
			radix2 #(.width(width)) rd_st7_2005  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[2005]), .rdlo_in(a7_wr[2013]),  .coef_in(coef[640]), .rdup_out(a8_wr[2005]), .rdlo_out(a8_wr[2013]));
			radix2 #(.width(width)) rd_st7_2006  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[2006]), .rdlo_in(a7_wr[2014]),  .coef_in(coef[768]), .rdup_out(a8_wr[2006]), .rdlo_out(a8_wr[2014]));
			radix2 #(.width(width)) rd_st7_2007  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[2007]), .rdlo_in(a7_wr[2015]),  .coef_in(coef[896]), .rdup_out(a8_wr[2007]), .rdlo_out(a8_wr[2015]));
			radix2 #(.width(width)) rd_st7_2016  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[2016]), .rdlo_in(a7_wr[2024]),  .coef_in(coef[0]), .rdup_out(a8_wr[2016]), .rdlo_out(a8_wr[2024]));
			radix2 #(.width(width)) rd_st7_2017  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[2017]), .rdlo_in(a7_wr[2025]),  .coef_in(coef[128]), .rdup_out(a8_wr[2017]), .rdlo_out(a8_wr[2025]));
			radix2 #(.width(width)) rd_st7_2018  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[2018]), .rdlo_in(a7_wr[2026]),  .coef_in(coef[256]), .rdup_out(a8_wr[2018]), .rdlo_out(a8_wr[2026]));
			radix2 #(.width(width)) rd_st7_2019  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[2019]), .rdlo_in(a7_wr[2027]),  .coef_in(coef[384]), .rdup_out(a8_wr[2019]), .rdlo_out(a8_wr[2027]));
			radix2 #(.width(width)) rd_st7_2020  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[2020]), .rdlo_in(a7_wr[2028]),  .coef_in(coef[512]), .rdup_out(a8_wr[2020]), .rdlo_out(a8_wr[2028]));
			radix2 #(.width(width)) rd_st7_2021  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[2021]), .rdlo_in(a7_wr[2029]),  .coef_in(coef[640]), .rdup_out(a8_wr[2021]), .rdlo_out(a8_wr[2029]));
			radix2 #(.width(width)) rd_st7_2022  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[2022]), .rdlo_in(a7_wr[2030]),  .coef_in(coef[768]), .rdup_out(a8_wr[2022]), .rdlo_out(a8_wr[2030]));
			radix2 #(.width(width)) rd_st7_2023  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[2023]), .rdlo_in(a7_wr[2031]),  .coef_in(coef[896]), .rdup_out(a8_wr[2023]), .rdlo_out(a8_wr[2031]));
			radix2 #(.width(width)) rd_st7_2032  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[2032]), .rdlo_in(a7_wr[2040]),  .coef_in(coef[0]), .rdup_out(a8_wr[2032]), .rdlo_out(a8_wr[2040]));
			radix2 #(.width(width)) rd_st7_2033  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[2033]), .rdlo_in(a7_wr[2041]),  .coef_in(coef[128]), .rdup_out(a8_wr[2033]), .rdlo_out(a8_wr[2041]));
			radix2 #(.width(width)) rd_st7_2034  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[2034]), .rdlo_in(a7_wr[2042]),  .coef_in(coef[256]), .rdup_out(a8_wr[2034]), .rdlo_out(a8_wr[2042]));
			radix2 #(.width(width)) rd_st7_2035  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[2035]), .rdlo_in(a7_wr[2043]),  .coef_in(coef[384]), .rdup_out(a8_wr[2035]), .rdlo_out(a8_wr[2043]));
			radix2 #(.width(width)) rd_st7_2036  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[2036]), .rdlo_in(a7_wr[2044]),  .coef_in(coef[512]), .rdup_out(a8_wr[2036]), .rdlo_out(a8_wr[2044]));
			radix2 #(.width(width)) rd_st7_2037  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[2037]), .rdlo_in(a7_wr[2045]),  .coef_in(coef[640]), .rdup_out(a8_wr[2037]), .rdlo_out(a8_wr[2045]));
			radix2 #(.width(width)) rd_st7_2038  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[2038]), .rdlo_in(a7_wr[2046]),  .coef_in(coef[768]), .rdup_out(a8_wr[2038]), .rdlo_out(a8_wr[2046]));
			radix2 #(.width(width)) rd_st7_2039  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a7_wr[2039]), .rdlo_in(a7_wr[2047]),  .coef_in(coef[896]), .rdup_out(a8_wr[2039]), .rdlo_out(a8_wr[2047]));

		//--- radix stage 8
			radix2 #(.width(width)) rd_st8_0   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[0]), .rdlo_in(a8_wr[4]),  .coef_in(coef[0]), .rdup_out(a9_wr[0]), .rdlo_out(a9_wr[4]));
			radix2 #(.width(width)) rd_st8_1   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1]), .rdlo_in(a8_wr[5]),  .coef_in(coef[256]), .rdup_out(a9_wr[1]), .rdlo_out(a9_wr[5]));
			radix2 #(.width(width)) rd_st8_2   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[2]), .rdlo_in(a8_wr[6]),  .coef_in(coef[512]), .rdup_out(a9_wr[2]), .rdlo_out(a9_wr[6]));
			radix2 #(.width(width)) rd_st8_3   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[3]), .rdlo_in(a8_wr[7]),  .coef_in(coef[768]), .rdup_out(a9_wr[3]), .rdlo_out(a9_wr[7]));
			radix2 #(.width(width)) rd_st8_8   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[8]), .rdlo_in(a8_wr[12]),  .coef_in(coef[0]), .rdup_out(a9_wr[8]), .rdlo_out(a9_wr[12]));
			radix2 #(.width(width)) rd_st8_9   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[9]), .rdlo_in(a8_wr[13]),  .coef_in(coef[256]), .rdup_out(a9_wr[9]), .rdlo_out(a9_wr[13]));
			radix2 #(.width(width)) rd_st8_10  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[10]), .rdlo_in(a8_wr[14]),  .coef_in(coef[512]), .rdup_out(a9_wr[10]), .rdlo_out(a9_wr[14]));
			radix2 #(.width(width)) rd_st8_11  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[11]), .rdlo_in(a8_wr[15]),  .coef_in(coef[768]), .rdup_out(a9_wr[11]), .rdlo_out(a9_wr[15]));
			radix2 #(.width(width)) rd_st8_16  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[16]), .rdlo_in(a8_wr[20]),  .coef_in(coef[0]), .rdup_out(a9_wr[16]), .rdlo_out(a9_wr[20]));
			radix2 #(.width(width)) rd_st8_17  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[17]), .rdlo_in(a8_wr[21]),  .coef_in(coef[256]), .rdup_out(a9_wr[17]), .rdlo_out(a9_wr[21]));
			radix2 #(.width(width)) rd_st8_18  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[18]), .rdlo_in(a8_wr[22]),  .coef_in(coef[512]), .rdup_out(a9_wr[18]), .rdlo_out(a9_wr[22]));
			radix2 #(.width(width)) rd_st8_19  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[19]), .rdlo_in(a8_wr[23]),  .coef_in(coef[768]), .rdup_out(a9_wr[19]), .rdlo_out(a9_wr[23]));
			radix2 #(.width(width)) rd_st8_24  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[24]), .rdlo_in(a8_wr[28]),  .coef_in(coef[0]), .rdup_out(a9_wr[24]), .rdlo_out(a9_wr[28]));
			radix2 #(.width(width)) rd_st8_25  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[25]), .rdlo_in(a8_wr[29]),  .coef_in(coef[256]), .rdup_out(a9_wr[25]), .rdlo_out(a9_wr[29]));
			radix2 #(.width(width)) rd_st8_26  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[26]), .rdlo_in(a8_wr[30]),  .coef_in(coef[512]), .rdup_out(a9_wr[26]), .rdlo_out(a9_wr[30]));
			radix2 #(.width(width)) rd_st8_27  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[27]), .rdlo_in(a8_wr[31]),  .coef_in(coef[768]), .rdup_out(a9_wr[27]), .rdlo_out(a9_wr[31]));
			radix2 #(.width(width)) rd_st8_32  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[32]), .rdlo_in(a8_wr[36]),  .coef_in(coef[0]), .rdup_out(a9_wr[32]), .rdlo_out(a9_wr[36]));
			radix2 #(.width(width)) rd_st8_33  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[33]), .rdlo_in(a8_wr[37]),  .coef_in(coef[256]), .rdup_out(a9_wr[33]), .rdlo_out(a9_wr[37]));
			radix2 #(.width(width)) rd_st8_34  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[34]), .rdlo_in(a8_wr[38]),  .coef_in(coef[512]), .rdup_out(a9_wr[34]), .rdlo_out(a9_wr[38]));
			radix2 #(.width(width)) rd_st8_35  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[35]), .rdlo_in(a8_wr[39]),  .coef_in(coef[768]), .rdup_out(a9_wr[35]), .rdlo_out(a9_wr[39]));
			radix2 #(.width(width)) rd_st8_40  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[40]), .rdlo_in(a8_wr[44]),  .coef_in(coef[0]), .rdup_out(a9_wr[40]), .rdlo_out(a9_wr[44]));
			radix2 #(.width(width)) rd_st8_41  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[41]), .rdlo_in(a8_wr[45]),  .coef_in(coef[256]), .rdup_out(a9_wr[41]), .rdlo_out(a9_wr[45]));
			radix2 #(.width(width)) rd_st8_42  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[42]), .rdlo_in(a8_wr[46]),  .coef_in(coef[512]), .rdup_out(a9_wr[42]), .rdlo_out(a9_wr[46]));
			radix2 #(.width(width)) rd_st8_43  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[43]), .rdlo_in(a8_wr[47]),  .coef_in(coef[768]), .rdup_out(a9_wr[43]), .rdlo_out(a9_wr[47]));
			radix2 #(.width(width)) rd_st8_48  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[48]), .rdlo_in(a8_wr[52]),  .coef_in(coef[0]), .rdup_out(a9_wr[48]), .rdlo_out(a9_wr[52]));
			radix2 #(.width(width)) rd_st8_49  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[49]), .rdlo_in(a8_wr[53]),  .coef_in(coef[256]), .rdup_out(a9_wr[49]), .rdlo_out(a9_wr[53]));
			radix2 #(.width(width)) rd_st8_50  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[50]), .rdlo_in(a8_wr[54]),  .coef_in(coef[512]), .rdup_out(a9_wr[50]), .rdlo_out(a9_wr[54]));
			radix2 #(.width(width)) rd_st8_51  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[51]), .rdlo_in(a8_wr[55]),  .coef_in(coef[768]), .rdup_out(a9_wr[51]), .rdlo_out(a9_wr[55]));
			radix2 #(.width(width)) rd_st8_56  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[56]), .rdlo_in(a8_wr[60]),  .coef_in(coef[0]), .rdup_out(a9_wr[56]), .rdlo_out(a9_wr[60]));
			radix2 #(.width(width)) rd_st8_57  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[57]), .rdlo_in(a8_wr[61]),  .coef_in(coef[256]), .rdup_out(a9_wr[57]), .rdlo_out(a9_wr[61]));
			radix2 #(.width(width)) rd_st8_58  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[58]), .rdlo_in(a8_wr[62]),  .coef_in(coef[512]), .rdup_out(a9_wr[58]), .rdlo_out(a9_wr[62]));
			radix2 #(.width(width)) rd_st8_59  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[59]), .rdlo_in(a8_wr[63]),  .coef_in(coef[768]), .rdup_out(a9_wr[59]), .rdlo_out(a9_wr[63]));
			radix2 #(.width(width)) rd_st8_64  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[64]), .rdlo_in(a8_wr[68]),  .coef_in(coef[0]), .rdup_out(a9_wr[64]), .rdlo_out(a9_wr[68]));
			radix2 #(.width(width)) rd_st8_65  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[65]), .rdlo_in(a8_wr[69]),  .coef_in(coef[256]), .rdup_out(a9_wr[65]), .rdlo_out(a9_wr[69]));
			radix2 #(.width(width)) rd_st8_66  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[66]), .rdlo_in(a8_wr[70]),  .coef_in(coef[512]), .rdup_out(a9_wr[66]), .rdlo_out(a9_wr[70]));
			radix2 #(.width(width)) rd_st8_67  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[67]), .rdlo_in(a8_wr[71]),  .coef_in(coef[768]), .rdup_out(a9_wr[67]), .rdlo_out(a9_wr[71]));
			radix2 #(.width(width)) rd_st8_72  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[72]), .rdlo_in(a8_wr[76]),  .coef_in(coef[0]), .rdup_out(a9_wr[72]), .rdlo_out(a9_wr[76]));
			radix2 #(.width(width)) rd_st8_73  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[73]), .rdlo_in(a8_wr[77]),  .coef_in(coef[256]), .rdup_out(a9_wr[73]), .rdlo_out(a9_wr[77]));
			radix2 #(.width(width)) rd_st8_74  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[74]), .rdlo_in(a8_wr[78]),  .coef_in(coef[512]), .rdup_out(a9_wr[74]), .rdlo_out(a9_wr[78]));
			radix2 #(.width(width)) rd_st8_75  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[75]), .rdlo_in(a8_wr[79]),  .coef_in(coef[768]), .rdup_out(a9_wr[75]), .rdlo_out(a9_wr[79]));
			radix2 #(.width(width)) rd_st8_80  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[80]), .rdlo_in(a8_wr[84]),  .coef_in(coef[0]), .rdup_out(a9_wr[80]), .rdlo_out(a9_wr[84]));
			radix2 #(.width(width)) rd_st8_81  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[81]), .rdlo_in(a8_wr[85]),  .coef_in(coef[256]), .rdup_out(a9_wr[81]), .rdlo_out(a9_wr[85]));
			radix2 #(.width(width)) rd_st8_82  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[82]), .rdlo_in(a8_wr[86]),  .coef_in(coef[512]), .rdup_out(a9_wr[82]), .rdlo_out(a9_wr[86]));
			radix2 #(.width(width)) rd_st8_83  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[83]), .rdlo_in(a8_wr[87]),  .coef_in(coef[768]), .rdup_out(a9_wr[83]), .rdlo_out(a9_wr[87]));
			radix2 #(.width(width)) rd_st8_88  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[88]), .rdlo_in(a8_wr[92]),  .coef_in(coef[0]), .rdup_out(a9_wr[88]), .rdlo_out(a9_wr[92]));
			radix2 #(.width(width)) rd_st8_89  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[89]), .rdlo_in(a8_wr[93]),  .coef_in(coef[256]), .rdup_out(a9_wr[89]), .rdlo_out(a9_wr[93]));
			radix2 #(.width(width)) rd_st8_90  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[90]), .rdlo_in(a8_wr[94]),  .coef_in(coef[512]), .rdup_out(a9_wr[90]), .rdlo_out(a9_wr[94]));
			radix2 #(.width(width)) rd_st8_91  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[91]), .rdlo_in(a8_wr[95]),  .coef_in(coef[768]), .rdup_out(a9_wr[91]), .rdlo_out(a9_wr[95]));
			radix2 #(.width(width)) rd_st8_96  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[96]), .rdlo_in(a8_wr[100]),  .coef_in(coef[0]), .rdup_out(a9_wr[96]), .rdlo_out(a9_wr[100]));
			radix2 #(.width(width)) rd_st8_97  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[97]), .rdlo_in(a8_wr[101]),  .coef_in(coef[256]), .rdup_out(a9_wr[97]), .rdlo_out(a9_wr[101]));
			radix2 #(.width(width)) rd_st8_98  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[98]), .rdlo_in(a8_wr[102]),  .coef_in(coef[512]), .rdup_out(a9_wr[98]), .rdlo_out(a9_wr[102]));
			radix2 #(.width(width)) rd_st8_99  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[99]), .rdlo_in(a8_wr[103]),  .coef_in(coef[768]), .rdup_out(a9_wr[99]), .rdlo_out(a9_wr[103]));
			radix2 #(.width(width)) rd_st8_104  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[104]), .rdlo_in(a8_wr[108]),  .coef_in(coef[0]), .rdup_out(a9_wr[104]), .rdlo_out(a9_wr[108]));
			radix2 #(.width(width)) rd_st8_105  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[105]), .rdlo_in(a8_wr[109]),  .coef_in(coef[256]), .rdup_out(a9_wr[105]), .rdlo_out(a9_wr[109]));
			radix2 #(.width(width)) rd_st8_106  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[106]), .rdlo_in(a8_wr[110]),  .coef_in(coef[512]), .rdup_out(a9_wr[106]), .rdlo_out(a9_wr[110]));
			radix2 #(.width(width)) rd_st8_107  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[107]), .rdlo_in(a8_wr[111]),  .coef_in(coef[768]), .rdup_out(a9_wr[107]), .rdlo_out(a9_wr[111]));
			radix2 #(.width(width)) rd_st8_112  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[112]), .rdlo_in(a8_wr[116]),  .coef_in(coef[0]), .rdup_out(a9_wr[112]), .rdlo_out(a9_wr[116]));
			radix2 #(.width(width)) rd_st8_113  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[113]), .rdlo_in(a8_wr[117]),  .coef_in(coef[256]), .rdup_out(a9_wr[113]), .rdlo_out(a9_wr[117]));
			radix2 #(.width(width)) rd_st8_114  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[114]), .rdlo_in(a8_wr[118]),  .coef_in(coef[512]), .rdup_out(a9_wr[114]), .rdlo_out(a9_wr[118]));
			radix2 #(.width(width)) rd_st8_115  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[115]), .rdlo_in(a8_wr[119]),  .coef_in(coef[768]), .rdup_out(a9_wr[115]), .rdlo_out(a9_wr[119]));
			radix2 #(.width(width)) rd_st8_120  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[120]), .rdlo_in(a8_wr[124]),  .coef_in(coef[0]), .rdup_out(a9_wr[120]), .rdlo_out(a9_wr[124]));
			radix2 #(.width(width)) rd_st8_121  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[121]), .rdlo_in(a8_wr[125]),  .coef_in(coef[256]), .rdup_out(a9_wr[121]), .rdlo_out(a9_wr[125]));
			radix2 #(.width(width)) rd_st8_122  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[122]), .rdlo_in(a8_wr[126]),  .coef_in(coef[512]), .rdup_out(a9_wr[122]), .rdlo_out(a9_wr[126]));
			radix2 #(.width(width)) rd_st8_123  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[123]), .rdlo_in(a8_wr[127]),  .coef_in(coef[768]), .rdup_out(a9_wr[123]), .rdlo_out(a9_wr[127]));
			radix2 #(.width(width)) rd_st8_128  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[128]), .rdlo_in(a8_wr[132]),  .coef_in(coef[0]), .rdup_out(a9_wr[128]), .rdlo_out(a9_wr[132]));
			radix2 #(.width(width)) rd_st8_129  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[129]), .rdlo_in(a8_wr[133]),  .coef_in(coef[256]), .rdup_out(a9_wr[129]), .rdlo_out(a9_wr[133]));
			radix2 #(.width(width)) rd_st8_130  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[130]), .rdlo_in(a8_wr[134]),  .coef_in(coef[512]), .rdup_out(a9_wr[130]), .rdlo_out(a9_wr[134]));
			radix2 #(.width(width)) rd_st8_131  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[131]), .rdlo_in(a8_wr[135]),  .coef_in(coef[768]), .rdup_out(a9_wr[131]), .rdlo_out(a9_wr[135]));
			radix2 #(.width(width)) rd_st8_136  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[136]), .rdlo_in(a8_wr[140]),  .coef_in(coef[0]), .rdup_out(a9_wr[136]), .rdlo_out(a9_wr[140]));
			radix2 #(.width(width)) rd_st8_137  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[137]), .rdlo_in(a8_wr[141]),  .coef_in(coef[256]), .rdup_out(a9_wr[137]), .rdlo_out(a9_wr[141]));
			radix2 #(.width(width)) rd_st8_138  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[138]), .rdlo_in(a8_wr[142]),  .coef_in(coef[512]), .rdup_out(a9_wr[138]), .rdlo_out(a9_wr[142]));
			radix2 #(.width(width)) rd_st8_139  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[139]), .rdlo_in(a8_wr[143]),  .coef_in(coef[768]), .rdup_out(a9_wr[139]), .rdlo_out(a9_wr[143]));
			radix2 #(.width(width)) rd_st8_144  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[144]), .rdlo_in(a8_wr[148]),  .coef_in(coef[0]), .rdup_out(a9_wr[144]), .rdlo_out(a9_wr[148]));
			radix2 #(.width(width)) rd_st8_145  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[145]), .rdlo_in(a8_wr[149]),  .coef_in(coef[256]), .rdup_out(a9_wr[145]), .rdlo_out(a9_wr[149]));
			radix2 #(.width(width)) rd_st8_146  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[146]), .rdlo_in(a8_wr[150]),  .coef_in(coef[512]), .rdup_out(a9_wr[146]), .rdlo_out(a9_wr[150]));
			radix2 #(.width(width)) rd_st8_147  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[147]), .rdlo_in(a8_wr[151]),  .coef_in(coef[768]), .rdup_out(a9_wr[147]), .rdlo_out(a9_wr[151]));
			radix2 #(.width(width)) rd_st8_152  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[152]), .rdlo_in(a8_wr[156]),  .coef_in(coef[0]), .rdup_out(a9_wr[152]), .rdlo_out(a9_wr[156]));
			radix2 #(.width(width)) rd_st8_153  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[153]), .rdlo_in(a8_wr[157]),  .coef_in(coef[256]), .rdup_out(a9_wr[153]), .rdlo_out(a9_wr[157]));
			radix2 #(.width(width)) rd_st8_154  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[154]), .rdlo_in(a8_wr[158]),  .coef_in(coef[512]), .rdup_out(a9_wr[154]), .rdlo_out(a9_wr[158]));
			radix2 #(.width(width)) rd_st8_155  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[155]), .rdlo_in(a8_wr[159]),  .coef_in(coef[768]), .rdup_out(a9_wr[155]), .rdlo_out(a9_wr[159]));
			radix2 #(.width(width)) rd_st8_160  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[160]), .rdlo_in(a8_wr[164]),  .coef_in(coef[0]), .rdup_out(a9_wr[160]), .rdlo_out(a9_wr[164]));
			radix2 #(.width(width)) rd_st8_161  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[161]), .rdlo_in(a8_wr[165]),  .coef_in(coef[256]), .rdup_out(a9_wr[161]), .rdlo_out(a9_wr[165]));
			radix2 #(.width(width)) rd_st8_162  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[162]), .rdlo_in(a8_wr[166]),  .coef_in(coef[512]), .rdup_out(a9_wr[162]), .rdlo_out(a9_wr[166]));
			radix2 #(.width(width)) rd_st8_163  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[163]), .rdlo_in(a8_wr[167]),  .coef_in(coef[768]), .rdup_out(a9_wr[163]), .rdlo_out(a9_wr[167]));
			radix2 #(.width(width)) rd_st8_168  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[168]), .rdlo_in(a8_wr[172]),  .coef_in(coef[0]), .rdup_out(a9_wr[168]), .rdlo_out(a9_wr[172]));
			radix2 #(.width(width)) rd_st8_169  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[169]), .rdlo_in(a8_wr[173]),  .coef_in(coef[256]), .rdup_out(a9_wr[169]), .rdlo_out(a9_wr[173]));
			radix2 #(.width(width)) rd_st8_170  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[170]), .rdlo_in(a8_wr[174]),  .coef_in(coef[512]), .rdup_out(a9_wr[170]), .rdlo_out(a9_wr[174]));
			radix2 #(.width(width)) rd_st8_171  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[171]), .rdlo_in(a8_wr[175]),  .coef_in(coef[768]), .rdup_out(a9_wr[171]), .rdlo_out(a9_wr[175]));
			radix2 #(.width(width)) rd_st8_176  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[176]), .rdlo_in(a8_wr[180]),  .coef_in(coef[0]), .rdup_out(a9_wr[176]), .rdlo_out(a9_wr[180]));
			radix2 #(.width(width)) rd_st8_177  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[177]), .rdlo_in(a8_wr[181]),  .coef_in(coef[256]), .rdup_out(a9_wr[177]), .rdlo_out(a9_wr[181]));
			radix2 #(.width(width)) rd_st8_178  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[178]), .rdlo_in(a8_wr[182]),  .coef_in(coef[512]), .rdup_out(a9_wr[178]), .rdlo_out(a9_wr[182]));
			radix2 #(.width(width)) rd_st8_179  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[179]), .rdlo_in(a8_wr[183]),  .coef_in(coef[768]), .rdup_out(a9_wr[179]), .rdlo_out(a9_wr[183]));
			radix2 #(.width(width)) rd_st8_184  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[184]), .rdlo_in(a8_wr[188]),  .coef_in(coef[0]), .rdup_out(a9_wr[184]), .rdlo_out(a9_wr[188]));
			radix2 #(.width(width)) rd_st8_185  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[185]), .rdlo_in(a8_wr[189]),  .coef_in(coef[256]), .rdup_out(a9_wr[185]), .rdlo_out(a9_wr[189]));
			radix2 #(.width(width)) rd_st8_186  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[186]), .rdlo_in(a8_wr[190]),  .coef_in(coef[512]), .rdup_out(a9_wr[186]), .rdlo_out(a9_wr[190]));
			radix2 #(.width(width)) rd_st8_187  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[187]), .rdlo_in(a8_wr[191]),  .coef_in(coef[768]), .rdup_out(a9_wr[187]), .rdlo_out(a9_wr[191]));
			radix2 #(.width(width)) rd_st8_192  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[192]), .rdlo_in(a8_wr[196]),  .coef_in(coef[0]), .rdup_out(a9_wr[192]), .rdlo_out(a9_wr[196]));
			radix2 #(.width(width)) rd_st8_193  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[193]), .rdlo_in(a8_wr[197]),  .coef_in(coef[256]), .rdup_out(a9_wr[193]), .rdlo_out(a9_wr[197]));
			radix2 #(.width(width)) rd_st8_194  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[194]), .rdlo_in(a8_wr[198]),  .coef_in(coef[512]), .rdup_out(a9_wr[194]), .rdlo_out(a9_wr[198]));
			radix2 #(.width(width)) rd_st8_195  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[195]), .rdlo_in(a8_wr[199]),  .coef_in(coef[768]), .rdup_out(a9_wr[195]), .rdlo_out(a9_wr[199]));
			radix2 #(.width(width)) rd_st8_200  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[200]), .rdlo_in(a8_wr[204]),  .coef_in(coef[0]), .rdup_out(a9_wr[200]), .rdlo_out(a9_wr[204]));
			radix2 #(.width(width)) rd_st8_201  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[201]), .rdlo_in(a8_wr[205]),  .coef_in(coef[256]), .rdup_out(a9_wr[201]), .rdlo_out(a9_wr[205]));
			radix2 #(.width(width)) rd_st8_202  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[202]), .rdlo_in(a8_wr[206]),  .coef_in(coef[512]), .rdup_out(a9_wr[202]), .rdlo_out(a9_wr[206]));
			radix2 #(.width(width)) rd_st8_203  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[203]), .rdlo_in(a8_wr[207]),  .coef_in(coef[768]), .rdup_out(a9_wr[203]), .rdlo_out(a9_wr[207]));
			radix2 #(.width(width)) rd_st8_208  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[208]), .rdlo_in(a8_wr[212]),  .coef_in(coef[0]), .rdup_out(a9_wr[208]), .rdlo_out(a9_wr[212]));
			radix2 #(.width(width)) rd_st8_209  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[209]), .rdlo_in(a8_wr[213]),  .coef_in(coef[256]), .rdup_out(a9_wr[209]), .rdlo_out(a9_wr[213]));
			radix2 #(.width(width)) rd_st8_210  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[210]), .rdlo_in(a8_wr[214]),  .coef_in(coef[512]), .rdup_out(a9_wr[210]), .rdlo_out(a9_wr[214]));
			radix2 #(.width(width)) rd_st8_211  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[211]), .rdlo_in(a8_wr[215]),  .coef_in(coef[768]), .rdup_out(a9_wr[211]), .rdlo_out(a9_wr[215]));
			radix2 #(.width(width)) rd_st8_216  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[216]), .rdlo_in(a8_wr[220]),  .coef_in(coef[0]), .rdup_out(a9_wr[216]), .rdlo_out(a9_wr[220]));
			radix2 #(.width(width)) rd_st8_217  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[217]), .rdlo_in(a8_wr[221]),  .coef_in(coef[256]), .rdup_out(a9_wr[217]), .rdlo_out(a9_wr[221]));
			radix2 #(.width(width)) rd_st8_218  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[218]), .rdlo_in(a8_wr[222]),  .coef_in(coef[512]), .rdup_out(a9_wr[218]), .rdlo_out(a9_wr[222]));
			radix2 #(.width(width)) rd_st8_219  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[219]), .rdlo_in(a8_wr[223]),  .coef_in(coef[768]), .rdup_out(a9_wr[219]), .rdlo_out(a9_wr[223]));
			radix2 #(.width(width)) rd_st8_224  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[224]), .rdlo_in(a8_wr[228]),  .coef_in(coef[0]), .rdup_out(a9_wr[224]), .rdlo_out(a9_wr[228]));
			radix2 #(.width(width)) rd_st8_225  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[225]), .rdlo_in(a8_wr[229]),  .coef_in(coef[256]), .rdup_out(a9_wr[225]), .rdlo_out(a9_wr[229]));
			radix2 #(.width(width)) rd_st8_226  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[226]), .rdlo_in(a8_wr[230]),  .coef_in(coef[512]), .rdup_out(a9_wr[226]), .rdlo_out(a9_wr[230]));
			radix2 #(.width(width)) rd_st8_227  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[227]), .rdlo_in(a8_wr[231]),  .coef_in(coef[768]), .rdup_out(a9_wr[227]), .rdlo_out(a9_wr[231]));
			radix2 #(.width(width)) rd_st8_232  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[232]), .rdlo_in(a8_wr[236]),  .coef_in(coef[0]), .rdup_out(a9_wr[232]), .rdlo_out(a9_wr[236]));
			radix2 #(.width(width)) rd_st8_233  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[233]), .rdlo_in(a8_wr[237]),  .coef_in(coef[256]), .rdup_out(a9_wr[233]), .rdlo_out(a9_wr[237]));
			radix2 #(.width(width)) rd_st8_234  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[234]), .rdlo_in(a8_wr[238]),  .coef_in(coef[512]), .rdup_out(a9_wr[234]), .rdlo_out(a9_wr[238]));
			radix2 #(.width(width)) rd_st8_235  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[235]), .rdlo_in(a8_wr[239]),  .coef_in(coef[768]), .rdup_out(a9_wr[235]), .rdlo_out(a9_wr[239]));
			radix2 #(.width(width)) rd_st8_240  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[240]), .rdlo_in(a8_wr[244]),  .coef_in(coef[0]), .rdup_out(a9_wr[240]), .rdlo_out(a9_wr[244]));
			radix2 #(.width(width)) rd_st8_241  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[241]), .rdlo_in(a8_wr[245]),  .coef_in(coef[256]), .rdup_out(a9_wr[241]), .rdlo_out(a9_wr[245]));
			radix2 #(.width(width)) rd_st8_242  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[242]), .rdlo_in(a8_wr[246]),  .coef_in(coef[512]), .rdup_out(a9_wr[242]), .rdlo_out(a9_wr[246]));
			radix2 #(.width(width)) rd_st8_243  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[243]), .rdlo_in(a8_wr[247]),  .coef_in(coef[768]), .rdup_out(a9_wr[243]), .rdlo_out(a9_wr[247]));
			radix2 #(.width(width)) rd_st8_248  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[248]), .rdlo_in(a8_wr[252]),  .coef_in(coef[0]), .rdup_out(a9_wr[248]), .rdlo_out(a9_wr[252]));
			radix2 #(.width(width)) rd_st8_249  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[249]), .rdlo_in(a8_wr[253]),  .coef_in(coef[256]), .rdup_out(a9_wr[249]), .rdlo_out(a9_wr[253]));
			radix2 #(.width(width)) rd_st8_250  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[250]), .rdlo_in(a8_wr[254]),  .coef_in(coef[512]), .rdup_out(a9_wr[250]), .rdlo_out(a9_wr[254]));
			radix2 #(.width(width)) rd_st8_251  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[251]), .rdlo_in(a8_wr[255]),  .coef_in(coef[768]), .rdup_out(a9_wr[251]), .rdlo_out(a9_wr[255]));
			radix2 #(.width(width)) rd_st8_256  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[256]), .rdlo_in(a8_wr[260]),  .coef_in(coef[0]), .rdup_out(a9_wr[256]), .rdlo_out(a9_wr[260]));
			radix2 #(.width(width)) rd_st8_257  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[257]), .rdlo_in(a8_wr[261]),  .coef_in(coef[256]), .rdup_out(a9_wr[257]), .rdlo_out(a9_wr[261]));
			radix2 #(.width(width)) rd_st8_258  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[258]), .rdlo_in(a8_wr[262]),  .coef_in(coef[512]), .rdup_out(a9_wr[258]), .rdlo_out(a9_wr[262]));
			radix2 #(.width(width)) rd_st8_259  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[259]), .rdlo_in(a8_wr[263]),  .coef_in(coef[768]), .rdup_out(a9_wr[259]), .rdlo_out(a9_wr[263]));
			radix2 #(.width(width)) rd_st8_264  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[264]), .rdlo_in(a8_wr[268]),  .coef_in(coef[0]), .rdup_out(a9_wr[264]), .rdlo_out(a9_wr[268]));
			radix2 #(.width(width)) rd_st8_265  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[265]), .rdlo_in(a8_wr[269]),  .coef_in(coef[256]), .rdup_out(a9_wr[265]), .rdlo_out(a9_wr[269]));
			radix2 #(.width(width)) rd_st8_266  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[266]), .rdlo_in(a8_wr[270]),  .coef_in(coef[512]), .rdup_out(a9_wr[266]), .rdlo_out(a9_wr[270]));
			radix2 #(.width(width)) rd_st8_267  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[267]), .rdlo_in(a8_wr[271]),  .coef_in(coef[768]), .rdup_out(a9_wr[267]), .rdlo_out(a9_wr[271]));
			radix2 #(.width(width)) rd_st8_272  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[272]), .rdlo_in(a8_wr[276]),  .coef_in(coef[0]), .rdup_out(a9_wr[272]), .rdlo_out(a9_wr[276]));
			radix2 #(.width(width)) rd_st8_273  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[273]), .rdlo_in(a8_wr[277]),  .coef_in(coef[256]), .rdup_out(a9_wr[273]), .rdlo_out(a9_wr[277]));
			radix2 #(.width(width)) rd_st8_274  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[274]), .rdlo_in(a8_wr[278]),  .coef_in(coef[512]), .rdup_out(a9_wr[274]), .rdlo_out(a9_wr[278]));
			radix2 #(.width(width)) rd_st8_275  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[275]), .rdlo_in(a8_wr[279]),  .coef_in(coef[768]), .rdup_out(a9_wr[275]), .rdlo_out(a9_wr[279]));
			radix2 #(.width(width)) rd_st8_280  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[280]), .rdlo_in(a8_wr[284]),  .coef_in(coef[0]), .rdup_out(a9_wr[280]), .rdlo_out(a9_wr[284]));
			radix2 #(.width(width)) rd_st8_281  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[281]), .rdlo_in(a8_wr[285]),  .coef_in(coef[256]), .rdup_out(a9_wr[281]), .rdlo_out(a9_wr[285]));
			radix2 #(.width(width)) rd_st8_282  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[282]), .rdlo_in(a8_wr[286]),  .coef_in(coef[512]), .rdup_out(a9_wr[282]), .rdlo_out(a9_wr[286]));
			radix2 #(.width(width)) rd_st8_283  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[283]), .rdlo_in(a8_wr[287]),  .coef_in(coef[768]), .rdup_out(a9_wr[283]), .rdlo_out(a9_wr[287]));
			radix2 #(.width(width)) rd_st8_288  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[288]), .rdlo_in(a8_wr[292]),  .coef_in(coef[0]), .rdup_out(a9_wr[288]), .rdlo_out(a9_wr[292]));
			radix2 #(.width(width)) rd_st8_289  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[289]), .rdlo_in(a8_wr[293]),  .coef_in(coef[256]), .rdup_out(a9_wr[289]), .rdlo_out(a9_wr[293]));
			radix2 #(.width(width)) rd_st8_290  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[290]), .rdlo_in(a8_wr[294]),  .coef_in(coef[512]), .rdup_out(a9_wr[290]), .rdlo_out(a9_wr[294]));
			radix2 #(.width(width)) rd_st8_291  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[291]), .rdlo_in(a8_wr[295]),  .coef_in(coef[768]), .rdup_out(a9_wr[291]), .rdlo_out(a9_wr[295]));
			radix2 #(.width(width)) rd_st8_296  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[296]), .rdlo_in(a8_wr[300]),  .coef_in(coef[0]), .rdup_out(a9_wr[296]), .rdlo_out(a9_wr[300]));
			radix2 #(.width(width)) rd_st8_297  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[297]), .rdlo_in(a8_wr[301]),  .coef_in(coef[256]), .rdup_out(a9_wr[297]), .rdlo_out(a9_wr[301]));
			radix2 #(.width(width)) rd_st8_298  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[298]), .rdlo_in(a8_wr[302]),  .coef_in(coef[512]), .rdup_out(a9_wr[298]), .rdlo_out(a9_wr[302]));
			radix2 #(.width(width)) rd_st8_299  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[299]), .rdlo_in(a8_wr[303]),  .coef_in(coef[768]), .rdup_out(a9_wr[299]), .rdlo_out(a9_wr[303]));
			radix2 #(.width(width)) rd_st8_304  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[304]), .rdlo_in(a8_wr[308]),  .coef_in(coef[0]), .rdup_out(a9_wr[304]), .rdlo_out(a9_wr[308]));
			radix2 #(.width(width)) rd_st8_305  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[305]), .rdlo_in(a8_wr[309]),  .coef_in(coef[256]), .rdup_out(a9_wr[305]), .rdlo_out(a9_wr[309]));
			radix2 #(.width(width)) rd_st8_306  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[306]), .rdlo_in(a8_wr[310]),  .coef_in(coef[512]), .rdup_out(a9_wr[306]), .rdlo_out(a9_wr[310]));
			radix2 #(.width(width)) rd_st8_307  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[307]), .rdlo_in(a8_wr[311]),  .coef_in(coef[768]), .rdup_out(a9_wr[307]), .rdlo_out(a9_wr[311]));
			radix2 #(.width(width)) rd_st8_312  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[312]), .rdlo_in(a8_wr[316]),  .coef_in(coef[0]), .rdup_out(a9_wr[312]), .rdlo_out(a9_wr[316]));
			radix2 #(.width(width)) rd_st8_313  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[313]), .rdlo_in(a8_wr[317]),  .coef_in(coef[256]), .rdup_out(a9_wr[313]), .rdlo_out(a9_wr[317]));
			radix2 #(.width(width)) rd_st8_314  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[314]), .rdlo_in(a8_wr[318]),  .coef_in(coef[512]), .rdup_out(a9_wr[314]), .rdlo_out(a9_wr[318]));
			radix2 #(.width(width)) rd_st8_315  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[315]), .rdlo_in(a8_wr[319]),  .coef_in(coef[768]), .rdup_out(a9_wr[315]), .rdlo_out(a9_wr[319]));
			radix2 #(.width(width)) rd_st8_320  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[320]), .rdlo_in(a8_wr[324]),  .coef_in(coef[0]), .rdup_out(a9_wr[320]), .rdlo_out(a9_wr[324]));
			radix2 #(.width(width)) rd_st8_321  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[321]), .rdlo_in(a8_wr[325]),  .coef_in(coef[256]), .rdup_out(a9_wr[321]), .rdlo_out(a9_wr[325]));
			radix2 #(.width(width)) rd_st8_322  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[322]), .rdlo_in(a8_wr[326]),  .coef_in(coef[512]), .rdup_out(a9_wr[322]), .rdlo_out(a9_wr[326]));
			radix2 #(.width(width)) rd_st8_323  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[323]), .rdlo_in(a8_wr[327]),  .coef_in(coef[768]), .rdup_out(a9_wr[323]), .rdlo_out(a9_wr[327]));
			radix2 #(.width(width)) rd_st8_328  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[328]), .rdlo_in(a8_wr[332]),  .coef_in(coef[0]), .rdup_out(a9_wr[328]), .rdlo_out(a9_wr[332]));
			radix2 #(.width(width)) rd_st8_329  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[329]), .rdlo_in(a8_wr[333]),  .coef_in(coef[256]), .rdup_out(a9_wr[329]), .rdlo_out(a9_wr[333]));
			radix2 #(.width(width)) rd_st8_330  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[330]), .rdlo_in(a8_wr[334]),  .coef_in(coef[512]), .rdup_out(a9_wr[330]), .rdlo_out(a9_wr[334]));
			radix2 #(.width(width)) rd_st8_331  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[331]), .rdlo_in(a8_wr[335]),  .coef_in(coef[768]), .rdup_out(a9_wr[331]), .rdlo_out(a9_wr[335]));
			radix2 #(.width(width)) rd_st8_336  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[336]), .rdlo_in(a8_wr[340]),  .coef_in(coef[0]), .rdup_out(a9_wr[336]), .rdlo_out(a9_wr[340]));
			radix2 #(.width(width)) rd_st8_337  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[337]), .rdlo_in(a8_wr[341]),  .coef_in(coef[256]), .rdup_out(a9_wr[337]), .rdlo_out(a9_wr[341]));
			radix2 #(.width(width)) rd_st8_338  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[338]), .rdlo_in(a8_wr[342]),  .coef_in(coef[512]), .rdup_out(a9_wr[338]), .rdlo_out(a9_wr[342]));
			radix2 #(.width(width)) rd_st8_339  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[339]), .rdlo_in(a8_wr[343]),  .coef_in(coef[768]), .rdup_out(a9_wr[339]), .rdlo_out(a9_wr[343]));
			radix2 #(.width(width)) rd_st8_344  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[344]), .rdlo_in(a8_wr[348]),  .coef_in(coef[0]), .rdup_out(a9_wr[344]), .rdlo_out(a9_wr[348]));
			radix2 #(.width(width)) rd_st8_345  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[345]), .rdlo_in(a8_wr[349]),  .coef_in(coef[256]), .rdup_out(a9_wr[345]), .rdlo_out(a9_wr[349]));
			radix2 #(.width(width)) rd_st8_346  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[346]), .rdlo_in(a8_wr[350]),  .coef_in(coef[512]), .rdup_out(a9_wr[346]), .rdlo_out(a9_wr[350]));
			radix2 #(.width(width)) rd_st8_347  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[347]), .rdlo_in(a8_wr[351]),  .coef_in(coef[768]), .rdup_out(a9_wr[347]), .rdlo_out(a9_wr[351]));
			radix2 #(.width(width)) rd_st8_352  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[352]), .rdlo_in(a8_wr[356]),  .coef_in(coef[0]), .rdup_out(a9_wr[352]), .rdlo_out(a9_wr[356]));
			radix2 #(.width(width)) rd_st8_353  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[353]), .rdlo_in(a8_wr[357]),  .coef_in(coef[256]), .rdup_out(a9_wr[353]), .rdlo_out(a9_wr[357]));
			radix2 #(.width(width)) rd_st8_354  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[354]), .rdlo_in(a8_wr[358]),  .coef_in(coef[512]), .rdup_out(a9_wr[354]), .rdlo_out(a9_wr[358]));
			radix2 #(.width(width)) rd_st8_355  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[355]), .rdlo_in(a8_wr[359]),  .coef_in(coef[768]), .rdup_out(a9_wr[355]), .rdlo_out(a9_wr[359]));
			radix2 #(.width(width)) rd_st8_360  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[360]), .rdlo_in(a8_wr[364]),  .coef_in(coef[0]), .rdup_out(a9_wr[360]), .rdlo_out(a9_wr[364]));
			radix2 #(.width(width)) rd_st8_361  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[361]), .rdlo_in(a8_wr[365]),  .coef_in(coef[256]), .rdup_out(a9_wr[361]), .rdlo_out(a9_wr[365]));
			radix2 #(.width(width)) rd_st8_362  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[362]), .rdlo_in(a8_wr[366]),  .coef_in(coef[512]), .rdup_out(a9_wr[362]), .rdlo_out(a9_wr[366]));
			radix2 #(.width(width)) rd_st8_363  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[363]), .rdlo_in(a8_wr[367]),  .coef_in(coef[768]), .rdup_out(a9_wr[363]), .rdlo_out(a9_wr[367]));
			radix2 #(.width(width)) rd_st8_368  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[368]), .rdlo_in(a8_wr[372]),  .coef_in(coef[0]), .rdup_out(a9_wr[368]), .rdlo_out(a9_wr[372]));
			radix2 #(.width(width)) rd_st8_369  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[369]), .rdlo_in(a8_wr[373]),  .coef_in(coef[256]), .rdup_out(a9_wr[369]), .rdlo_out(a9_wr[373]));
			radix2 #(.width(width)) rd_st8_370  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[370]), .rdlo_in(a8_wr[374]),  .coef_in(coef[512]), .rdup_out(a9_wr[370]), .rdlo_out(a9_wr[374]));
			radix2 #(.width(width)) rd_st8_371  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[371]), .rdlo_in(a8_wr[375]),  .coef_in(coef[768]), .rdup_out(a9_wr[371]), .rdlo_out(a9_wr[375]));
			radix2 #(.width(width)) rd_st8_376  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[376]), .rdlo_in(a8_wr[380]),  .coef_in(coef[0]), .rdup_out(a9_wr[376]), .rdlo_out(a9_wr[380]));
			radix2 #(.width(width)) rd_st8_377  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[377]), .rdlo_in(a8_wr[381]),  .coef_in(coef[256]), .rdup_out(a9_wr[377]), .rdlo_out(a9_wr[381]));
			radix2 #(.width(width)) rd_st8_378  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[378]), .rdlo_in(a8_wr[382]),  .coef_in(coef[512]), .rdup_out(a9_wr[378]), .rdlo_out(a9_wr[382]));
			radix2 #(.width(width)) rd_st8_379  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[379]), .rdlo_in(a8_wr[383]),  .coef_in(coef[768]), .rdup_out(a9_wr[379]), .rdlo_out(a9_wr[383]));
			radix2 #(.width(width)) rd_st8_384  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[384]), .rdlo_in(a8_wr[388]),  .coef_in(coef[0]), .rdup_out(a9_wr[384]), .rdlo_out(a9_wr[388]));
			radix2 #(.width(width)) rd_st8_385  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[385]), .rdlo_in(a8_wr[389]),  .coef_in(coef[256]), .rdup_out(a9_wr[385]), .rdlo_out(a9_wr[389]));
			radix2 #(.width(width)) rd_st8_386  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[386]), .rdlo_in(a8_wr[390]),  .coef_in(coef[512]), .rdup_out(a9_wr[386]), .rdlo_out(a9_wr[390]));
			radix2 #(.width(width)) rd_st8_387  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[387]), .rdlo_in(a8_wr[391]),  .coef_in(coef[768]), .rdup_out(a9_wr[387]), .rdlo_out(a9_wr[391]));
			radix2 #(.width(width)) rd_st8_392  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[392]), .rdlo_in(a8_wr[396]),  .coef_in(coef[0]), .rdup_out(a9_wr[392]), .rdlo_out(a9_wr[396]));
			radix2 #(.width(width)) rd_st8_393  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[393]), .rdlo_in(a8_wr[397]),  .coef_in(coef[256]), .rdup_out(a9_wr[393]), .rdlo_out(a9_wr[397]));
			radix2 #(.width(width)) rd_st8_394  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[394]), .rdlo_in(a8_wr[398]),  .coef_in(coef[512]), .rdup_out(a9_wr[394]), .rdlo_out(a9_wr[398]));
			radix2 #(.width(width)) rd_st8_395  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[395]), .rdlo_in(a8_wr[399]),  .coef_in(coef[768]), .rdup_out(a9_wr[395]), .rdlo_out(a9_wr[399]));
			radix2 #(.width(width)) rd_st8_400  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[400]), .rdlo_in(a8_wr[404]),  .coef_in(coef[0]), .rdup_out(a9_wr[400]), .rdlo_out(a9_wr[404]));
			radix2 #(.width(width)) rd_st8_401  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[401]), .rdlo_in(a8_wr[405]),  .coef_in(coef[256]), .rdup_out(a9_wr[401]), .rdlo_out(a9_wr[405]));
			radix2 #(.width(width)) rd_st8_402  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[402]), .rdlo_in(a8_wr[406]),  .coef_in(coef[512]), .rdup_out(a9_wr[402]), .rdlo_out(a9_wr[406]));
			radix2 #(.width(width)) rd_st8_403  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[403]), .rdlo_in(a8_wr[407]),  .coef_in(coef[768]), .rdup_out(a9_wr[403]), .rdlo_out(a9_wr[407]));
			radix2 #(.width(width)) rd_st8_408  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[408]), .rdlo_in(a8_wr[412]),  .coef_in(coef[0]), .rdup_out(a9_wr[408]), .rdlo_out(a9_wr[412]));
			radix2 #(.width(width)) rd_st8_409  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[409]), .rdlo_in(a8_wr[413]),  .coef_in(coef[256]), .rdup_out(a9_wr[409]), .rdlo_out(a9_wr[413]));
			radix2 #(.width(width)) rd_st8_410  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[410]), .rdlo_in(a8_wr[414]),  .coef_in(coef[512]), .rdup_out(a9_wr[410]), .rdlo_out(a9_wr[414]));
			radix2 #(.width(width)) rd_st8_411  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[411]), .rdlo_in(a8_wr[415]),  .coef_in(coef[768]), .rdup_out(a9_wr[411]), .rdlo_out(a9_wr[415]));
			radix2 #(.width(width)) rd_st8_416  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[416]), .rdlo_in(a8_wr[420]),  .coef_in(coef[0]), .rdup_out(a9_wr[416]), .rdlo_out(a9_wr[420]));
			radix2 #(.width(width)) rd_st8_417  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[417]), .rdlo_in(a8_wr[421]),  .coef_in(coef[256]), .rdup_out(a9_wr[417]), .rdlo_out(a9_wr[421]));
			radix2 #(.width(width)) rd_st8_418  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[418]), .rdlo_in(a8_wr[422]),  .coef_in(coef[512]), .rdup_out(a9_wr[418]), .rdlo_out(a9_wr[422]));
			radix2 #(.width(width)) rd_st8_419  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[419]), .rdlo_in(a8_wr[423]),  .coef_in(coef[768]), .rdup_out(a9_wr[419]), .rdlo_out(a9_wr[423]));
			radix2 #(.width(width)) rd_st8_424  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[424]), .rdlo_in(a8_wr[428]),  .coef_in(coef[0]), .rdup_out(a9_wr[424]), .rdlo_out(a9_wr[428]));
			radix2 #(.width(width)) rd_st8_425  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[425]), .rdlo_in(a8_wr[429]),  .coef_in(coef[256]), .rdup_out(a9_wr[425]), .rdlo_out(a9_wr[429]));
			radix2 #(.width(width)) rd_st8_426  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[426]), .rdlo_in(a8_wr[430]),  .coef_in(coef[512]), .rdup_out(a9_wr[426]), .rdlo_out(a9_wr[430]));
			radix2 #(.width(width)) rd_st8_427  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[427]), .rdlo_in(a8_wr[431]),  .coef_in(coef[768]), .rdup_out(a9_wr[427]), .rdlo_out(a9_wr[431]));
			radix2 #(.width(width)) rd_st8_432  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[432]), .rdlo_in(a8_wr[436]),  .coef_in(coef[0]), .rdup_out(a9_wr[432]), .rdlo_out(a9_wr[436]));
			radix2 #(.width(width)) rd_st8_433  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[433]), .rdlo_in(a8_wr[437]),  .coef_in(coef[256]), .rdup_out(a9_wr[433]), .rdlo_out(a9_wr[437]));
			radix2 #(.width(width)) rd_st8_434  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[434]), .rdlo_in(a8_wr[438]),  .coef_in(coef[512]), .rdup_out(a9_wr[434]), .rdlo_out(a9_wr[438]));
			radix2 #(.width(width)) rd_st8_435  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[435]), .rdlo_in(a8_wr[439]),  .coef_in(coef[768]), .rdup_out(a9_wr[435]), .rdlo_out(a9_wr[439]));
			radix2 #(.width(width)) rd_st8_440  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[440]), .rdlo_in(a8_wr[444]),  .coef_in(coef[0]), .rdup_out(a9_wr[440]), .rdlo_out(a9_wr[444]));
			radix2 #(.width(width)) rd_st8_441  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[441]), .rdlo_in(a8_wr[445]),  .coef_in(coef[256]), .rdup_out(a9_wr[441]), .rdlo_out(a9_wr[445]));
			radix2 #(.width(width)) rd_st8_442  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[442]), .rdlo_in(a8_wr[446]),  .coef_in(coef[512]), .rdup_out(a9_wr[442]), .rdlo_out(a9_wr[446]));
			radix2 #(.width(width)) rd_st8_443  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[443]), .rdlo_in(a8_wr[447]),  .coef_in(coef[768]), .rdup_out(a9_wr[443]), .rdlo_out(a9_wr[447]));
			radix2 #(.width(width)) rd_st8_448  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[448]), .rdlo_in(a8_wr[452]),  .coef_in(coef[0]), .rdup_out(a9_wr[448]), .rdlo_out(a9_wr[452]));
			radix2 #(.width(width)) rd_st8_449  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[449]), .rdlo_in(a8_wr[453]),  .coef_in(coef[256]), .rdup_out(a9_wr[449]), .rdlo_out(a9_wr[453]));
			radix2 #(.width(width)) rd_st8_450  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[450]), .rdlo_in(a8_wr[454]),  .coef_in(coef[512]), .rdup_out(a9_wr[450]), .rdlo_out(a9_wr[454]));
			radix2 #(.width(width)) rd_st8_451  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[451]), .rdlo_in(a8_wr[455]),  .coef_in(coef[768]), .rdup_out(a9_wr[451]), .rdlo_out(a9_wr[455]));
			radix2 #(.width(width)) rd_st8_456  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[456]), .rdlo_in(a8_wr[460]),  .coef_in(coef[0]), .rdup_out(a9_wr[456]), .rdlo_out(a9_wr[460]));
			radix2 #(.width(width)) rd_st8_457  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[457]), .rdlo_in(a8_wr[461]),  .coef_in(coef[256]), .rdup_out(a9_wr[457]), .rdlo_out(a9_wr[461]));
			radix2 #(.width(width)) rd_st8_458  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[458]), .rdlo_in(a8_wr[462]),  .coef_in(coef[512]), .rdup_out(a9_wr[458]), .rdlo_out(a9_wr[462]));
			radix2 #(.width(width)) rd_st8_459  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[459]), .rdlo_in(a8_wr[463]),  .coef_in(coef[768]), .rdup_out(a9_wr[459]), .rdlo_out(a9_wr[463]));
			radix2 #(.width(width)) rd_st8_464  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[464]), .rdlo_in(a8_wr[468]),  .coef_in(coef[0]), .rdup_out(a9_wr[464]), .rdlo_out(a9_wr[468]));
			radix2 #(.width(width)) rd_st8_465  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[465]), .rdlo_in(a8_wr[469]),  .coef_in(coef[256]), .rdup_out(a9_wr[465]), .rdlo_out(a9_wr[469]));
			radix2 #(.width(width)) rd_st8_466  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[466]), .rdlo_in(a8_wr[470]),  .coef_in(coef[512]), .rdup_out(a9_wr[466]), .rdlo_out(a9_wr[470]));
			radix2 #(.width(width)) rd_st8_467  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[467]), .rdlo_in(a8_wr[471]),  .coef_in(coef[768]), .rdup_out(a9_wr[467]), .rdlo_out(a9_wr[471]));
			radix2 #(.width(width)) rd_st8_472  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[472]), .rdlo_in(a8_wr[476]),  .coef_in(coef[0]), .rdup_out(a9_wr[472]), .rdlo_out(a9_wr[476]));
			radix2 #(.width(width)) rd_st8_473  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[473]), .rdlo_in(a8_wr[477]),  .coef_in(coef[256]), .rdup_out(a9_wr[473]), .rdlo_out(a9_wr[477]));
			radix2 #(.width(width)) rd_st8_474  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[474]), .rdlo_in(a8_wr[478]),  .coef_in(coef[512]), .rdup_out(a9_wr[474]), .rdlo_out(a9_wr[478]));
			radix2 #(.width(width)) rd_st8_475  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[475]), .rdlo_in(a8_wr[479]),  .coef_in(coef[768]), .rdup_out(a9_wr[475]), .rdlo_out(a9_wr[479]));
			radix2 #(.width(width)) rd_st8_480  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[480]), .rdlo_in(a8_wr[484]),  .coef_in(coef[0]), .rdup_out(a9_wr[480]), .rdlo_out(a9_wr[484]));
			radix2 #(.width(width)) rd_st8_481  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[481]), .rdlo_in(a8_wr[485]),  .coef_in(coef[256]), .rdup_out(a9_wr[481]), .rdlo_out(a9_wr[485]));
			radix2 #(.width(width)) rd_st8_482  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[482]), .rdlo_in(a8_wr[486]),  .coef_in(coef[512]), .rdup_out(a9_wr[482]), .rdlo_out(a9_wr[486]));
			radix2 #(.width(width)) rd_st8_483  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[483]), .rdlo_in(a8_wr[487]),  .coef_in(coef[768]), .rdup_out(a9_wr[483]), .rdlo_out(a9_wr[487]));
			radix2 #(.width(width)) rd_st8_488  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[488]), .rdlo_in(a8_wr[492]),  .coef_in(coef[0]), .rdup_out(a9_wr[488]), .rdlo_out(a9_wr[492]));
			radix2 #(.width(width)) rd_st8_489  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[489]), .rdlo_in(a8_wr[493]),  .coef_in(coef[256]), .rdup_out(a9_wr[489]), .rdlo_out(a9_wr[493]));
			radix2 #(.width(width)) rd_st8_490  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[490]), .rdlo_in(a8_wr[494]),  .coef_in(coef[512]), .rdup_out(a9_wr[490]), .rdlo_out(a9_wr[494]));
			radix2 #(.width(width)) rd_st8_491  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[491]), .rdlo_in(a8_wr[495]),  .coef_in(coef[768]), .rdup_out(a9_wr[491]), .rdlo_out(a9_wr[495]));
			radix2 #(.width(width)) rd_st8_496  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[496]), .rdlo_in(a8_wr[500]),  .coef_in(coef[0]), .rdup_out(a9_wr[496]), .rdlo_out(a9_wr[500]));
			radix2 #(.width(width)) rd_st8_497  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[497]), .rdlo_in(a8_wr[501]),  .coef_in(coef[256]), .rdup_out(a9_wr[497]), .rdlo_out(a9_wr[501]));
			radix2 #(.width(width)) rd_st8_498  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[498]), .rdlo_in(a8_wr[502]),  .coef_in(coef[512]), .rdup_out(a9_wr[498]), .rdlo_out(a9_wr[502]));
			radix2 #(.width(width)) rd_st8_499  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[499]), .rdlo_in(a8_wr[503]),  .coef_in(coef[768]), .rdup_out(a9_wr[499]), .rdlo_out(a9_wr[503]));
			radix2 #(.width(width)) rd_st8_504  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[504]), .rdlo_in(a8_wr[508]),  .coef_in(coef[0]), .rdup_out(a9_wr[504]), .rdlo_out(a9_wr[508]));
			radix2 #(.width(width)) rd_st8_505  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[505]), .rdlo_in(a8_wr[509]),  .coef_in(coef[256]), .rdup_out(a9_wr[505]), .rdlo_out(a9_wr[509]));
			radix2 #(.width(width)) rd_st8_506  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[506]), .rdlo_in(a8_wr[510]),  .coef_in(coef[512]), .rdup_out(a9_wr[506]), .rdlo_out(a9_wr[510]));
			radix2 #(.width(width)) rd_st8_507  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[507]), .rdlo_in(a8_wr[511]),  .coef_in(coef[768]), .rdup_out(a9_wr[507]), .rdlo_out(a9_wr[511]));
			radix2 #(.width(width)) rd_st8_512  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[512]), .rdlo_in(a8_wr[516]),  .coef_in(coef[0]), .rdup_out(a9_wr[512]), .rdlo_out(a9_wr[516]));
			radix2 #(.width(width)) rd_st8_513  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[513]), .rdlo_in(a8_wr[517]),  .coef_in(coef[256]), .rdup_out(a9_wr[513]), .rdlo_out(a9_wr[517]));
			radix2 #(.width(width)) rd_st8_514  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[514]), .rdlo_in(a8_wr[518]),  .coef_in(coef[512]), .rdup_out(a9_wr[514]), .rdlo_out(a9_wr[518]));
			radix2 #(.width(width)) rd_st8_515  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[515]), .rdlo_in(a8_wr[519]),  .coef_in(coef[768]), .rdup_out(a9_wr[515]), .rdlo_out(a9_wr[519]));
			radix2 #(.width(width)) rd_st8_520  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[520]), .rdlo_in(a8_wr[524]),  .coef_in(coef[0]), .rdup_out(a9_wr[520]), .rdlo_out(a9_wr[524]));
			radix2 #(.width(width)) rd_st8_521  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[521]), .rdlo_in(a8_wr[525]),  .coef_in(coef[256]), .rdup_out(a9_wr[521]), .rdlo_out(a9_wr[525]));
			radix2 #(.width(width)) rd_st8_522  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[522]), .rdlo_in(a8_wr[526]),  .coef_in(coef[512]), .rdup_out(a9_wr[522]), .rdlo_out(a9_wr[526]));
			radix2 #(.width(width)) rd_st8_523  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[523]), .rdlo_in(a8_wr[527]),  .coef_in(coef[768]), .rdup_out(a9_wr[523]), .rdlo_out(a9_wr[527]));
			radix2 #(.width(width)) rd_st8_528  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[528]), .rdlo_in(a8_wr[532]),  .coef_in(coef[0]), .rdup_out(a9_wr[528]), .rdlo_out(a9_wr[532]));
			radix2 #(.width(width)) rd_st8_529  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[529]), .rdlo_in(a8_wr[533]),  .coef_in(coef[256]), .rdup_out(a9_wr[529]), .rdlo_out(a9_wr[533]));
			radix2 #(.width(width)) rd_st8_530  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[530]), .rdlo_in(a8_wr[534]),  .coef_in(coef[512]), .rdup_out(a9_wr[530]), .rdlo_out(a9_wr[534]));
			radix2 #(.width(width)) rd_st8_531  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[531]), .rdlo_in(a8_wr[535]),  .coef_in(coef[768]), .rdup_out(a9_wr[531]), .rdlo_out(a9_wr[535]));
			radix2 #(.width(width)) rd_st8_536  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[536]), .rdlo_in(a8_wr[540]),  .coef_in(coef[0]), .rdup_out(a9_wr[536]), .rdlo_out(a9_wr[540]));
			radix2 #(.width(width)) rd_st8_537  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[537]), .rdlo_in(a8_wr[541]),  .coef_in(coef[256]), .rdup_out(a9_wr[537]), .rdlo_out(a9_wr[541]));
			radix2 #(.width(width)) rd_st8_538  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[538]), .rdlo_in(a8_wr[542]),  .coef_in(coef[512]), .rdup_out(a9_wr[538]), .rdlo_out(a9_wr[542]));
			radix2 #(.width(width)) rd_st8_539  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[539]), .rdlo_in(a8_wr[543]),  .coef_in(coef[768]), .rdup_out(a9_wr[539]), .rdlo_out(a9_wr[543]));
			radix2 #(.width(width)) rd_st8_544  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[544]), .rdlo_in(a8_wr[548]),  .coef_in(coef[0]), .rdup_out(a9_wr[544]), .rdlo_out(a9_wr[548]));
			radix2 #(.width(width)) rd_st8_545  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[545]), .rdlo_in(a8_wr[549]),  .coef_in(coef[256]), .rdup_out(a9_wr[545]), .rdlo_out(a9_wr[549]));
			radix2 #(.width(width)) rd_st8_546  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[546]), .rdlo_in(a8_wr[550]),  .coef_in(coef[512]), .rdup_out(a9_wr[546]), .rdlo_out(a9_wr[550]));
			radix2 #(.width(width)) rd_st8_547  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[547]), .rdlo_in(a8_wr[551]),  .coef_in(coef[768]), .rdup_out(a9_wr[547]), .rdlo_out(a9_wr[551]));
			radix2 #(.width(width)) rd_st8_552  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[552]), .rdlo_in(a8_wr[556]),  .coef_in(coef[0]), .rdup_out(a9_wr[552]), .rdlo_out(a9_wr[556]));
			radix2 #(.width(width)) rd_st8_553  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[553]), .rdlo_in(a8_wr[557]),  .coef_in(coef[256]), .rdup_out(a9_wr[553]), .rdlo_out(a9_wr[557]));
			radix2 #(.width(width)) rd_st8_554  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[554]), .rdlo_in(a8_wr[558]),  .coef_in(coef[512]), .rdup_out(a9_wr[554]), .rdlo_out(a9_wr[558]));
			radix2 #(.width(width)) rd_st8_555  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[555]), .rdlo_in(a8_wr[559]),  .coef_in(coef[768]), .rdup_out(a9_wr[555]), .rdlo_out(a9_wr[559]));
			radix2 #(.width(width)) rd_st8_560  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[560]), .rdlo_in(a8_wr[564]),  .coef_in(coef[0]), .rdup_out(a9_wr[560]), .rdlo_out(a9_wr[564]));
			radix2 #(.width(width)) rd_st8_561  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[561]), .rdlo_in(a8_wr[565]),  .coef_in(coef[256]), .rdup_out(a9_wr[561]), .rdlo_out(a9_wr[565]));
			radix2 #(.width(width)) rd_st8_562  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[562]), .rdlo_in(a8_wr[566]),  .coef_in(coef[512]), .rdup_out(a9_wr[562]), .rdlo_out(a9_wr[566]));
			radix2 #(.width(width)) rd_st8_563  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[563]), .rdlo_in(a8_wr[567]),  .coef_in(coef[768]), .rdup_out(a9_wr[563]), .rdlo_out(a9_wr[567]));
			radix2 #(.width(width)) rd_st8_568  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[568]), .rdlo_in(a8_wr[572]),  .coef_in(coef[0]), .rdup_out(a9_wr[568]), .rdlo_out(a9_wr[572]));
			radix2 #(.width(width)) rd_st8_569  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[569]), .rdlo_in(a8_wr[573]),  .coef_in(coef[256]), .rdup_out(a9_wr[569]), .rdlo_out(a9_wr[573]));
			radix2 #(.width(width)) rd_st8_570  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[570]), .rdlo_in(a8_wr[574]),  .coef_in(coef[512]), .rdup_out(a9_wr[570]), .rdlo_out(a9_wr[574]));
			radix2 #(.width(width)) rd_st8_571  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[571]), .rdlo_in(a8_wr[575]),  .coef_in(coef[768]), .rdup_out(a9_wr[571]), .rdlo_out(a9_wr[575]));
			radix2 #(.width(width)) rd_st8_576  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[576]), .rdlo_in(a8_wr[580]),  .coef_in(coef[0]), .rdup_out(a9_wr[576]), .rdlo_out(a9_wr[580]));
			radix2 #(.width(width)) rd_st8_577  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[577]), .rdlo_in(a8_wr[581]),  .coef_in(coef[256]), .rdup_out(a9_wr[577]), .rdlo_out(a9_wr[581]));
			radix2 #(.width(width)) rd_st8_578  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[578]), .rdlo_in(a8_wr[582]),  .coef_in(coef[512]), .rdup_out(a9_wr[578]), .rdlo_out(a9_wr[582]));
			radix2 #(.width(width)) rd_st8_579  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[579]), .rdlo_in(a8_wr[583]),  .coef_in(coef[768]), .rdup_out(a9_wr[579]), .rdlo_out(a9_wr[583]));
			radix2 #(.width(width)) rd_st8_584  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[584]), .rdlo_in(a8_wr[588]),  .coef_in(coef[0]), .rdup_out(a9_wr[584]), .rdlo_out(a9_wr[588]));
			radix2 #(.width(width)) rd_st8_585  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[585]), .rdlo_in(a8_wr[589]),  .coef_in(coef[256]), .rdup_out(a9_wr[585]), .rdlo_out(a9_wr[589]));
			radix2 #(.width(width)) rd_st8_586  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[586]), .rdlo_in(a8_wr[590]),  .coef_in(coef[512]), .rdup_out(a9_wr[586]), .rdlo_out(a9_wr[590]));
			radix2 #(.width(width)) rd_st8_587  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[587]), .rdlo_in(a8_wr[591]),  .coef_in(coef[768]), .rdup_out(a9_wr[587]), .rdlo_out(a9_wr[591]));
			radix2 #(.width(width)) rd_st8_592  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[592]), .rdlo_in(a8_wr[596]),  .coef_in(coef[0]), .rdup_out(a9_wr[592]), .rdlo_out(a9_wr[596]));
			radix2 #(.width(width)) rd_st8_593  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[593]), .rdlo_in(a8_wr[597]),  .coef_in(coef[256]), .rdup_out(a9_wr[593]), .rdlo_out(a9_wr[597]));
			radix2 #(.width(width)) rd_st8_594  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[594]), .rdlo_in(a8_wr[598]),  .coef_in(coef[512]), .rdup_out(a9_wr[594]), .rdlo_out(a9_wr[598]));
			radix2 #(.width(width)) rd_st8_595  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[595]), .rdlo_in(a8_wr[599]),  .coef_in(coef[768]), .rdup_out(a9_wr[595]), .rdlo_out(a9_wr[599]));
			radix2 #(.width(width)) rd_st8_600  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[600]), .rdlo_in(a8_wr[604]),  .coef_in(coef[0]), .rdup_out(a9_wr[600]), .rdlo_out(a9_wr[604]));
			radix2 #(.width(width)) rd_st8_601  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[601]), .rdlo_in(a8_wr[605]),  .coef_in(coef[256]), .rdup_out(a9_wr[601]), .rdlo_out(a9_wr[605]));
			radix2 #(.width(width)) rd_st8_602  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[602]), .rdlo_in(a8_wr[606]),  .coef_in(coef[512]), .rdup_out(a9_wr[602]), .rdlo_out(a9_wr[606]));
			radix2 #(.width(width)) rd_st8_603  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[603]), .rdlo_in(a8_wr[607]),  .coef_in(coef[768]), .rdup_out(a9_wr[603]), .rdlo_out(a9_wr[607]));
			radix2 #(.width(width)) rd_st8_608  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[608]), .rdlo_in(a8_wr[612]),  .coef_in(coef[0]), .rdup_out(a9_wr[608]), .rdlo_out(a9_wr[612]));
			radix2 #(.width(width)) rd_st8_609  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[609]), .rdlo_in(a8_wr[613]),  .coef_in(coef[256]), .rdup_out(a9_wr[609]), .rdlo_out(a9_wr[613]));
			radix2 #(.width(width)) rd_st8_610  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[610]), .rdlo_in(a8_wr[614]),  .coef_in(coef[512]), .rdup_out(a9_wr[610]), .rdlo_out(a9_wr[614]));
			radix2 #(.width(width)) rd_st8_611  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[611]), .rdlo_in(a8_wr[615]),  .coef_in(coef[768]), .rdup_out(a9_wr[611]), .rdlo_out(a9_wr[615]));
			radix2 #(.width(width)) rd_st8_616  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[616]), .rdlo_in(a8_wr[620]),  .coef_in(coef[0]), .rdup_out(a9_wr[616]), .rdlo_out(a9_wr[620]));
			radix2 #(.width(width)) rd_st8_617  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[617]), .rdlo_in(a8_wr[621]),  .coef_in(coef[256]), .rdup_out(a9_wr[617]), .rdlo_out(a9_wr[621]));
			radix2 #(.width(width)) rd_st8_618  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[618]), .rdlo_in(a8_wr[622]),  .coef_in(coef[512]), .rdup_out(a9_wr[618]), .rdlo_out(a9_wr[622]));
			radix2 #(.width(width)) rd_st8_619  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[619]), .rdlo_in(a8_wr[623]),  .coef_in(coef[768]), .rdup_out(a9_wr[619]), .rdlo_out(a9_wr[623]));
			radix2 #(.width(width)) rd_st8_624  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[624]), .rdlo_in(a8_wr[628]),  .coef_in(coef[0]), .rdup_out(a9_wr[624]), .rdlo_out(a9_wr[628]));
			radix2 #(.width(width)) rd_st8_625  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[625]), .rdlo_in(a8_wr[629]),  .coef_in(coef[256]), .rdup_out(a9_wr[625]), .rdlo_out(a9_wr[629]));
			radix2 #(.width(width)) rd_st8_626  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[626]), .rdlo_in(a8_wr[630]),  .coef_in(coef[512]), .rdup_out(a9_wr[626]), .rdlo_out(a9_wr[630]));
			radix2 #(.width(width)) rd_st8_627  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[627]), .rdlo_in(a8_wr[631]),  .coef_in(coef[768]), .rdup_out(a9_wr[627]), .rdlo_out(a9_wr[631]));
			radix2 #(.width(width)) rd_st8_632  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[632]), .rdlo_in(a8_wr[636]),  .coef_in(coef[0]), .rdup_out(a9_wr[632]), .rdlo_out(a9_wr[636]));
			radix2 #(.width(width)) rd_st8_633  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[633]), .rdlo_in(a8_wr[637]),  .coef_in(coef[256]), .rdup_out(a9_wr[633]), .rdlo_out(a9_wr[637]));
			radix2 #(.width(width)) rd_st8_634  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[634]), .rdlo_in(a8_wr[638]),  .coef_in(coef[512]), .rdup_out(a9_wr[634]), .rdlo_out(a9_wr[638]));
			radix2 #(.width(width)) rd_st8_635  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[635]), .rdlo_in(a8_wr[639]),  .coef_in(coef[768]), .rdup_out(a9_wr[635]), .rdlo_out(a9_wr[639]));
			radix2 #(.width(width)) rd_st8_640  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[640]), .rdlo_in(a8_wr[644]),  .coef_in(coef[0]), .rdup_out(a9_wr[640]), .rdlo_out(a9_wr[644]));
			radix2 #(.width(width)) rd_st8_641  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[641]), .rdlo_in(a8_wr[645]),  .coef_in(coef[256]), .rdup_out(a9_wr[641]), .rdlo_out(a9_wr[645]));
			radix2 #(.width(width)) rd_st8_642  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[642]), .rdlo_in(a8_wr[646]),  .coef_in(coef[512]), .rdup_out(a9_wr[642]), .rdlo_out(a9_wr[646]));
			radix2 #(.width(width)) rd_st8_643  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[643]), .rdlo_in(a8_wr[647]),  .coef_in(coef[768]), .rdup_out(a9_wr[643]), .rdlo_out(a9_wr[647]));
			radix2 #(.width(width)) rd_st8_648  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[648]), .rdlo_in(a8_wr[652]),  .coef_in(coef[0]), .rdup_out(a9_wr[648]), .rdlo_out(a9_wr[652]));
			radix2 #(.width(width)) rd_st8_649  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[649]), .rdlo_in(a8_wr[653]),  .coef_in(coef[256]), .rdup_out(a9_wr[649]), .rdlo_out(a9_wr[653]));
			radix2 #(.width(width)) rd_st8_650  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[650]), .rdlo_in(a8_wr[654]),  .coef_in(coef[512]), .rdup_out(a9_wr[650]), .rdlo_out(a9_wr[654]));
			radix2 #(.width(width)) rd_st8_651  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[651]), .rdlo_in(a8_wr[655]),  .coef_in(coef[768]), .rdup_out(a9_wr[651]), .rdlo_out(a9_wr[655]));
			radix2 #(.width(width)) rd_st8_656  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[656]), .rdlo_in(a8_wr[660]),  .coef_in(coef[0]), .rdup_out(a9_wr[656]), .rdlo_out(a9_wr[660]));
			radix2 #(.width(width)) rd_st8_657  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[657]), .rdlo_in(a8_wr[661]),  .coef_in(coef[256]), .rdup_out(a9_wr[657]), .rdlo_out(a9_wr[661]));
			radix2 #(.width(width)) rd_st8_658  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[658]), .rdlo_in(a8_wr[662]),  .coef_in(coef[512]), .rdup_out(a9_wr[658]), .rdlo_out(a9_wr[662]));
			radix2 #(.width(width)) rd_st8_659  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[659]), .rdlo_in(a8_wr[663]),  .coef_in(coef[768]), .rdup_out(a9_wr[659]), .rdlo_out(a9_wr[663]));
			radix2 #(.width(width)) rd_st8_664  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[664]), .rdlo_in(a8_wr[668]),  .coef_in(coef[0]), .rdup_out(a9_wr[664]), .rdlo_out(a9_wr[668]));
			radix2 #(.width(width)) rd_st8_665  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[665]), .rdlo_in(a8_wr[669]),  .coef_in(coef[256]), .rdup_out(a9_wr[665]), .rdlo_out(a9_wr[669]));
			radix2 #(.width(width)) rd_st8_666  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[666]), .rdlo_in(a8_wr[670]),  .coef_in(coef[512]), .rdup_out(a9_wr[666]), .rdlo_out(a9_wr[670]));
			radix2 #(.width(width)) rd_st8_667  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[667]), .rdlo_in(a8_wr[671]),  .coef_in(coef[768]), .rdup_out(a9_wr[667]), .rdlo_out(a9_wr[671]));
			radix2 #(.width(width)) rd_st8_672  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[672]), .rdlo_in(a8_wr[676]),  .coef_in(coef[0]), .rdup_out(a9_wr[672]), .rdlo_out(a9_wr[676]));
			radix2 #(.width(width)) rd_st8_673  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[673]), .rdlo_in(a8_wr[677]),  .coef_in(coef[256]), .rdup_out(a9_wr[673]), .rdlo_out(a9_wr[677]));
			radix2 #(.width(width)) rd_st8_674  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[674]), .rdlo_in(a8_wr[678]),  .coef_in(coef[512]), .rdup_out(a9_wr[674]), .rdlo_out(a9_wr[678]));
			radix2 #(.width(width)) rd_st8_675  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[675]), .rdlo_in(a8_wr[679]),  .coef_in(coef[768]), .rdup_out(a9_wr[675]), .rdlo_out(a9_wr[679]));
			radix2 #(.width(width)) rd_st8_680  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[680]), .rdlo_in(a8_wr[684]),  .coef_in(coef[0]), .rdup_out(a9_wr[680]), .rdlo_out(a9_wr[684]));
			radix2 #(.width(width)) rd_st8_681  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[681]), .rdlo_in(a8_wr[685]),  .coef_in(coef[256]), .rdup_out(a9_wr[681]), .rdlo_out(a9_wr[685]));
			radix2 #(.width(width)) rd_st8_682  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[682]), .rdlo_in(a8_wr[686]),  .coef_in(coef[512]), .rdup_out(a9_wr[682]), .rdlo_out(a9_wr[686]));
			radix2 #(.width(width)) rd_st8_683  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[683]), .rdlo_in(a8_wr[687]),  .coef_in(coef[768]), .rdup_out(a9_wr[683]), .rdlo_out(a9_wr[687]));
			radix2 #(.width(width)) rd_st8_688  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[688]), .rdlo_in(a8_wr[692]),  .coef_in(coef[0]), .rdup_out(a9_wr[688]), .rdlo_out(a9_wr[692]));
			radix2 #(.width(width)) rd_st8_689  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[689]), .rdlo_in(a8_wr[693]),  .coef_in(coef[256]), .rdup_out(a9_wr[689]), .rdlo_out(a9_wr[693]));
			radix2 #(.width(width)) rd_st8_690  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[690]), .rdlo_in(a8_wr[694]),  .coef_in(coef[512]), .rdup_out(a9_wr[690]), .rdlo_out(a9_wr[694]));
			radix2 #(.width(width)) rd_st8_691  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[691]), .rdlo_in(a8_wr[695]),  .coef_in(coef[768]), .rdup_out(a9_wr[691]), .rdlo_out(a9_wr[695]));
			radix2 #(.width(width)) rd_st8_696  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[696]), .rdlo_in(a8_wr[700]),  .coef_in(coef[0]), .rdup_out(a9_wr[696]), .rdlo_out(a9_wr[700]));
			radix2 #(.width(width)) rd_st8_697  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[697]), .rdlo_in(a8_wr[701]),  .coef_in(coef[256]), .rdup_out(a9_wr[697]), .rdlo_out(a9_wr[701]));
			radix2 #(.width(width)) rd_st8_698  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[698]), .rdlo_in(a8_wr[702]),  .coef_in(coef[512]), .rdup_out(a9_wr[698]), .rdlo_out(a9_wr[702]));
			radix2 #(.width(width)) rd_st8_699  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[699]), .rdlo_in(a8_wr[703]),  .coef_in(coef[768]), .rdup_out(a9_wr[699]), .rdlo_out(a9_wr[703]));
			radix2 #(.width(width)) rd_st8_704  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[704]), .rdlo_in(a8_wr[708]),  .coef_in(coef[0]), .rdup_out(a9_wr[704]), .rdlo_out(a9_wr[708]));
			radix2 #(.width(width)) rd_st8_705  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[705]), .rdlo_in(a8_wr[709]),  .coef_in(coef[256]), .rdup_out(a9_wr[705]), .rdlo_out(a9_wr[709]));
			radix2 #(.width(width)) rd_st8_706  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[706]), .rdlo_in(a8_wr[710]),  .coef_in(coef[512]), .rdup_out(a9_wr[706]), .rdlo_out(a9_wr[710]));
			radix2 #(.width(width)) rd_st8_707  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[707]), .rdlo_in(a8_wr[711]),  .coef_in(coef[768]), .rdup_out(a9_wr[707]), .rdlo_out(a9_wr[711]));
			radix2 #(.width(width)) rd_st8_712  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[712]), .rdlo_in(a8_wr[716]),  .coef_in(coef[0]), .rdup_out(a9_wr[712]), .rdlo_out(a9_wr[716]));
			radix2 #(.width(width)) rd_st8_713  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[713]), .rdlo_in(a8_wr[717]),  .coef_in(coef[256]), .rdup_out(a9_wr[713]), .rdlo_out(a9_wr[717]));
			radix2 #(.width(width)) rd_st8_714  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[714]), .rdlo_in(a8_wr[718]),  .coef_in(coef[512]), .rdup_out(a9_wr[714]), .rdlo_out(a9_wr[718]));
			radix2 #(.width(width)) rd_st8_715  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[715]), .rdlo_in(a8_wr[719]),  .coef_in(coef[768]), .rdup_out(a9_wr[715]), .rdlo_out(a9_wr[719]));
			radix2 #(.width(width)) rd_st8_720  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[720]), .rdlo_in(a8_wr[724]),  .coef_in(coef[0]), .rdup_out(a9_wr[720]), .rdlo_out(a9_wr[724]));
			radix2 #(.width(width)) rd_st8_721  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[721]), .rdlo_in(a8_wr[725]),  .coef_in(coef[256]), .rdup_out(a9_wr[721]), .rdlo_out(a9_wr[725]));
			radix2 #(.width(width)) rd_st8_722  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[722]), .rdlo_in(a8_wr[726]),  .coef_in(coef[512]), .rdup_out(a9_wr[722]), .rdlo_out(a9_wr[726]));
			radix2 #(.width(width)) rd_st8_723  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[723]), .rdlo_in(a8_wr[727]),  .coef_in(coef[768]), .rdup_out(a9_wr[723]), .rdlo_out(a9_wr[727]));
			radix2 #(.width(width)) rd_st8_728  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[728]), .rdlo_in(a8_wr[732]),  .coef_in(coef[0]), .rdup_out(a9_wr[728]), .rdlo_out(a9_wr[732]));
			radix2 #(.width(width)) rd_st8_729  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[729]), .rdlo_in(a8_wr[733]),  .coef_in(coef[256]), .rdup_out(a9_wr[729]), .rdlo_out(a9_wr[733]));
			radix2 #(.width(width)) rd_st8_730  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[730]), .rdlo_in(a8_wr[734]),  .coef_in(coef[512]), .rdup_out(a9_wr[730]), .rdlo_out(a9_wr[734]));
			radix2 #(.width(width)) rd_st8_731  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[731]), .rdlo_in(a8_wr[735]),  .coef_in(coef[768]), .rdup_out(a9_wr[731]), .rdlo_out(a9_wr[735]));
			radix2 #(.width(width)) rd_st8_736  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[736]), .rdlo_in(a8_wr[740]),  .coef_in(coef[0]), .rdup_out(a9_wr[736]), .rdlo_out(a9_wr[740]));
			radix2 #(.width(width)) rd_st8_737  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[737]), .rdlo_in(a8_wr[741]),  .coef_in(coef[256]), .rdup_out(a9_wr[737]), .rdlo_out(a9_wr[741]));
			radix2 #(.width(width)) rd_st8_738  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[738]), .rdlo_in(a8_wr[742]),  .coef_in(coef[512]), .rdup_out(a9_wr[738]), .rdlo_out(a9_wr[742]));
			radix2 #(.width(width)) rd_st8_739  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[739]), .rdlo_in(a8_wr[743]),  .coef_in(coef[768]), .rdup_out(a9_wr[739]), .rdlo_out(a9_wr[743]));
			radix2 #(.width(width)) rd_st8_744  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[744]), .rdlo_in(a8_wr[748]),  .coef_in(coef[0]), .rdup_out(a9_wr[744]), .rdlo_out(a9_wr[748]));
			radix2 #(.width(width)) rd_st8_745  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[745]), .rdlo_in(a8_wr[749]),  .coef_in(coef[256]), .rdup_out(a9_wr[745]), .rdlo_out(a9_wr[749]));
			radix2 #(.width(width)) rd_st8_746  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[746]), .rdlo_in(a8_wr[750]),  .coef_in(coef[512]), .rdup_out(a9_wr[746]), .rdlo_out(a9_wr[750]));
			radix2 #(.width(width)) rd_st8_747  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[747]), .rdlo_in(a8_wr[751]),  .coef_in(coef[768]), .rdup_out(a9_wr[747]), .rdlo_out(a9_wr[751]));
			radix2 #(.width(width)) rd_st8_752  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[752]), .rdlo_in(a8_wr[756]),  .coef_in(coef[0]), .rdup_out(a9_wr[752]), .rdlo_out(a9_wr[756]));
			radix2 #(.width(width)) rd_st8_753  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[753]), .rdlo_in(a8_wr[757]),  .coef_in(coef[256]), .rdup_out(a9_wr[753]), .rdlo_out(a9_wr[757]));
			radix2 #(.width(width)) rd_st8_754  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[754]), .rdlo_in(a8_wr[758]),  .coef_in(coef[512]), .rdup_out(a9_wr[754]), .rdlo_out(a9_wr[758]));
			radix2 #(.width(width)) rd_st8_755  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[755]), .rdlo_in(a8_wr[759]),  .coef_in(coef[768]), .rdup_out(a9_wr[755]), .rdlo_out(a9_wr[759]));
			radix2 #(.width(width)) rd_st8_760  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[760]), .rdlo_in(a8_wr[764]),  .coef_in(coef[0]), .rdup_out(a9_wr[760]), .rdlo_out(a9_wr[764]));
			radix2 #(.width(width)) rd_st8_761  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[761]), .rdlo_in(a8_wr[765]),  .coef_in(coef[256]), .rdup_out(a9_wr[761]), .rdlo_out(a9_wr[765]));
			radix2 #(.width(width)) rd_st8_762  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[762]), .rdlo_in(a8_wr[766]),  .coef_in(coef[512]), .rdup_out(a9_wr[762]), .rdlo_out(a9_wr[766]));
			radix2 #(.width(width)) rd_st8_763  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[763]), .rdlo_in(a8_wr[767]),  .coef_in(coef[768]), .rdup_out(a9_wr[763]), .rdlo_out(a9_wr[767]));
			radix2 #(.width(width)) rd_st8_768  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[768]), .rdlo_in(a8_wr[772]),  .coef_in(coef[0]), .rdup_out(a9_wr[768]), .rdlo_out(a9_wr[772]));
			radix2 #(.width(width)) rd_st8_769  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[769]), .rdlo_in(a8_wr[773]),  .coef_in(coef[256]), .rdup_out(a9_wr[769]), .rdlo_out(a9_wr[773]));
			radix2 #(.width(width)) rd_st8_770  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[770]), .rdlo_in(a8_wr[774]),  .coef_in(coef[512]), .rdup_out(a9_wr[770]), .rdlo_out(a9_wr[774]));
			radix2 #(.width(width)) rd_st8_771  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[771]), .rdlo_in(a8_wr[775]),  .coef_in(coef[768]), .rdup_out(a9_wr[771]), .rdlo_out(a9_wr[775]));
			radix2 #(.width(width)) rd_st8_776  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[776]), .rdlo_in(a8_wr[780]),  .coef_in(coef[0]), .rdup_out(a9_wr[776]), .rdlo_out(a9_wr[780]));
			radix2 #(.width(width)) rd_st8_777  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[777]), .rdlo_in(a8_wr[781]),  .coef_in(coef[256]), .rdup_out(a9_wr[777]), .rdlo_out(a9_wr[781]));
			radix2 #(.width(width)) rd_st8_778  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[778]), .rdlo_in(a8_wr[782]),  .coef_in(coef[512]), .rdup_out(a9_wr[778]), .rdlo_out(a9_wr[782]));
			radix2 #(.width(width)) rd_st8_779  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[779]), .rdlo_in(a8_wr[783]),  .coef_in(coef[768]), .rdup_out(a9_wr[779]), .rdlo_out(a9_wr[783]));
			radix2 #(.width(width)) rd_st8_784  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[784]), .rdlo_in(a8_wr[788]),  .coef_in(coef[0]), .rdup_out(a9_wr[784]), .rdlo_out(a9_wr[788]));
			radix2 #(.width(width)) rd_st8_785  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[785]), .rdlo_in(a8_wr[789]),  .coef_in(coef[256]), .rdup_out(a9_wr[785]), .rdlo_out(a9_wr[789]));
			radix2 #(.width(width)) rd_st8_786  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[786]), .rdlo_in(a8_wr[790]),  .coef_in(coef[512]), .rdup_out(a9_wr[786]), .rdlo_out(a9_wr[790]));
			radix2 #(.width(width)) rd_st8_787  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[787]), .rdlo_in(a8_wr[791]),  .coef_in(coef[768]), .rdup_out(a9_wr[787]), .rdlo_out(a9_wr[791]));
			radix2 #(.width(width)) rd_st8_792  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[792]), .rdlo_in(a8_wr[796]),  .coef_in(coef[0]), .rdup_out(a9_wr[792]), .rdlo_out(a9_wr[796]));
			radix2 #(.width(width)) rd_st8_793  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[793]), .rdlo_in(a8_wr[797]),  .coef_in(coef[256]), .rdup_out(a9_wr[793]), .rdlo_out(a9_wr[797]));
			radix2 #(.width(width)) rd_st8_794  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[794]), .rdlo_in(a8_wr[798]),  .coef_in(coef[512]), .rdup_out(a9_wr[794]), .rdlo_out(a9_wr[798]));
			radix2 #(.width(width)) rd_st8_795  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[795]), .rdlo_in(a8_wr[799]),  .coef_in(coef[768]), .rdup_out(a9_wr[795]), .rdlo_out(a9_wr[799]));
			radix2 #(.width(width)) rd_st8_800  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[800]), .rdlo_in(a8_wr[804]),  .coef_in(coef[0]), .rdup_out(a9_wr[800]), .rdlo_out(a9_wr[804]));
			radix2 #(.width(width)) rd_st8_801  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[801]), .rdlo_in(a8_wr[805]),  .coef_in(coef[256]), .rdup_out(a9_wr[801]), .rdlo_out(a9_wr[805]));
			radix2 #(.width(width)) rd_st8_802  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[802]), .rdlo_in(a8_wr[806]),  .coef_in(coef[512]), .rdup_out(a9_wr[802]), .rdlo_out(a9_wr[806]));
			radix2 #(.width(width)) rd_st8_803  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[803]), .rdlo_in(a8_wr[807]),  .coef_in(coef[768]), .rdup_out(a9_wr[803]), .rdlo_out(a9_wr[807]));
			radix2 #(.width(width)) rd_st8_808  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[808]), .rdlo_in(a8_wr[812]),  .coef_in(coef[0]), .rdup_out(a9_wr[808]), .rdlo_out(a9_wr[812]));
			radix2 #(.width(width)) rd_st8_809  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[809]), .rdlo_in(a8_wr[813]),  .coef_in(coef[256]), .rdup_out(a9_wr[809]), .rdlo_out(a9_wr[813]));
			radix2 #(.width(width)) rd_st8_810  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[810]), .rdlo_in(a8_wr[814]),  .coef_in(coef[512]), .rdup_out(a9_wr[810]), .rdlo_out(a9_wr[814]));
			radix2 #(.width(width)) rd_st8_811  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[811]), .rdlo_in(a8_wr[815]),  .coef_in(coef[768]), .rdup_out(a9_wr[811]), .rdlo_out(a9_wr[815]));
			radix2 #(.width(width)) rd_st8_816  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[816]), .rdlo_in(a8_wr[820]),  .coef_in(coef[0]), .rdup_out(a9_wr[816]), .rdlo_out(a9_wr[820]));
			radix2 #(.width(width)) rd_st8_817  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[817]), .rdlo_in(a8_wr[821]),  .coef_in(coef[256]), .rdup_out(a9_wr[817]), .rdlo_out(a9_wr[821]));
			radix2 #(.width(width)) rd_st8_818  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[818]), .rdlo_in(a8_wr[822]),  .coef_in(coef[512]), .rdup_out(a9_wr[818]), .rdlo_out(a9_wr[822]));
			radix2 #(.width(width)) rd_st8_819  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[819]), .rdlo_in(a8_wr[823]),  .coef_in(coef[768]), .rdup_out(a9_wr[819]), .rdlo_out(a9_wr[823]));
			radix2 #(.width(width)) rd_st8_824  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[824]), .rdlo_in(a8_wr[828]),  .coef_in(coef[0]), .rdup_out(a9_wr[824]), .rdlo_out(a9_wr[828]));
			radix2 #(.width(width)) rd_st8_825  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[825]), .rdlo_in(a8_wr[829]),  .coef_in(coef[256]), .rdup_out(a9_wr[825]), .rdlo_out(a9_wr[829]));
			radix2 #(.width(width)) rd_st8_826  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[826]), .rdlo_in(a8_wr[830]),  .coef_in(coef[512]), .rdup_out(a9_wr[826]), .rdlo_out(a9_wr[830]));
			radix2 #(.width(width)) rd_st8_827  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[827]), .rdlo_in(a8_wr[831]),  .coef_in(coef[768]), .rdup_out(a9_wr[827]), .rdlo_out(a9_wr[831]));
			radix2 #(.width(width)) rd_st8_832  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[832]), .rdlo_in(a8_wr[836]),  .coef_in(coef[0]), .rdup_out(a9_wr[832]), .rdlo_out(a9_wr[836]));
			radix2 #(.width(width)) rd_st8_833  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[833]), .rdlo_in(a8_wr[837]),  .coef_in(coef[256]), .rdup_out(a9_wr[833]), .rdlo_out(a9_wr[837]));
			radix2 #(.width(width)) rd_st8_834  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[834]), .rdlo_in(a8_wr[838]),  .coef_in(coef[512]), .rdup_out(a9_wr[834]), .rdlo_out(a9_wr[838]));
			radix2 #(.width(width)) rd_st8_835  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[835]), .rdlo_in(a8_wr[839]),  .coef_in(coef[768]), .rdup_out(a9_wr[835]), .rdlo_out(a9_wr[839]));
			radix2 #(.width(width)) rd_st8_840  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[840]), .rdlo_in(a8_wr[844]),  .coef_in(coef[0]), .rdup_out(a9_wr[840]), .rdlo_out(a9_wr[844]));
			radix2 #(.width(width)) rd_st8_841  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[841]), .rdlo_in(a8_wr[845]),  .coef_in(coef[256]), .rdup_out(a9_wr[841]), .rdlo_out(a9_wr[845]));
			radix2 #(.width(width)) rd_st8_842  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[842]), .rdlo_in(a8_wr[846]),  .coef_in(coef[512]), .rdup_out(a9_wr[842]), .rdlo_out(a9_wr[846]));
			radix2 #(.width(width)) rd_st8_843  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[843]), .rdlo_in(a8_wr[847]),  .coef_in(coef[768]), .rdup_out(a9_wr[843]), .rdlo_out(a9_wr[847]));
			radix2 #(.width(width)) rd_st8_848  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[848]), .rdlo_in(a8_wr[852]),  .coef_in(coef[0]), .rdup_out(a9_wr[848]), .rdlo_out(a9_wr[852]));
			radix2 #(.width(width)) rd_st8_849  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[849]), .rdlo_in(a8_wr[853]),  .coef_in(coef[256]), .rdup_out(a9_wr[849]), .rdlo_out(a9_wr[853]));
			radix2 #(.width(width)) rd_st8_850  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[850]), .rdlo_in(a8_wr[854]),  .coef_in(coef[512]), .rdup_out(a9_wr[850]), .rdlo_out(a9_wr[854]));
			radix2 #(.width(width)) rd_st8_851  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[851]), .rdlo_in(a8_wr[855]),  .coef_in(coef[768]), .rdup_out(a9_wr[851]), .rdlo_out(a9_wr[855]));
			radix2 #(.width(width)) rd_st8_856  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[856]), .rdlo_in(a8_wr[860]),  .coef_in(coef[0]), .rdup_out(a9_wr[856]), .rdlo_out(a9_wr[860]));
			radix2 #(.width(width)) rd_st8_857  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[857]), .rdlo_in(a8_wr[861]),  .coef_in(coef[256]), .rdup_out(a9_wr[857]), .rdlo_out(a9_wr[861]));
			radix2 #(.width(width)) rd_st8_858  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[858]), .rdlo_in(a8_wr[862]),  .coef_in(coef[512]), .rdup_out(a9_wr[858]), .rdlo_out(a9_wr[862]));
			radix2 #(.width(width)) rd_st8_859  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[859]), .rdlo_in(a8_wr[863]),  .coef_in(coef[768]), .rdup_out(a9_wr[859]), .rdlo_out(a9_wr[863]));
			radix2 #(.width(width)) rd_st8_864  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[864]), .rdlo_in(a8_wr[868]),  .coef_in(coef[0]), .rdup_out(a9_wr[864]), .rdlo_out(a9_wr[868]));
			radix2 #(.width(width)) rd_st8_865  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[865]), .rdlo_in(a8_wr[869]),  .coef_in(coef[256]), .rdup_out(a9_wr[865]), .rdlo_out(a9_wr[869]));
			radix2 #(.width(width)) rd_st8_866  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[866]), .rdlo_in(a8_wr[870]),  .coef_in(coef[512]), .rdup_out(a9_wr[866]), .rdlo_out(a9_wr[870]));
			radix2 #(.width(width)) rd_st8_867  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[867]), .rdlo_in(a8_wr[871]),  .coef_in(coef[768]), .rdup_out(a9_wr[867]), .rdlo_out(a9_wr[871]));
			radix2 #(.width(width)) rd_st8_872  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[872]), .rdlo_in(a8_wr[876]),  .coef_in(coef[0]), .rdup_out(a9_wr[872]), .rdlo_out(a9_wr[876]));
			radix2 #(.width(width)) rd_st8_873  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[873]), .rdlo_in(a8_wr[877]),  .coef_in(coef[256]), .rdup_out(a9_wr[873]), .rdlo_out(a9_wr[877]));
			radix2 #(.width(width)) rd_st8_874  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[874]), .rdlo_in(a8_wr[878]),  .coef_in(coef[512]), .rdup_out(a9_wr[874]), .rdlo_out(a9_wr[878]));
			radix2 #(.width(width)) rd_st8_875  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[875]), .rdlo_in(a8_wr[879]),  .coef_in(coef[768]), .rdup_out(a9_wr[875]), .rdlo_out(a9_wr[879]));
			radix2 #(.width(width)) rd_st8_880  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[880]), .rdlo_in(a8_wr[884]),  .coef_in(coef[0]), .rdup_out(a9_wr[880]), .rdlo_out(a9_wr[884]));
			radix2 #(.width(width)) rd_st8_881  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[881]), .rdlo_in(a8_wr[885]),  .coef_in(coef[256]), .rdup_out(a9_wr[881]), .rdlo_out(a9_wr[885]));
			radix2 #(.width(width)) rd_st8_882  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[882]), .rdlo_in(a8_wr[886]),  .coef_in(coef[512]), .rdup_out(a9_wr[882]), .rdlo_out(a9_wr[886]));
			radix2 #(.width(width)) rd_st8_883  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[883]), .rdlo_in(a8_wr[887]),  .coef_in(coef[768]), .rdup_out(a9_wr[883]), .rdlo_out(a9_wr[887]));
			radix2 #(.width(width)) rd_st8_888  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[888]), .rdlo_in(a8_wr[892]),  .coef_in(coef[0]), .rdup_out(a9_wr[888]), .rdlo_out(a9_wr[892]));
			radix2 #(.width(width)) rd_st8_889  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[889]), .rdlo_in(a8_wr[893]),  .coef_in(coef[256]), .rdup_out(a9_wr[889]), .rdlo_out(a9_wr[893]));
			radix2 #(.width(width)) rd_st8_890  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[890]), .rdlo_in(a8_wr[894]),  .coef_in(coef[512]), .rdup_out(a9_wr[890]), .rdlo_out(a9_wr[894]));
			radix2 #(.width(width)) rd_st8_891  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[891]), .rdlo_in(a8_wr[895]),  .coef_in(coef[768]), .rdup_out(a9_wr[891]), .rdlo_out(a9_wr[895]));
			radix2 #(.width(width)) rd_st8_896  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[896]), .rdlo_in(a8_wr[900]),  .coef_in(coef[0]), .rdup_out(a9_wr[896]), .rdlo_out(a9_wr[900]));
			radix2 #(.width(width)) rd_st8_897  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[897]), .rdlo_in(a8_wr[901]),  .coef_in(coef[256]), .rdup_out(a9_wr[897]), .rdlo_out(a9_wr[901]));
			radix2 #(.width(width)) rd_st8_898  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[898]), .rdlo_in(a8_wr[902]),  .coef_in(coef[512]), .rdup_out(a9_wr[898]), .rdlo_out(a9_wr[902]));
			radix2 #(.width(width)) rd_st8_899  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[899]), .rdlo_in(a8_wr[903]),  .coef_in(coef[768]), .rdup_out(a9_wr[899]), .rdlo_out(a9_wr[903]));
			radix2 #(.width(width)) rd_st8_904  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[904]), .rdlo_in(a8_wr[908]),  .coef_in(coef[0]), .rdup_out(a9_wr[904]), .rdlo_out(a9_wr[908]));
			radix2 #(.width(width)) rd_st8_905  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[905]), .rdlo_in(a8_wr[909]),  .coef_in(coef[256]), .rdup_out(a9_wr[905]), .rdlo_out(a9_wr[909]));
			radix2 #(.width(width)) rd_st8_906  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[906]), .rdlo_in(a8_wr[910]),  .coef_in(coef[512]), .rdup_out(a9_wr[906]), .rdlo_out(a9_wr[910]));
			radix2 #(.width(width)) rd_st8_907  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[907]), .rdlo_in(a8_wr[911]),  .coef_in(coef[768]), .rdup_out(a9_wr[907]), .rdlo_out(a9_wr[911]));
			radix2 #(.width(width)) rd_st8_912  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[912]), .rdlo_in(a8_wr[916]),  .coef_in(coef[0]), .rdup_out(a9_wr[912]), .rdlo_out(a9_wr[916]));
			radix2 #(.width(width)) rd_st8_913  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[913]), .rdlo_in(a8_wr[917]),  .coef_in(coef[256]), .rdup_out(a9_wr[913]), .rdlo_out(a9_wr[917]));
			radix2 #(.width(width)) rd_st8_914  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[914]), .rdlo_in(a8_wr[918]),  .coef_in(coef[512]), .rdup_out(a9_wr[914]), .rdlo_out(a9_wr[918]));
			radix2 #(.width(width)) rd_st8_915  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[915]), .rdlo_in(a8_wr[919]),  .coef_in(coef[768]), .rdup_out(a9_wr[915]), .rdlo_out(a9_wr[919]));
			radix2 #(.width(width)) rd_st8_920  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[920]), .rdlo_in(a8_wr[924]),  .coef_in(coef[0]), .rdup_out(a9_wr[920]), .rdlo_out(a9_wr[924]));
			radix2 #(.width(width)) rd_st8_921  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[921]), .rdlo_in(a8_wr[925]),  .coef_in(coef[256]), .rdup_out(a9_wr[921]), .rdlo_out(a9_wr[925]));
			radix2 #(.width(width)) rd_st8_922  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[922]), .rdlo_in(a8_wr[926]),  .coef_in(coef[512]), .rdup_out(a9_wr[922]), .rdlo_out(a9_wr[926]));
			radix2 #(.width(width)) rd_st8_923  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[923]), .rdlo_in(a8_wr[927]),  .coef_in(coef[768]), .rdup_out(a9_wr[923]), .rdlo_out(a9_wr[927]));
			radix2 #(.width(width)) rd_st8_928  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[928]), .rdlo_in(a8_wr[932]),  .coef_in(coef[0]), .rdup_out(a9_wr[928]), .rdlo_out(a9_wr[932]));
			radix2 #(.width(width)) rd_st8_929  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[929]), .rdlo_in(a8_wr[933]),  .coef_in(coef[256]), .rdup_out(a9_wr[929]), .rdlo_out(a9_wr[933]));
			radix2 #(.width(width)) rd_st8_930  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[930]), .rdlo_in(a8_wr[934]),  .coef_in(coef[512]), .rdup_out(a9_wr[930]), .rdlo_out(a9_wr[934]));
			radix2 #(.width(width)) rd_st8_931  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[931]), .rdlo_in(a8_wr[935]),  .coef_in(coef[768]), .rdup_out(a9_wr[931]), .rdlo_out(a9_wr[935]));
			radix2 #(.width(width)) rd_st8_936  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[936]), .rdlo_in(a8_wr[940]),  .coef_in(coef[0]), .rdup_out(a9_wr[936]), .rdlo_out(a9_wr[940]));
			radix2 #(.width(width)) rd_st8_937  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[937]), .rdlo_in(a8_wr[941]),  .coef_in(coef[256]), .rdup_out(a9_wr[937]), .rdlo_out(a9_wr[941]));
			radix2 #(.width(width)) rd_st8_938  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[938]), .rdlo_in(a8_wr[942]),  .coef_in(coef[512]), .rdup_out(a9_wr[938]), .rdlo_out(a9_wr[942]));
			radix2 #(.width(width)) rd_st8_939  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[939]), .rdlo_in(a8_wr[943]),  .coef_in(coef[768]), .rdup_out(a9_wr[939]), .rdlo_out(a9_wr[943]));
			radix2 #(.width(width)) rd_st8_944  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[944]), .rdlo_in(a8_wr[948]),  .coef_in(coef[0]), .rdup_out(a9_wr[944]), .rdlo_out(a9_wr[948]));
			radix2 #(.width(width)) rd_st8_945  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[945]), .rdlo_in(a8_wr[949]),  .coef_in(coef[256]), .rdup_out(a9_wr[945]), .rdlo_out(a9_wr[949]));
			radix2 #(.width(width)) rd_st8_946  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[946]), .rdlo_in(a8_wr[950]),  .coef_in(coef[512]), .rdup_out(a9_wr[946]), .rdlo_out(a9_wr[950]));
			radix2 #(.width(width)) rd_st8_947  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[947]), .rdlo_in(a8_wr[951]),  .coef_in(coef[768]), .rdup_out(a9_wr[947]), .rdlo_out(a9_wr[951]));
			radix2 #(.width(width)) rd_st8_952  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[952]), .rdlo_in(a8_wr[956]),  .coef_in(coef[0]), .rdup_out(a9_wr[952]), .rdlo_out(a9_wr[956]));
			radix2 #(.width(width)) rd_st8_953  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[953]), .rdlo_in(a8_wr[957]),  .coef_in(coef[256]), .rdup_out(a9_wr[953]), .rdlo_out(a9_wr[957]));
			radix2 #(.width(width)) rd_st8_954  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[954]), .rdlo_in(a8_wr[958]),  .coef_in(coef[512]), .rdup_out(a9_wr[954]), .rdlo_out(a9_wr[958]));
			radix2 #(.width(width)) rd_st8_955  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[955]), .rdlo_in(a8_wr[959]),  .coef_in(coef[768]), .rdup_out(a9_wr[955]), .rdlo_out(a9_wr[959]));
			radix2 #(.width(width)) rd_st8_960  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[960]), .rdlo_in(a8_wr[964]),  .coef_in(coef[0]), .rdup_out(a9_wr[960]), .rdlo_out(a9_wr[964]));
			radix2 #(.width(width)) rd_st8_961  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[961]), .rdlo_in(a8_wr[965]),  .coef_in(coef[256]), .rdup_out(a9_wr[961]), .rdlo_out(a9_wr[965]));
			radix2 #(.width(width)) rd_st8_962  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[962]), .rdlo_in(a8_wr[966]),  .coef_in(coef[512]), .rdup_out(a9_wr[962]), .rdlo_out(a9_wr[966]));
			radix2 #(.width(width)) rd_st8_963  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[963]), .rdlo_in(a8_wr[967]),  .coef_in(coef[768]), .rdup_out(a9_wr[963]), .rdlo_out(a9_wr[967]));
			radix2 #(.width(width)) rd_st8_968  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[968]), .rdlo_in(a8_wr[972]),  .coef_in(coef[0]), .rdup_out(a9_wr[968]), .rdlo_out(a9_wr[972]));
			radix2 #(.width(width)) rd_st8_969  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[969]), .rdlo_in(a8_wr[973]),  .coef_in(coef[256]), .rdup_out(a9_wr[969]), .rdlo_out(a9_wr[973]));
			radix2 #(.width(width)) rd_st8_970  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[970]), .rdlo_in(a8_wr[974]),  .coef_in(coef[512]), .rdup_out(a9_wr[970]), .rdlo_out(a9_wr[974]));
			radix2 #(.width(width)) rd_st8_971  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[971]), .rdlo_in(a8_wr[975]),  .coef_in(coef[768]), .rdup_out(a9_wr[971]), .rdlo_out(a9_wr[975]));
			radix2 #(.width(width)) rd_st8_976  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[976]), .rdlo_in(a8_wr[980]),  .coef_in(coef[0]), .rdup_out(a9_wr[976]), .rdlo_out(a9_wr[980]));
			radix2 #(.width(width)) rd_st8_977  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[977]), .rdlo_in(a8_wr[981]),  .coef_in(coef[256]), .rdup_out(a9_wr[977]), .rdlo_out(a9_wr[981]));
			radix2 #(.width(width)) rd_st8_978  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[978]), .rdlo_in(a8_wr[982]),  .coef_in(coef[512]), .rdup_out(a9_wr[978]), .rdlo_out(a9_wr[982]));
			radix2 #(.width(width)) rd_st8_979  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[979]), .rdlo_in(a8_wr[983]),  .coef_in(coef[768]), .rdup_out(a9_wr[979]), .rdlo_out(a9_wr[983]));
			radix2 #(.width(width)) rd_st8_984  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[984]), .rdlo_in(a8_wr[988]),  .coef_in(coef[0]), .rdup_out(a9_wr[984]), .rdlo_out(a9_wr[988]));
			radix2 #(.width(width)) rd_st8_985  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[985]), .rdlo_in(a8_wr[989]),  .coef_in(coef[256]), .rdup_out(a9_wr[985]), .rdlo_out(a9_wr[989]));
			radix2 #(.width(width)) rd_st8_986  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[986]), .rdlo_in(a8_wr[990]),  .coef_in(coef[512]), .rdup_out(a9_wr[986]), .rdlo_out(a9_wr[990]));
			radix2 #(.width(width)) rd_st8_987  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[987]), .rdlo_in(a8_wr[991]),  .coef_in(coef[768]), .rdup_out(a9_wr[987]), .rdlo_out(a9_wr[991]));
			radix2 #(.width(width)) rd_st8_992  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[992]), .rdlo_in(a8_wr[996]),  .coef_in(coef[0]), .rdup_out(a9_wr[992]), .rdlo_out(a9_wr[996]));
			radix2 #(.width(width)) rd_st8_993  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[993]), .rdlo_in(a8_wr[997]),  .coef_in(coef[256]), .rdup_out(a9_wr[993]), .rdlo_out(a9_wr[997]));
			radix2 #(.width(width)) rd_st8_994  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[994]), .rdlo_in(a8_wr[998]),  .coef_in(coef[512]), .rdup_out(a9_wr[994]), .rdlo_out(a9_wr[998]));
			radix2 #(.width(width)) rd_st8_995  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[995]), .rdlo_in(a8_wr[999]),  .coef_in(coef[768]), .rdup_out(a9_wr[995]), .rdlo_out(a9_wr[999]));
			radix2 #(.width(width)) rd_st8_1000  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1000]), .rdlo_in(a8_wr[1004]),  .coef_in(coef[0]), .rdup_out(a9_wr[1000]), .rdlo_out(a9_wr[1004]));
			radix2 #(.width(width)) rd_st8_1001  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1001]), .rdlo_in(a8_wr[1005]),  .coef_in(coef[256]), .rdup_out(a9_wr[1001]), .rdlo_out(a9_wr[1005]));
			radix2 #(.width(width)) rd_st8_1002  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1002]), .rdlo_in(a8_wr[1006]),  .coef_in(coef[512]), .rdup_out(a9_wr[1002]), .rdlo_out(a9_wr[1006]));
			radix2 #(.width(width)) rd_st8_1003  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1003]), .rdlo_in(a8_wr[1007]),  .coef_in(coef[768]), .rdup_out(a9_wr[1003]), .rdlo_out(a9_wr[1007]));
			radix2 #(.width(width)) rd_st8_1008  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1008]), .rdlo_in(a8_wr[1012]),  .coef_in(coef[0]), .rdup_out(a9_wr[1008]), .rdlo_out(a9_wr[1012]));
			radix2 #(.width(width)) rd_st8_1009  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1009]), .rdlo_in(a8_wr[1013]),  .coef_in(coef[256]), .rdup_out(a9_wr[1009]), .rdlo_out(a9_wr[1013]));
			radix2 #(.width(width)) rd_st8_1010  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1010]), .rdlo_in(a8_wr[1014]),  .coef_in(coef[512]), .rdup_out(a9_wr[1010]), .rdlo_out(a9_wr[1014]));
			radix2 #(.width(width)) rd_st8_1011  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1011]), .rdlo_in(a8_wr[1015]),  .coef_in(coef[768]), .rdup_out(a9_wr[1011]), .rdlo_out(a9_wr[1015]));
			radix2 #(.width(width)) rd_st8_1016  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1016]), .rdlo_in(a8_wr[1020]),  .coef_in(coef[0]), .rdup_out(a9_wr[1016]), .rdlo_out(a9_wr[1020]));
			radix2 #(.width(width)) rd_st8_1017  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1017]), .rdlo_in(a8_wr[1021]),  .coef_in(coef[256]), .rdup_out(a9_wr[1017]), .rdlo_out(a9_wr[1021]));
			radix2 #(.width(width)) rd_st8_1018  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1018]), .rdlo_in(a8_wr[1022]),  .coef_in(coef[512]), .rdup_out(a9_wr[1018]), .rdlo_out(a9_wr[1022]));
			radix2 #(.width(width)) rd_st8_1019  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1019]), .rdlo_in(a8_wr[1023]),  .coef_in(coef[768]), .rdup_out(a9_wr[1019]), .rdlo_out(a9_wr[1023]));
			radix2 #(.width(width)) rd_st8_1024  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1024]), .rdlo_in(a8_wr[1028]),  .coef_in(coef[0]), .rdup_out(a9_wr[1024]), .rdlo_out(a9_wr[1028]));
			radix2 #(.width(width)) rd_st8_1025  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1025]), .rdlo_in(a8_wr[1029]),  .coef_in(coef[256]), .rdup_out(a9_wr[1025]), .rdlo_out(a9_wr[1029]));
			radix2 #(.width(width)) rd_st8_1026  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1026]), .rdlo_in(a8_wr[1030]),  .coef_in(coef[512]), .rdup_out(a9_wr[1026]), .rdlo_out(a9_wr[1030]));
			radix2 #(.width(width)) rd_st8_1027  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1027]), .rdlo_in(a8_wr[1031]),  .coef_in(coef[768]), .rdup_out(a9_wr[1027]), .rdlo_out(a9_wr[1031]));
			radix2 #(.width(width)) rd_st8_1032  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1032]), .rdlo_in(a8_wr[1036]),  .coef_in(coef[0]), .rdup_out(a9_wr[1032]), .rdlo_out(a9_wr[1036]));
			radix2 #(.width(width)) rd_st8_1033  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1033]), .rdlo_in(a8_wr[1037]),  .coef_in(coef[256]), .rdup_out(a9_wr[1033]), .rdlo_out(a9_wr[1037]));
			radix2 #(.width(width)) rd_st8_1034  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1034]), .rdlo_in(a8_wr[1038]),  .coef_in(coef[512]), .rdup_out(a9_wr[1034]), .rdlo_out(a9_wr[1038]));
			radix2 #(.width(width)) rd_st8_1035  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1035]), .rdlo_in(a8_wr[1039]),  .coef_in(coef[768]), .rdup_out(a9_wr[1035]), .rdlo_out(a9_wr[1039]));
			radix2 #(.width(width)) rd_st8_1040  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1040]), .rdlo_in(a8_wr[1044]),  .coef_in(coef[0]), .rdup_out(a9_wr[1040]), .rdlo_out(a9_wr[1044]));
			radix2 #(.width(width)) rd_st8_1041  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1041]), .rdlo_in(a8_wr[1045]),  .coef_in(coef[256]), .rdup_out(a9_wr[1041]), .rdlo_out(a9_wr[1045]));
			radix2 #(.width(width)) rd_st8_1042  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1042]), .rdlo_in(a8_wr[1046]),  .coef_in(coef[512]), .rdup_out(a9_wr[1042]), .rdlo_out(a9_wr[1046]));
			radix2 #(.width(width)) rd_st8_1043  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1043]), .rdlo_in(a8_wr[1047]),  .coef_in(coef[768]), .rdup_out(a9_wr[1043]), .rdlo_out(a9_wr[1047]));
			radix2 #(.width(width)) rd_st8_1048  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1048]), .rdlo_in(a8_wr[1052]),  .coef_in(coef[0]), .rdup_out(a9_wr[1048]), .rdlo_out(a9_wr[1052]));
			radix2 #(.width(width)) rd_st8_1049  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1049]), .rdlo_in(a8_wr[1053]),  .coef_in(coef[256]), .rdup_out(a9_wr[1049]), .rdlo_out(a9_wr[1053]));
			radix2 #(.width(width)) rd_st8_1050  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1050]), .rdlo_in(a8_wr[1054]),  .coef_in(coef[512]), .rdup_out(a9_wr[1050]), .rdlo_out(a9_wr[1054]));
			radix2 #(.width(width)) rd_st8_1051  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1051]), .rdlo_in(a8_wr[1055]),  .coef_in(coef[768]), .rdup_out(a9_wr[1051]), .rdlo_out(a9_wr[1055]));
			radix2 #(.width(width)) rd_st8_1056  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1056]), .rdlo_in(a8_wr[1060]),  .coef_in(coef[0]), .rdup_out(a9_wr[1056]), .rdlo_out(a9_wr[1060]));
			radix2 #(.width(width)) rd_st8_1057  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1057]), .rdlo_in(a8_wr[1061]),  .coef_in(coef[256]), .rdup_out(a9_wr[1057]), .rdlo_out(a9_wr[1061]));
			radix2 #(.width(width)) rd_st8_1058  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1058]), .rdlo_in(a8_wr[1062]),  .coef_in(coef[512]), .rdup_out(a9_wr[1058]), .rdlo_out(a9_wr[1062]));
			radix2 #(.width(width)) rd_st8_1059  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1059]), .rdlo_in(a8_wr[1063]),  .coef_in(coef[768]), .rdup_out(a9_wr[1059]), .rdlo_out(a9_wr[1063]));
			radix2 #(.width(width)) rd_st8_1064  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1064]), .rdlo_in(a8_wr[1068]),  .coef_in(coef[0]), .rdup_out(a9_wr[1064]), .rdlo_out(a9_wr[1068]));
			radix2 #(.width(width)) rd_st8_1065  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1065]), .rdlo_in(a8_wr[1069]),  .coef_in(coef[256]), .rdup_out(a9_wr[1065]), .rdlo_out(a9_wr[1069]));
			radix2 #(.width(width)) rd_st8_1066  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1066]), .rdlo_in(a8_wr[1070]),  .coef_in(coef[512]), .rdup_out(a9_wr[1066]), .rdlo_out(a9_wr[1070]));
			radix2 #(.width(width)) rd_st8_1067  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1067]), .rdlo_in(a8_wr[1071]),  .coef_in(coef[768]), .rdup_out(a9_wr[1067]), .rdlo_out(a9_wr[1071]));
			radix2 #(.width(width)) rd_st8_1072  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1072]), .rdlo_in(a8_wr[1076]),  .coef_in(coef[0]), .rdup_out(a9_wr[1072]), .rdlo_out(a9_wr[1076]));
			radix2 #(.width(width)) rd_st8_1073  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1073]), .rdlo_in(a8_wr[1077]),  .coef_in(coef[256]), .rdup_out(a9_wr[1073]), .rdlo_out(a9_wr[1077]));
			radix2 #(.width(width)) rd_st8_1074  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1074]), .rdlo_in(a8_wr[1078]),  .coef_in(coef[512]), .rdup_out(a9_wr[1074]), .rdlo_out(a9_wr[1078]));
			radix2 #(.width(width)) rd_st8_1075  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1075]), .rdlo_in(a8_wr[1079]),  .coef_in(coef[768]), .rdup_out(a9_wr[1075]), .rdlo_out(a9_wr[1079]));
			radix2 #(.width(width)) rd_st8_1080  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1080]), .rdlo_in(a8_wr[1084]),  .coef_in(coef[0]), .rdup_out(a9_wr[1080]), .rdlo_out(a9_wr[1084]));
			radix2 #(.width(width)) rd_st8_1081  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1081]), .rdlo_in(a8_wr[1085]),  .coef_in(coef[256]), .rdup_out(a9_wr[1081]), .rdlo_out(a9_wr[1085]));
			radix2 #(.width(width)) rd_st8_1082  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1082]), .rdlo_in(a8_wr[1086]),  .coef_in(coef[512]), .rdup_out(a9_wr[1082]), .rdlo_out(a9_wr[1086]));
			radix2 #(.width(width)) rd_st8_1083  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1083]), .rdlo_in(a8_wr[1087]),  .coef_in(coef[768]), .rdup_out(a9_wr[1083]), .rdlo_out(a9_wr[1087]));
			radix2 #(.width(width)) rd_st8_1088  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1088]), .rdlo_in(a8_wr[1092]),  .coef_in(coef[0]), .rdup_out(a9_wr[1088]), .rdlo_out(a9_wr[1092]));
			radix2 #(.width(width)) rd_st8_1089  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1089]), .rdlo_in(a8_wr[1093]),  .coef_in(coef[256]), .rdup_out(a9_wr[1089]), .rdlo_out(a9_wr[1093]));
			radix2 #(.width(width)) rd_st8_1090  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1090]), .rdlo_in(a8_wr[1094]),  .coef_in(coef[512]), .rdup_out(a9_wr[1090]), .rdlo_out(a9_wr[1094]));
			radix2 #(.width(width)) rd_st8_1091  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1091]), .rdlo_in(a8_wr[1095]),  .coef_in(coef[768]), .rdup_out(a9_wr[1091]), .rdlo_out(a9_wr[1095]));
			radix2 #(.width(width)) rd_st8_1096  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1096]), .rdlo_in(a8_wr[1100]),  .coef_in(coef[0]), .rdup_out(a9_wr[1096]), .rdlo_out(a9_wr[1100]));
			radix2 #(.width(width)) rd_st8_1097  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1097]), .rdlo_in(a8_wr[1101]),  .coef_in(coef[256]), .rdup_out(a9_wr[1097]), .rdlo_out(a9_wr[1101]));
			radix2 #(.width(width)) rd_st8_1098  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1098]), .rdlo_in(a8_wr[1102]),  .coef_in(coef[512]), .rdup_out(a9_wr[1098]), .rdlo_out(a9_wr[1102]));
			radix2 #(.width(width)) rd_st8_1099  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1099]), .rdlo_in(a8_wr[1103]),  .coef_in(coef[768]), .rdup_out(a9_wr[1099]), .rdlo_out(a9_wr[1103]));
			radix2 #(.width(width)) rd_st8_1104  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1104]), .rdlo_in(a8_wr[1108]),  .coef_in(coef[0]), .rdup_out(a9_wr[1104]), .rdlo_out(a9_wr[1108]));
			radix2 #(.width(width)) rd_st8_1105  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1105]), .rdlo_in(a8_wr[1109]),  .coef_in(coef[256]), .rdup_out(a9_wr[1105]), .rdlo_out(a9_wr[1109]));
			radix2 #(.width(width)) rd_st8_1106  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1106]), .rdlo_in(a8_wr[1110]),  .coef_in(coef[512]), .rdup_out(a9_wr[1106]), .rdlo_out(a9_wr[1110]));
			radix2 #(.width(width)) rd_st8_1107  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1107]), .rdlo_in(a8_wr[1111]),  .coef_in(coef[768]), .rdup_out(a9_wr[1107]), .rdlo_out(a9_wr[1111]));
			radix2 #(.width(width)) rd_st8_1112  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1112]), .rdlo_in(a8_wr[1116]),  .coef_in(coef[0]), .rdup_out(a9_wr[1112]), .rdlo_out(a9_wr[1116]));
			radix2 #(.width(width)) rd_st8_1113  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1113]), .rdlo_in(a8_wr[1117]),  .coef_in(coef[256]), .rdup_out(a9_wr[1113]), .rdlo_out(a9_wr[1117]));
			radix2 #(.width(width)) rd_st8_1114  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1114]), .rdlo_in(a8_wr[1118]),  .coef_in(coef[512]), .rdup_out(a9_wr[1114]), .rdlo_out(a9_wr[1118]));
			radix2 #(.width(width)) rd_st8_1115  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1115]), .rdlo_in(a8_wr[1119]),  .coef_in(coef[768]), .rdup_out(a9_wr[1115]), .rdlo_out(a9_wr[1119]));
			radix2 #(.width(width)) rd_st8_1120  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1120]), .rdlo_in(a8_wr[1124]),  .coef_in(coef[0]), .rdup_out(a9_wr[1120]), .rdlo_out(a9_wr[1124]));
			radix2 #(.width(width)) rd_st8_1121  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1121]), .rdlo_in(a8_wr[1125]),  .coef_in(coef[256]), .rdup_out(a9_wr[1121]), .rdlo_out(a9_wr[1125]));
			radix2 #(.width(width)) rd_st8_1122  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1122]), .rdlo_in(a8_wr[1126]),  .coef_in(coef[512]), .rdup_out(a9_wr[1122]), .rdlo_out(a9_wr[1126]));
			radix2 #(.width(width)) rd_st8_1123  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1123]), .rdlo_in(a8_wr[1127]),  .coef_in(coef[768]), .rdup_out(a9_wr[1123]), .rdlo_out(a9_wr[1127]));
			radix2 #(.width(width)) rd_st8_1128  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1128]), .rdlo_in(a8_wr[1132]),  .coef_in(coef[0]), .rdup_out(a9_wr[1128]), .rdlo_out(a9_wr[1132]));
			radix2 #(.width(width)) rd_st8_1129  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1129]), .rdlo_in(a8_wr[1133]),  .coef_in(coef[256]), .rdup_out(a9_wr[1129]), .rdlo_out(a9_wr[1133]));
			radix2 #(.width(width)) rd_st8_1130  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1130]), .rdlo_in(a8_wr[1134]),  .coef_in(coef[512]), .rdup_out(a9_wr[1130]), .rdlo_out(a9_wr[1134]));
			radix2 #(.width(width)) rd_st8_1131  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1131]), .rdlo_in(a8_wr[1135]),  .coef_in(coef[768]), .rdup_out(a9_wr[1131]), .rdlo_out(a9_wr[1135]));
			radix2 #(.width(width)) rd_st8_1136  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1136]), .rdlo_in(a8_wr[1140]),  .coef_in(coef[0]), .rdup_out(a9_wr[1136]), .rdlo_out(a9_wr[1140]));
			radix2 #(.width(width)) rd_st8_1137  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1137]), .rdlo_in(a8_wr[1141]),  .coef_in(coef[256]), .rdup_out(a9_wr[1137]), .rdlo_out(a9_wr[1141]));
			radix2 #(.width(width)) rd_st8_1138  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1138]), .rdlo_in(a8_wr[1142]),  .coef_in(coef[512]), .rdup_out(a9_wr[1138]), .rdlo_out(a9_wr[1142]));
			radix2 #(.width(width)) rd_st8_1139  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1139]), .rdlo_in(a8_wr[1143]),  .coef_in(coef[768]), .rdup_out(a9_wr[1139]), .rdlo_out(a9_wr[1143]));
			radix2 #(.width(width)) rd_st8_1144  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1144]), .rdlo_in(a8_wr[1148]),  .coef_in(coef[0]), .rdup_out(a9_wr[1144]), .rdlo_out(a9_wr[1148]));
			radix2 #(.width(width)) rd_st8_1145  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1145]), .rdlo_in(a8_wr[1149]),  .coef_in(coef[256]), .rdup_out(a9_wr[1145]), .rdlo_out(a9_wr[1149]));
			radix2 #(.width(width)) rd_st8_1146  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1146]), .rdlo_in(a8_wr[1150]),  .coef_in(coef[512]), .rdup_out(a9_wr[1146]), .rdlo_out(a9_wr[1150]));
			radix2 #(.width(width)) rd_st8_1147  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1147]), .rdlo_in(a8_wr[1151]),  .coef_in(coef[768]), .rdup_out(a9_wr[1147]), .rdlo_out(a9_wr[1151]));
			radix2 #(.width(width)) rd_st8_1152  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1152]), .rdlo_in(a8_wr[1156]),  .coef_in(coef[0]), .rdup_out(a9_wr[1152]), .rdlo_out(a9_wr[1156]));
			radix2 #(.width(width)) rd_st8_1153  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1153]), .rdlo_in(a8_wr[1157]),  .coef_in(coef[256]), .rdup_out(a9_wr[1153]), .rdlo_out(a9_wr[1157]));
			radix2 #(.width(width)) rd_st8_1154  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1154]), .rdlo_in(a8_wr[1158]),  .coef_in(coef[512]), .rdup_out(a9_wr[1154]), .rdlo_out(a9_wr[1158]));
			radix2 #(.width(width)) rd_st8_1155  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1155]), .rdlo_in(a8_wr[1159]),  .coef_in(coef[768]), .rdup_out(a9_wr[1155]), .rdlo_out(a9_wr[1159]));
			radix2 #(.width(width)) rd_st8_1160  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1160]), .rdlo_in(a8_wr[1164]),  .coef_in(coef[0]), .rdup_out(a9_wr[1160]), .rdlo_out(a9_wr[1164]));
			radix2 #(.width(width)) rd_st8_1161  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1161]), .rdlo_in(a8_wr[1165]),  .coef_in(coef[256]), .rdup_out(a9_wr[1161]), .rdlo_out(a9_wr[1165]));
			radix2 #(.width(width)) rd_st8_1162  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1162]), .rdlo_in(a8_wr[1166]),  .coef_in(coef[512]), .rdup_out(a9_wr[1162]), .rdlo_out(a9_wr[1166]));
			radix2 #(.width(width)) rd_st8_1163  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1163]), .rdlo_in(a8_wr[1167]),  .coef_in(coef[768]), .rdup_out(a9_wr[1163]), .rdlo_out(a9_wr[1167]));
			radix2 #(.width(width)) rd_st8_1168  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1168]), .rdlo_in(a8_wr[1172]),  .coef_in(coef[0]), .rdup_out(a9_wr[1168]), .rdlo_out(a9_wr[1172]));
			radix2 #(.width(width)) rd_st8_1169  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1169]), .rdlo_in(a8_wr[1173]),  .coef_in(coef[256]), .rdup_out(a9_wr[1169]), .rdlo_out(a9_wr[1173]));
			radix2 #(.width(width)) rd_st8_1170  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1170]), .rdlo_in(a8_wr[1174]),  .coef_in(coef[512]), .rdup_out(a9_wr[1170]), .rdlo_out(a9_wr[1174]));
			radix2 #(.width(width)) rd_st8_1171  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1171]), .rdlo_in(a8_wr[1175]),  .coef_in(coef[768]), .rdup_out(a9_wr[1171]), .rdlo_out(a9_wr[1175]));
			radix2 #(.width(width)) rd_st8_1176  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1176]), .rdlo_in(a8_wr[1180]),  .coef_in(coef[0]), .rdup_out(a9_wr[1176]), .rdlo_out(a9_wr[1180]));
			radix2 #(.width(width)) rd_st8_1177  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1177]), .rdlo_in(a8_wr[1181]),  .coef_in(coef[256]), .rdup_out(a9_wr[1177]), .rdlo_out(a9_wr[1181]));
			radix2 #(.width(width)) rd_st8_1178  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1178]), .rdlo_in(a8_wr[1182]),  .coef_in(coef[512]), .rdup_out(a9_wr[1178]), .rdlo_out(a9_wr[1182]));
			radix2 #(.width(width)) rd_st8_1179  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1179]), .rdlo_in(a8_wr[1183]),  .coef_in(coef[768]), .rdup_out(a9_wr[1179]), .rdlo_out(a9_wr[1183]));
			radix2 #(.width(width)) rd_st8_1184  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1184]), .rdlo_in(a8_wr[1188]),  .coef_in(coef[0]), .rdup_out(a9_wr[1184]), .rdlo_out(a9_wr[1188]));
			radix2 #(.width(width)) rd_st8_1185  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1185]), .rdlo_in(a8_wr[1189]),  .coef_in(coef[256]), .rdup_out(a9_wr[1185]), .rdlo_out(a9_wr[1189]));
			radix2 #(.width(width)) rd_st8_1186  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1186]), .rdlo_in(a8_wr[1190]),  .coef_in(coef[512]), .rdup_out(a9_wr[1186]), .rdlo_out(a9_wr[1190]));
			radix2 #(.width(width)) rd_st8_1187  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1187]), .rdlo_in(a8_wr[1191]),  .coef_in(coef[768]), .rdup_out(a9_wr[1187]), .rdlo_out(a9_wr[1191]));
			radix2 #(.width(width)) rd_st8_1192  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1192]), .rdlo_in(a8_wr[1196]),  .coef_in(coef[0]), .rdup_out(a9_wr[1192]), .rdlo_out(a9_wr[1196]));
			radix2 #(.width(width)) rd_st8_1193  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1193]), .rdlo_in(a8_wr[1197]),  .coef_in(coef[256]), .rdup_out(a9_wr[1193]), .rdlo_out(a9_wr[1197]));
			radix2 #(.width(width)) rd_st8_1194  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1194]), .rdlo_in(a8_wr[1198]),  .coef_in(coef[512]), .rdup_out(a9_wr[1194]), .rdlo_out(a9_wr[1198]));
			radix2 #(.width(width)) rd_st8_1195  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1195]), .rdlo_in(a8_wr[1199]),  .coef_in(coef[768]), .rdup_out(a9_wr[1195]), .rdlo_out(a9_wr[1199]));
			radix2 #(.width(width)) rd_st8_1200  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1200]), .rdlo_in(a8_wr[1204]),  .coef_in(coef[0]), .rdup_out(a9_wr[1200]), .rdlo_out(a9_wr[1204]));
			radix2 #(.width(width)) rd_st8_1201  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1201]), .rdlo_in(a8_wr[1205]),  .coef_in(coef[256]), .rdup_out(a9_wr[1201]), .rdlo_out(a9_wr[1205]));
			radix2 #(.width(width)) rd_st8_1202  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1202]), .rdlo_in(a8_wr[1206]),  .coef_in(coef[512]), .rdup_out(a9_wr[1202]), .rdlo_out(a9_wr[1206]));
			radix2 #(.width(width)) rd_st8_1203  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1203]), .rdlo_in(a8_wr[1207]),  .coef_in(coef[768]), .rdup_out(a9_wr[1203]), .rdlo_out(a9_wr[1207]));
			radix2 #(.width(width)) rd_st8_1208  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1208]), .rdlo_in(a8_wr[1212]),  .coef_in(coef[0]), .rdup_out(a9_wr[1208]), .rdlo_out(a9_wr[1212]));
			radix2 #(.width(width)) rd_st8_1209  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1209]), .rdlo_in(a8_wr[1213]),  .coef_in(coef[256]), .rdup_out(a9_wr[1209]), .rdlo_out(a9_wr[1213]));
			radix2 #(.width(width)) rd_st8_1210  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1210]), .rdlo_in(a8_wr[1214]),  .coef_in(coef[512]), .rdup_out(a9_wr[1210]), .rdlo_out(a9_wr[1214]));
			radix2 #(.width(width)) rd_st8_1211  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1211]), .rdlo_in(a8_wr[1215]),  .coef_in(coef[768]), .rdup_out(a9_wr[1211]), .rdlo_out(a9_wr[1215]));
			radix2 #(.width(width)) rd_st8_1216  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1216]), .rdlo_in(a8_wr[1220]),  .coef_in(coef[0]), .rdup_out(a9_wr[1216]), .rdlo_out(a9_wr[1220]));
			radix2 #(.width(width)) rd_st8_1217  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1217]), .rdlo_in(a8_wr[1221]),  .coef_in(coef[256]), .rdup_out(a9_wr[1217]), .rdlo_out(a9_wr[1221]));
			radix2 #(.width(width)) rd_st8_1218  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1218]), .rdlo_in(a8_wr[1222]),  .coef_in(coef[512]), .rdup_out(a9_wr[1218]), .rdlo_out(a9_wr[1222]));
			radix2 #(.width(width)) rd_st8_1219  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1219]), .rdlo_in(a8_wr[1223]),  .coef_in(coef[768]), .rdup_out(a9_wr[1219]), .rdlo_out(a9_wr[1223]));
			radix2 #(.width(width)) rd_st8_1224  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1224]), .rdlo_in(a8_wr[1228]),  .coef_in(coef[0]), .rdup_out(a9_wr[1224]), .rdlo_out(a9_wr[1228]));
			radix2 #(.width(width)) rd_st8_1225  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1225]), .rdlo_in(a8_wr[1229]),  .coef_in(coef[256]), .rdup_out(a9_wr[1225]), .rdlo_out(a9_wr[1229]));
			radix2 #(.width(width)) rd_st8_1226  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1226]), .rdlo_in(a8_wr[1230]),  .coef_in(coef[512]), .rdup_out(a9_wr[1226]), .rdlo_out(a9_wr[1230]));
			radix2 #(.width(width)) rd_st8_1227  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1227]), .rdlo_in(a8_wr[1231]),  .coef_in(coef[768]), .rdup_out(a9_wr[1227]), .rdlo_out(a9_wr[1231]));
			radix2 #(.width(width)) rd_st8_1232  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1232]), .rdlo_in(a8_wr[1236]),  .coef_in(coef[0]), .rdup_out(a9_wr[1232]), .rdlo_out(a9_wr[1236]));
			radix2 #(.width(width)) rd_st8_1233  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1233]), .rdlo_in(a8_wr[1237]),  .coef_in(coef[256]), .rdup_out(a9_wr[1233]), .rdlo_out(a9_wr[1237]));
			radix2 #(.width(width)) rd_st8_1234  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1234]), .rdlo_in(a8_wr[1238]),  .coef_in(coef[512]), .rdup_out(a9_wr[1234]), .rdlo_out(a9_wr[1238]));
			radix2 #(.width(width)) rd_st8_1235  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1235]), .rdlo_in(a8_wr[1239]),  .coef_in(coef[768]), .rdup_out(a9_wr[1235]), .rdlo_out(a9_wr[1239]));
			radix2 #(.width(width)) rd_st8_1240  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1240]), .rdlo_in(a8_wr[1244]),  .coef_in(coef[0]), .rdup_out(a9_wr[1240]), .rdlo_out(a9_wr[1244]));
			radix2 #(.width(width)) rd_st8_1241  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1241]), .rdlo_in(a8_wr[1245]),  .coef_in(coef[256]), .rdup_out(a9_wr[1241]), .rdlo_out(a9_wr[1245]));
			radix2 #(.width(width)) rd_st8_1242  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1242]), .rdlo_in(a8_wr[1246]),  .coef_in(coef[512]), .rdup_out(a9_wr[1242]), .rdlo_out(a9_wr[1246]));
			radix2 #(.width(width)) rd_st8_1243  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1243]), .rdlo_in(a8_wr[1247]),  .coef_in(coef[768]), .rdup_out(a9_wr[1243]), .rdlo_out(a9_wr[1247]));
			radix2 #(.width(width)) rd_st8_1248  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1248]), .rdlo_in(a8_wr[1252]),  .coef_in(coef[0]), .rdup_out(a9_wr[1248]), .rdlo_out(a9_wr[1252]));
			radix2 #(.width(width)) rd_st8_1249  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1249]), .rdlo_in(a8_wr[1253]),  .coef_in(coef[256]), .rdup_out(a9_wr[1249]), .rdlo_out(a9_wr[1253]));
			radix2 #(.width(width)) rd_st8_1250  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1250]), .rdlo_in(a8_wr[1254]),  .coef_in(coef[512]), .rdup_out(a9_wr[1250]), .rdlo_out(a9_wr[1254]));
			radix2 #(.width(width)) rd_st8_1251  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1251]), .rdlo_in(a8_wr[1255]),  .coef_in(coef[768]), .rdup_out(a9_wr[1251]), .rdlo_out(a9_wr[1255]));
			radix2 #(.width(width)) rd_st8_1256  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1256]), .rdlo_in(a8_wr[1260]),  .coef_in(coef[0]), .rdup_out(a9_wr[1256]), .rdlo_out(a9_wr[1260]));
			radix2 #(.width(width)) rd_st8_1257  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1257]), .rdlo_in(a8_wr[1261]),  .coef_in(coef[256]), .rdup_out(a9_wr[1257]), .rdlo_out(a9_wr[1261]));
			radix2 #(.width(width)) rd_st8_1258  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1258]), .rdlo_in(a8_wr[1262]),  .coef_in(coef[512]), .rdup_out(a9_wr[1258]), .rdlo_out(a9_wr[1262]));
			radix2 #(.width(width)) rd_st8_1259  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1259]), .rdlo_in(a8_wr[1263]),  .coef_in(coef[768]), .rdup_out(a9_wr[1259]), .rdlo_out(a9_wr[1263]));
			radix2 #(.width(width)) rd_st8_1264  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1264]), .rdlo_in(a8_wr[1268]),  .coef_in(coef[0]), .rdup_out(a9_wr[1264]), .rdlo_out(a9_wr[1268]));
			radix2 #(.width(width)) rd_st8_1265  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1265]), .rdlo_in(a8_wr[1269]),  .coef_in(coef[256]), .rdup_out(a9_wr[1265]), .rdlo_out(a9_wr[1269]));
			radix2 #(.width(width)) rd_st8_1266  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1266]), .rdlo_in(a8_wr[1270]),  .coef_in(coef[512]), .rdup_out(a9_wr[1266]), .rdlo_out(a9_wr[1270]));
			radix2 #(.width(width)) rd_st8_1267  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1267]), .rdlo_in(a8_wr[1271]),  .coef_in(coef[768]), .rdup_out(a9_wr[1267]), .rdlo_out(a9_wr[1271]));
			radix2 #(.width(width)) rd_st8_1272  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1272]), .rdlo_in(a8_wr[1276]),  .coef_in(coef[0]), .rdup_out(a9_wr[1272]), .rdlo_out(a9_wr[1276]));
			radix2 #(.width(width)) rd_st8_1273  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1273]), .rdlo_in(a8_wr[1277]),  .coef_in(coef[256]), .rdup_out(a9_wr[1273]), .rdlo_out(a9_wr[1277]));
			radix2 #(.width(width)) rd_st8_1274  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1274]), .rdlo_in(a8_wr[1278]),  .coef_in(coef[512]), .rdup_out(a9_wr[1274]), .rdlo_out(a9_wr[1278]));
			radix2 #(.width(width)) rd_st8_1275  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1275]), .rdlo_in(a8_wr[1279]),  .coef_in(coef[768]), .rdup_out(a9_wr[1275]), .rdlo_out(a9_wr[1279]));
			radix2 #(.width(width)) rd_st8_1280  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1280]), .rdlo_in(a8_wr[1284]),  .coef_in(coef[0]), .rdup_out(a9_wr[1280]), .rdlo_out(a9_wr[1284]));
			radix2 #(.width(width)) rd_st8_1281  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1281]), .rdlo_in(a8_wr[1285]),  .coef_in(coef[256]), .rdup_out(a9_wr[1281]), .rdlo_out(a9_wr[1285]));
			radix2 #(.width(width)) rd_st8_1282  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1282]), .rdlo_in(a8_wr[1286]),  .coef_in(coef[512]), .rdup_out(a9_wr[1282]), .rdlo_out(a9_wr[1286]));
			radix2 #(.width(width)) rd_st8_1283  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1283]), .rdlo_in(a8_wr[1287]),  .coef_in(coef[768]), .rdup_out(a9_wr[1283]), .rdlo_out(a9_wr[1287]));
			radix2 #(.width(width)) rd_st8_1288  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1288]), .rdlo_in(a8_wr[1292]),  .coef_in(coef[0]), .rdup_out(a9_wr[1288]), .rdlo_out(a9_wr[1292]));
			radix2 #(.width(width)) rd_st8_1289  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1289]), .rdlo_in(a8_wr[1293]),  .coef_in(coef[256]), .rdup_out(a9_wr[1289]), .rdlo_out(a9_wr[1293]));
			radix2 #(.width(width)) rd_st8_1290  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1290]), .rdlo_in(a8_wr[1294]),  .coef_in(coef[512]), .rdup_out(a9_wr[1290]), .rdlo_out(a9_wr[1294]));
			radix2 #(.width(width)) rd_st8_1291  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1291]), .rdlo_in(a8_wr[1295]),  .coef_in(coef[768]), .rdup_out(a9_wr[1291]), .rdlo_out(a9_wr[1295]));
			radix2 #(.width(width)) rd_st8_1296  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1296]), .rdlo_in(a8_wr[1300]),  .coef_in(coef[0]), .rdup_out(a9_wr[1296]), .rdlo_out(a9_wr[1300]));
			radix2 #(.width(width)) rd_st8_1297  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1297]), .rdlo_in(a8_wr[1301]),  .coef_in(coef[256]), .rdup_out(a9_wr[1297]), .rdlo_out(a9_wr[1301]));
			radix2 #(.width(width)) rd_st8_1298  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1298]), .rdlo_in(a8_wr[1302]),  .coef_in(coef[512]), .rdup_out(a9_wr[1298]), .rdlo_out(a9_wr[1302]));
			radix2 #(.width(width)) rd_st8_1299  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1299]), .rdlo_in(a8_wr[1303]),  .coef_in(coef[768]), .rdup_out(a9_wr[1299]), .rdlo_out(a9_wr[1303]));
			radix2 #(.width(width)) rd_st8_1304  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1304]), .rdlo_in(a8_wr[1308]),  .coef_in(coef[0]), .rdup_out(a9_wr[1304]), .rdlo_out(a9_wr[1308]));
			radix2 #(.width(width)) rd_st8_1305  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1305]), .rdlo_in(a8_wr[1309]),  .coef_in(coef[256]), .rdup_out(a9_wr[1305]), .rdlo_out(a9_wr[1309]));
			radix2 #(.width(width)) rd_st8_1306  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1306]), .rdlo_in(a8_wr[1310]),  .coef_in(coef[512]), .rdup_out(a9_wr[1306]), .rdlo_out(a9_wr[1310]));
			radix2 #(.width(width)) rd_st8_1307  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1307]), .rdlo_in(a8_wr[1311]),  .coef_in(coef[768]), .rdup_out(a9_wr[1307]), .rdlo_out(a9_wr[1311]));
			radix2 #(.width(width)) rd_st8_1312  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1312]), .rdlo_in(a8_wr[1316]),  .coef_in(coef[0]), .rdup_out(a9_wr[1312]), .rdlo_out(a9_wr[1316]));
			radix2 #(.width(width)) rd_st8_1313  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1313]), .rdlo_in(a8_wr[1317]),  .coef_in(coef[256]), .rdup_out(a9_wr[1313]), .rdlo_out(a9_wr[1317]));
			radix2 #(.width(width)) rd_st8_1314  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1314]), .rdlo_in(a8_wr[1318]),  .coef_in(coef[512]), .rdup_out(a9_wr[1314]), .rdlo_out(a9_wr[1318]));
			radix2 #(.width(width)) rd_st8_1315  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1315]), .rdlo_in(a8_wr[1319]),  .coef_in(coef[768]), .rdup_out(a9_wr[1315]), .rdlo_out(a9_wr[1319]));
			radix2 #(.width(width)) rd_st8_1320  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1320]), .rdlo_in(a8_wr[1324]),  .coef_in(coef[0]), .rdup_out(a9_wr[1320]), .rdlo_out(a9_wr[1324]));
			radix2 #(.width(width)) rd_st8_1321  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1321]), .rdlo_in(a8_wr[1325]),  .coef_in(coef[256]), .rdup_out(a9_wr[1321]), .rdlo_out(a9_wr[1325]));
			radix2 #(.width(width)) rd_st8_1322  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1322]), .rdlo_in(a8_wr[1326]),  .coef_in(coef[512]), .rdup_out(a9_wr[1322]), .rdlo_out(a9_wr[1326]));
			radix2 #(.width(width)) rd_st8_1323  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1323]), .rdlo_in(a8_wr[1327]),  .coef_in(coef[768]), .rdup_out(a9_wr[1323]), .rdlo_out(a9_wr[1327]));
			radix2 #(.width(width)) rd_st8_1328  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1328]), .rdlo_in(a8_wr[1332]),  .coef_in(coef[0]), .rdup_out(a9_wr[1328]), .rdlo_out(a9_wr[1332]));
			radix2 #(.width(width)) rd_st8_1329  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1329]), .rdlo_in(a8_wr[1333]),  .coef_in(coef[256]), .rdup_out(a9_wr[1329]), .rdlo_out(a9_wr[1333]));
			radix2 #(.width(width)) rd_st8_1330  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1330]), .rdlo_in(a8_wr[1334]),  .coef_in(coef[512]), .rdup_out(a9_wr[1330]), .rdlo_out(a9_wr[1334]));
			radix2 #(.width(width)) rd_st8_1331  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1331]), .rdlo_in(a8_wr[1335]),  .coef_in(coef[768]), .rdup_out(a9_wr[1331]), .rdlo_out(a9_wr[1335]));
			radix2 #(.width(width)) rd_st8_1336  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1336]), .rdlo_in(a8_wr[1340]),  .coef_in(coef[0]), .rdup_out(a9_wr[1336]), .rdlo_out(a9_wr[1340]));
			radix2 #(.width(width)) rd_st8_1337  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1337]), .rdlo_in(a8_wr[1341]),  .coef_in(coef[256]), .rdup_out(a9_wr[1337]), .rdlo_out(a9_wr[1341]));
			radix2 #(.width(width)) rd_st8_1338  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1338]), .rdlo_in(a8_wr[1342]),  .coef_in(coef[512]), .rdup_out(a9_wr[1338]), .rdlo_out(a9_wr[1342]));
			radix2 #(.width(width)) rd_st8_1339  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1339]), .rdlo_in(a8_wr[1343]),  .coef_in(coef[768]), .rdup_out(a9_wr[1339]), .rdlo_out(a9_wr[1343]));
			radix2 #(.width(width)) rd_st8_1344  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1344]), .rdlo_in(a8_wr[1348]),  .coef_in(coef[0]), .rdup_out(a9_wr[1344]), .rdlo_out(a9_wr[1348]));
			radix2 #(.width(width)) rd_st8_1345  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1345]), .rdlo_in(a8_wr[1349]),  .coef_in(coef[256]), .rdup_out(a9_wr[1345]), .rdlo_out(a9_wr[1349]));
			radix2 #(.width(width)) rd_st8_1346  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1346]), .rdlo_in(a8_wr[1350]),  .coef_in(coef[512]), .rdup_out(a9_wr[1346]), .rdlo_out(a9_wr[1350]));
			radix2 #(.width(width)) rd_st8_1347  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1347]), .rdlo_in(a8_wr[1351]),  .coef_in(coef[768]), .rdup_out(a9_wr[1347]), .rdlo_out(a9_wr[1351]));
			radix2 #(.width(width)) rd_st8_1352  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1352]), .rdlo_in(a8_wr[1356]),  .coef_in(coef[0]), .rdup_out(a9_wr[1352]), .rdlo_out(a9_wr[1356]));
			radix2 #(.width(width)) rd_st8_1353  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1353]), .rdlo_in(a8_wr[1357]),  .coef_in(coef[256]), .rdup_out(a9_wr[1353]), .rdlo_out(a9_wr[1357]));
			radix2 #(.width(width)) rd_st8_1354  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1354]), .rdlo_in(a8_wr[1358]),  .coef_in(coef[512]), .rdup_out(a9_wr[1354]), .rdlo_out(a9_wr[1358]));
			radix2 #(.width(width)) rd_st8_1355  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1355]), .rdlo_in(a8_wr[1359]),  .coef_in(coef[768]), .rdup_out(a9_wr[1355]), .rdlo_out(a9_wr[1359]));
			radix2 #(.width(width)) rd_st8_1360  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1360]), .rdlo_in(a8_wr[1364]),  .coef_in(coef[0]), .rdup_out(a9_wr[1360]), .rdlo_out(a9_wr[1364]));
			radix2 #(.width(width)) rd_st8_1361  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1361]), .rdlo_in(a8_wr[1365]),  .coef_in(coef[256]), .rdup_out(a9_wr[1361]), .rdlo_out(a9_wr[1365]));
			radix2 #(.width(width)) rd_st8_1362  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1362]), .rdlo_in(a8_wr[1366]),  .coef_in(coef[512]), .rdup_out(a9_wr[1362]), .rdlo_out(a9_wr[1366]));
			radix2 #(.width(width)) rd_st8_1363  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1363]), .rdlo_in(a8_wr[1367]),  .coef_in(coef[768]), .rdup_out(a9_wr[1363]), .rdlo_out(a9_wr[1367]));
			radix2 #(.width(width)) rd_st8_1368  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1368]), .rdlo_in(a8_wr[1372]),  .coef_in(coef[0]), .rdup_out(a9_wr[1368]), .rdlo_out(a9_wr[1372]));
			radix2 #(.width(width)) rd_st8_1369  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1369]), .rdlo_in(a8_wr[1373]),  .coef_in(coef[256]), .rdup_out(a9_wr[1369]), .rdlo_out(a9_wr[1373]));
			radix2 #(.width(width)) rd_st8_1370  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1370]), .rdlo_in(a8_wr[1374]),  .coef_in(coef[512]), .rdup_out(a9_wr[1370]), .rdlo_out(a9_wr[1374]));
			radix2 #(.width(width)) rd_st8_1371  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1371]), .rdlo_in(a8_wr[1375]),  .coef_in(coef[768]), .rdup_out(a9_wr[1371]), .rdlo_out(a9_wr[1375]));
			radix2 #(.width(width)) rd_st8_1376  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1376]), .rdlo_in(a8_wr[1380]),  .coef_in(coef[0]), .rdup_out(a9_wr[1376]), .rdlo_out(a9_wr[1380]));
			radix2 #(.width(width)) rd_st8_1377  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1377]), .rdlo_in(a8_wr[1381]),  .coef_in(coef[256]), .rdup_out(a9_wr[1377]), .rdlo_out(a9_wr[1381]));
			radix2 #(.width(width)) rd_st8_1378  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1378]), .rdlo_in(a8_wr[1382]),  .coef_in(coef[512]), .rdup_out(a9_wr[1378]), .rdlo_out(a9_wr[1382]));
			radix2 #(.width(width)) rd_st8_1379  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1379]), .rdlo_in(a8_wr[1383]),  .coef_in(coef[768]), .rdup_out(a9_wr[1379]), .rdlo_out(a9_wr[1383]));
			radix2 #(.width(width)) rd_st8_1384  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1384]), .rdlo_in(a8_wr[1388]),  .coef_in(coef[0]), .rdup_out(a9_wr[1384]), .rdlo_out(a9_wr[1388]));
			radix2 #(.width(width)) rd_st8_1385  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1385]), .rdlo_in(a8_wr[1389]),  .coef_in(coef[256]), .rdup_out(a9_wr[1385]), .rdlo_out(a9_wr[1389]));
			radix2 #(.width(width)) rd_st8_1386  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1386]), .rdlo_in(a8_wr[1390]),  .coef_in(coef[512]), .rdup_out(a9_wr[1386]), .rdlo_out(a9_wr[1390]));
			radix2 #(.width(width)) rd_st8_1387  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1387]), .rdlo_in(a8_wr[1391]),  .coef_in(coef[768]), .rdup_out(a9_wr[1387]), .rdlo_out(a9_wr[1391]));
			radix2 #(.width(width)) rd_st8_1392  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1392]), .rdlo_in(a8_wr[1396]),  .coef_in(coef[0]), .rdup_out(a9_wr[1392]), .rdlo_out(a9_wr[1396]));
			radix2 #(.width(width)) rd_st8_1393  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1393]), .rdlo_in(a8_wr[1397]),  .coef_in(coef[256]), .rdup_out(a9_wr[1393]), .rdlo_out(a9_wr[1397]));
			radix2 #(.width(width)) rd_st8_1394  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1394]), .rdlo_in(a8_wr[1398]),  .coef_in(coef[512]), .rdup_out(a9_wr[1394]), .rdlo_out(a9_wr[1398]));
			radix2 #(.width(width)) rd_st8_1395  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1395]), .rdlo_in(a8_wr[1399]),  .coef_in(coef[768]), .rdup_out(a9_wr[1395]), .rdlo_out(a9_wr[1399]));
			radix2 #(.width(width)) rd_st8_1400  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1400]), .rdlo_in(a8_wr[1404]),  .coef_in(coef[0]), .rdup_out(a9_wr[1400]), .rdlo_out(a9_wr[1404]));
			radix2 #(.width(width)) rd_st8_1401  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1401]), .rdlo_in(a8_wr[1405]),  .coef_in(coef[256]), .rdup_out(a9_wr[1401]), .rdlo_out(a9_wr[1405]));
			radix2 #(.width(width)) rd_st8_1402  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1402]), .rdlo_in(a8_wr[1406]),  .coef_in(coef[512]), .rdup_out(a9_wr[1402]), .rdlo_out(a9_wr[1406]));
			radix2 #(.width(width)) rd_st8_1403  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1403]), .rdlo_in(a8_wr[1407]),  .coef_in(coef[768]), .rdup_out(a9_wr[1403]), .rdlo_out(a9_wr[1407]));
			radix2 #(.width(width)) rd_st8_1408  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1408]), .rdlo_in(a8_wr[1412]),  .coef_in(coef[0]), .rdup_out(a9_wr[1408]), .rdlo_out(a9_wr[1412]));
			radix2 #(.width(width)) rd_st8_1409  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1409]), .rdlo_in(a8_wr[1413]),  .coef_in(coef[256]), .rdup_out(a9_wr[1409]), .rdlo_out(a9_wr[1413]));
			radix2 #(.width(width)) rd_st8_1410  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1410]), .rdlo_in(a8_wr[1414]),  .coef_in(coef[512]), .rdup_out(a9_wr[1410]), .rdlo_out(a9_wr[1414]));
			radix2 #(.width(width)) rd_st8_1411  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1411]), .rdlo_in(a8_wr[1415]),  .coef_in(coef[768]), .rdup_out(a9_wr[1411]), .rdlo_out(a9_wr[1415]));
			radix2 #(.width(width)) rd_st8_1416  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1416]), .rdlo_in(a8_wr[1420]),  .coef_in(coef[0]), .rdup_out(a9_wr[1416]), .rdlo_out(a9_wr[1420]));
			radix2 #(.width(width)) rd_st8_1417  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1417]), .rdlo_in(a8_wr[1421]),  .coef_in(coef[256]), .rdup_out(a9_wr[1417]), .rdlo_out(a9_wr[1421]));
			radix2 #(.width(width)) rd_st8_1418  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1418]), .rdlo_in(a8_wr[1422]),  .coef_in(coef[512]), .rdup_out(a9_wr[1418]), .rdlo_out(a9_wr[1422]));
			radix2 #(.width(width)) rd_st8_1419  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1419]), .rdlo_in(a8_wr[1423]),  .coef_in(coef[768]), .rdup_out(a9_wr[1419]), .rdlo_out(a9_wr[1423]));
			radix2 #(.width(width)) rd_st8_1424  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1424]), .rdlo_in(a8_wr[1428]),  .coef_in(coef[0]), .rdup_out(a9_wr[1424]), .rdlo_out(a9_wr[1428]));
			radix2 #(.width(width)) rd_st8_1425  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1425]), .rdlo_in(a8_wr[1429]),  .coef_in(coef[256]), .rdup_out(a9_wr[1425]), .rdlo_out(a9_wr[1429]));
			radix2 #(.width(width)) rd_st8_1426  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1426]), .rdlo_in(a8_wr[1430]),  .coef_in(coef[512]), .rdup_out(a9_wr[1426]), .rdlo_out(a9_wr[1430]));
			radix2 #(.width(width)) rd_st8_1427  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1427]), .rdlo_in(a8_wr[1431]),  .coef_in(coef[768]), .rdup_out(a9_wr[1427]), .rdlo_out(a9_wr[1431]));
			radix2 #(.width(width)) rd_st8_1432  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1432]), .rdlo_in(a8_wr[1436]),  .coef_in(coef[0]), .rdup_out(a9_wr[1432]), .rdlo_out(a9_wr[1436]));
			radix2 #(.width(width)) rd_st8_1433  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1433]), .rdlo_in(a8_wr[1437]),  .coef_in(coef[256]), .rdup_out(a9_wr[1433]), .rdlo_out(a9_wr[1437]));
			radix2 #(.width(width)) rd_st8_1434  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1434]), .rdlo_in(a8_wr[1438]),  .coef_in(coef[512]), .rdup_out(a9_wr[1434]), .rdlo_out(a9_wr[1438]));
			radix2 #(.width(width)) rd_st8_1435  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1435]), .rdlo_in(a8_wr[1439]),  .coef_in(coef[768]), .rdup_out(a9_wr[1435]), .rdlo_out(a9_wr[1439]));
			radix2 #(.width(width)) rd_st8_1440  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1440]), .rdlo_in(a8_wr[1444]),  .coef_in(coef[0]), .rdup_out(a9_wr[1440]), .rdlo_out(a9_wr[1444]));
			radix2 #(.width(width)) rd_st8_1441  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1441]), .rdlo_in(a8_wr[1445]),  .coef_in(coef[256]), .rdup_out(a9_wr[1441]), .rdlo_out(a9_wr[1445]));
			radix2 #(.width(width)) rd_st8_1442  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1442]), .rdlo_in(a8_wr[1446]),  .coef_in(coef[512]), .rdup_out(a9_wr[1442]), .rdlo_out(a9_wr[1446]));
			radix2 #(.width(width)) rd_st8_1443  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1443]), .rdlo_in(a8_wr[1447]),  .coef_in(coef[768]), .rdup_out(a9_wr[1443]), .rdlo_out(a9_wr[1447]));
			radix2 #(.width(width)) rd_st8_1448  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1448]), .rdlo_in(a8_wr[1452]),  .coef_in(coef[0]), .rdup_out(a9_wr[1448]), .rdlo_out(a9_wr[1452]));
			radix2 #(.width(width)) rd_st8_1449  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1449]), .rdlo_in(a8_wr[1453]),  .coef_in(coef[256]), .rdup_out(a9_wr[1449]), .rdlo_out(a9_wr[1453]));
			radix2 #(.width(width)) rd_st8_1450  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1450]), .rdlo_in(a8_wr[1454]),  .coef_in(coef[512]), .rdup_out(a9_wr[1450]), .rdlo_out(a9_wr[1454]));
			radix2 #(.width(width)) rd_st8_1451  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1451]), .rdlo_in(a8_wr[1455]),  .coef_in(coef[768]), .rdup_out(a9_wr[1451]), .rdlo_out(a9_wr[1455]));
			radix2 #(.width(width)) rd_st8_1456  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1456]), .rdlo_in(a8_wr[1460]),  .coef_in(coef[0]), .rdup_out(a9_wr[1456]), .rdlo_out(a9_wr[1460]));
			radix2 #(.width(width)) rd_st8_1457  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1457]), .rdlo_in(a8_wr[1461]),  .coef_in(coef[256]), .rdup_out(a9_wr[1457]), .rdlo_out(a9_wr[1461]));
			radix2 #(.width(width)) rd_st8_1458  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1458]), .rdlo_in(a8_wr[1462]),  .coef_in(coef[512]), .rdup_out(a9_wr[1458]), .rdlo_out(a9_wr[1462]));
			radix2 #(.width(width)) rd_st8_1459  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1459]), .rdlo_in(a8_wr[1463]),  .coef_in(coef[768]), .rdup_out(a9_wr[1459]), .rdlo_out(a9_wr[1463]));
			radix2 #(.width(width)) rd_st8_1464  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1464]), .rdlo_in(a8_wr[1468]),  .coef_in(coef[0]), .rdup_out(a9_wr[1464]), .rdlo_out(a9_wr[1468]));
			radix2 #(.width(width)) rd_st8_1465  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1465]), .rdlo_in(a8_wr[1469]),  .coef_in(coef[256]), .rdup_out(a9_wr[1465]), .rdlo_out(a9_wr[1469]));
			radix2 #(.width(width)) rd_st8_1466  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1466]), .rdlo_in(a8_wr[1470]),  .coef_in(coef[512]), .rdup_out(a9_wr[1466]), .rdlo_out(a9_wr[1470]));
			radix2 #(.width(width)) rd_st8_1467  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1467]), .rdlo_in(a8_wr[1471]),  .coef_in(coef[768]), .rdup_out(a9_wr[1467]), .rdlo_out(a9_wr[1471]));
			radix2 #(.width(width)) rd_st8_1472  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1472]), .rdlo_in(a8_wr[1476]),  .coef_in(coef[0]), .rdup_out(a9_wr[1472]), .rdlo_out(a9_wr[1476]));
			radix2 #(.width(width)) rd_st8_1473  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1473]), .rdlo_in(a8_wr[1477]),  .coef_in(coef[256]), .rdup_out(a9_wr[1473]), .rdlo_out(a9_wr[1477]));
			radix2 #(.width(width)) rd_st8_1474  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1474]), .rdlo_in(a8_wr[1478]),  .coef_in(coef[512]), .rdup_out(a9_wr[1474]), .rdlo_out(a9_wr[1478]));
			radix2 #(.width(width)) rd_st8_1475  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1475]), .rdlo_in(a8_wr[1479]),  .coef_in(coef[768]), .rdup_out(a9_wr[1475]), .rdlo_out(a9_wr[1479]));
			radix2 #(.width(width)) rd_st8_1480  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1480]), .rdlo_in(a8_wr[1484]),  .coef_in(coef[0]), .rdup_out(a9_wr[1480]), .rdlo_out(a9_wr[1484]));
			radix2 #(.width(width)) rd_st8_1481  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1481]), .rdlo_in(a8_wr[1485]),  .coef_in(coef[256]), .rdup_out(a9_wr[1481]), .rdlo_out(a9_wr[1485]));
			radix2 #(.width(width)) rd_st8_1482  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1482]), .rdlo_in(a8_wr[1486]),  .coef_in(coef[512]), .rdup_out(a9_wr[1482]), .rdlo_out(a9_wr[1486]));
			radix2 #(.width(width)) rd_st8_1483  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1483]), .rdlo_in(a8_wr[1487]),  .coef_in(coef[768]), .rdup_out(a9_wr[1483]), .rdlo_out(a9_wr[1487]));
			radix2 #(.width(width)) rd_st8_1488  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1488]), .rdlo_in(a8_wr[1492]),  .coef_in(coef[0]), .rdup_out(a9_wr[1488]), .rdlo_out(a9_wr[1492]));
			radix2 #(.width(width)) rd_st8_1489  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1489]), .rdlo_in(a8_wr[1493]),  .coef_in(coef[256]), .rdup_out(a9_wr[1489]), .rdlo_out(a9_wr[1493]));
			radix2 #(.width(width)) rd_st8_1490  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1490]), .rdlo_in(a8_wr[1494]),  .coef_in(coef[512]), .rdup_out(a9_wr[1490]), .rdlo_out(a9_wr[1494]));
			radix2 #(.width(width)) rd_st8_1491  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1491]), .rdlo_in(a8_wr[1495]),  .coef_in(coef[768]), .rdup_out(a9_wr[1491]), .rdlo_out(a9_wr[1495]));
			radix2 #(.width(width)) rd_st8_1496  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1496]), .rdlo_in(a8_wr[1500]),  .coef_in(coef[0]), .rdup_out(a9_wr[1496]), .rdlo_out(a9_wr[1500]));
			radix2 #(.width(width)) rd_st8_1497  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1497]), .rdlo_in(a8_wr[1501]),  .coef_in(coef[256]), .rdup_out(a9_wr[1497]), .rdlo_out(a9_wr[1501]));
			radix2 #(.width(width)) rd_st8_1498  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1498]), .rdlo_in(a8_wr[1502]),  .coef_in(coef[512]), .rdup_out(a9_wr[1498]), .rdlo_out(a9_wr[1502]));
			radix2 #(.width(width)) rd_st8_1499  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1499]), .rdlo_in(a8_wr[1503]),  .coef_in(coef[768]), .rdup_out(a9_wr[1499]), .rdlo_out(a9_wr[1503]));
			radix2 #(.width(width)) rd_st8_1504  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1504]), .rdlo_in(a8_wr[1508]),  .coef_in(coef[0]), .rdup_out(a9_wr[1504]), .rdlo_out(a9_wr[1508]));
			radix2 #(.width(width)) rd_st8_1505  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1505]), .rdlo_in(a8_wr[1509]),  .coef_in(coef[256]), .rdup_out(a9_wr[1505]), .rdlo_out(a9_wr[1509]));
			radix2 #(.width(width)) rd_st8_1506  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1506]), .rdlo_in(a8_wr[1510]),  .coef_in(coef[512]), .rdup_out(a9_wr[1506]), .rdlo_out(a9_wr[1510]));
			radix2 #(.width(width)) rd_st8_1507  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1507]), .rdlo_in(a8_wr[1511]),  .coef_in(coef[768]), .rdup_out(a9_wr[1507]), .rdlo_out(a9_wr[1511]));
			radix2 #(.width(width)) rd_st8_1512  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1512]), .rdlo_in(a8_wr[1516]),  .coef_in(coef[0]), .rdup_out(a9_wr[1512]), .rdlo_out(a9_wr[1516]));
			radix2 #(.width(width)) rd_st8_1513  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1513]), .rdlo_in(a8_wr[1517]),  .coef_in(coef[256]), .rdup_out(a9_wr[1513]), .rdlo_out(a9_wr[1517]));
			radix2 #(.width(width)) rd_st8_1514  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1514]), .rdlo_in(a8_wr[1518]),  .coef_in(coef[512]), .rdup_out(a9_wr[1514]), .rdlo_out(a9_wr[1518]));
			radix2 #(.width(width)) rd_st8_1515  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1515]), .rdlo_in(a8_wr[1519]),  .coef_in(coef[768]), .rdup_out(a9_wr[1515]), .rdlo_out(a9_wr[1519]));
			radix2 #(.width(width)) rd_st8_1520  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1520]), .rdlo_in(a8_wr[1524]),  .coef_in(coef[0]), .rdup_out(a9_wr[1520]), .rdlo_out(a9_wr[1524]));
			radix2 #(.width(width)) rd_st8_1521  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1521]), .rdlo_in(a8_wr[1525]),  .coef_in(coef[256]), .rdup_out(a9_wr[1521]), .rdlo_out(a9_wr[1525]));
			radix2 #(.width(width)) rd_st8_1522  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1522]), .rdlo_in(a8_wr[1526]),  .coef_in(coef[512]), .rdup_out(a9_wr[1522]), .rdlo_out(a9_wr[1526]));
			radix2 #(.width(width)) rd_st8_1523  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1523]), .rdlo_in(a8_wr[1527]),  .coef_in(coef[768]), .rdup_out(a9_wr[1523]), .rdlo_out(a9_wr[1527]));
			radix2 #(.width(width)) rd_st8_1528  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1528]), .rdlo_in(a8_wr[1532]),  .coef_in(coef[0]), .rdup_out(a9_wr[1528]), .rdlo_out(a9_wr[1532]));
			radix2 #(.width(width)) rd_st8_1529  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1529]), .rdlo_in(a8_wr[1533]),  .coef_in(coef[256]), .rdup_out(a9_wr[1529]), .rdlo_out(a9_wr[1533]));
			radix2 #(.width(width)) rd_st8_1530  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1530]), .rdlo_in(a8_wr[1534]),  .coef_in(coef[512]), .rdup_out(a9_wr[1530]), .rdlo_out(a9_wr[1534]));
			radix2 #(.width(width)) rd_st8_1531  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1531]), .rdlo_in(a8_wr[1535]),  .coef_in(coef[768]), .rdup_out(a9_wr[1531]), .rdlo_out(a9_wr[1535]));
			radix2 #(.width(width)) rd_st8_1536  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1536]), .rdlo_in(a8_wr[1540]),  .coef_in(coef[0]), .rdup_out(a9_wr[1536]), .rdlo_out(a9_wr[1540]));
			radix2 #(.width(width)) rd_st8_1537  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1537]), .rdlo_in(a8_wr[1541]),  .coef_in(coef[256]), .rdup_out(a9_wr[1537]), .rdlo_out(a9_wr[1541]));
			radix2 #(.width(width)) rd_st8_1538  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1538]), .rdlo_in(a8_wr[1542]),  .coef_in(coef[512]), .rdup_out(a9_wr[1538]), .rdlo_out(a9_wr[1542]));
			radix2 #(.width(width)) rd_st8_1539  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1539]), .rdlo_in(a8_wr[1543]),  .coef_in(coef[768]), .rdup_out(a9_wr[1539]), .rdlo_out(a9_wr[1543]));
			radix2 #(.width(width)) rd_st8_1544  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1544]), .rdlo_in(a8_wr[1548]),  .coef_in(coef[0]), .rdup_out(a9_wr[1544]), .rdlo_out(a9_wr[1548]));
			radix2 #(.width(width)) rd_st8_1545  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1545]), .rdlo_in(a8_wr[1549]),  .coef_in(coef[256]), .rdup_out(a9_wr[1545]), .rdlo_out(a9_wr[1549]));
			radix2 #(.width(width)) rd_st8_1546  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1546]), .rdlo_in(a8_wr[1550]),  .coef_in(coef[512]), .rdup_out(a9_wr[1546]), .rdlo_out(a9_wr[1550]));
			radix2 #(.width(width)) rd_st8_1547  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1547]), .rdlo_in(a8_wr[1551]),  .coef_in(coef[768]), .rdup_out(a9_wr[1547]), .rdlo_out(a9_wr[1551]));
			radix2 #(.width(width)) rd_st8_1552  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1552]), .rdlo_in(a8_wr[1556]),  .coef_in(coef[0]), .rdup_out(a9_wr[1552]), .rdlo_out(a9_wr[1556]));
			radix2 #(.width(width)) rd_st8_1553  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1553]), .rdlo_in(a8_wr[1557]),  .coef_in(coef[256]), .rdup_out(a9_wr[1553]), .rdlo_out(a9_wr[1557]));
			radix2 #(.width(width)) rd_st8_1554  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1554]), .rdlo_in(a8_wr[1558]),  .coef_in(coef[512]), .rdup_out(a9_wr[1554]), .rdlo_out(a9_wr[1558]));
			radix2 #(.width(width)) rd_st8_1555  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1555]), .rdlo_in(a8_wr[1559]),  .coef_in(coef[768]), .rdup_out(a9_wr[1555]), .rdlo_out(a9_wr[1559]));
			radix2 #(.width(width)) rd_st8_1560  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1560]), .rdlo_in(a8_wr[1564]),  .coef_in(coef[0]), .rdup_out(a9_wr[1560]), .rdlo_out(a9_wr[1564]));
			radix2 #(.width(width)) rd_st8_1561  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1561]), .rdlo_in(a8_wr[1565]),  .coef_in(coef[256]), .rdup_out(a9_wr[1561]), .rdlo_out(a9_wr[1565]));
			radix2 #(.width(width)) rd_st8_1562  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1562]), .rdlo_in(a8_wr[1566]),  .coef_in(coef[512]), .rdup_out(a9_wr[1562]), .rdlo_out(a9_wr[1566]));
			radix2 #(.width(width)) rd_st8_1563  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1563]), .rdlo_in(a8_wr[1567]),  .coef_in(coef[768]), .rdup_out(a9_wr[1563]), .rdlo_out(a9_wr[1567]));
			radix2 #(.width(width)) rd_st8_1568  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1568]), .rdlo_in(a8_wr[1572]),  .coef_in(coef[0]), .rdup_out(a9_wr[1568]), .rdlo_out(a9_wr[1572]));
			radix2 #(.width(width)) rd_st8_1569  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1569]), .rdlo_in(a8_wr[1573]),  .coef_in(coef[256]), .rdup_out(a9_wr[1569]), .rdlo_out(a9_wr[1573]));
			radix2 #(.width(width)) rd_st8_1570  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1570]), .rdlo_in(a8_wr[1574]),  .coef_in(coef[512]), .rdup_out(a9_wr[1570]), .rdlo_out(a9_wr[1574]));
			radix2 #(.width(width)) rd_st8_1571  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1571]), .rdlo_in(a8_wr[1575]),  .coef_in(coef[768]), .rdup_out(a9_wr[1571]), .rdlo_out(a9_wr[1575]));
			radix2 #(.width(width)) rd_st8_1576  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1576]), .rdlo_in(a8_wr[1580]),  .coef_in(coef[0]), .rdup_out(a9_wr[1576]), .rdlo_out(a9_wr[1580]));
			radix2 #(.width(width)) rd_st8_1577  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1577]), .rdlo_in(a8_wr[1581]),  .coef_in(coef[256]), .rdup_out(a9_wr[1577]), .rdlo_out(a9_wr[1581]));
			radix2 #(.width(width)) rd_st8_1578  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1578]), .rdlo_in(a8_wr[1582]),  .coef_in(coef[512]), .rdup_out(a9_wr[1578]), .rdlo_out(a9_wr[1582]));
			radix2 #(.width(width)) rd_st8_1579  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1579]), .rdlo_in(a8_wr[1583]),  .coef_in(coef[768]), .rdup_out(a9_wr[1579]), .rdlo_out(a9_wr[1583]));
			radix2 #(.width(width)) rd_st8_1584  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1584]), .rdlo_in(a8_wr[1588]),  .coef_in(coef[0]), .rdup_out(a9_wr[1584]), .rdlo_out(a9_wr[1588]));
			radix2 #(.width(width)) rd_st8_1585  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1585]), .rdlo_in(a8_wr[1589]),  .coef_in(coef[256]), .rdup_out(a9_wr[1585]), .rdlo_out(a9_wr[1589]));
			radix2 #(.width(width)) rd_st8_1586  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1586]), .rdlo_in(a8_wr[1590]),  .coef_in(coef[512]), .rdup_out(a9_wr[1586]), .rdlo_out(a9_wr[1590]));
			radix2 #(.width(width)) rd_st8_1587  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1587]), .rdlo_in(a8_wr[1591]),  .coef_in(coef[768]), .rdup_out(a9_wr[1587]), .rdlo_out(a9_wr[1591]));
			radix2 #(.width(width)) rd_st8_1592  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1592]), .rdlo_in(a8_wr[1596]),  .coef_in(coef[0]), .rdup_out(a9_wr[1592]), .rdlo_out(a9_wr[1596]));
			radix2 #(.width(width)) rd_st8_1593  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1593]), .rdlo_in(a8_wr[1597]),  .coef_in(coef[256]), .rdup_out(a9_wr[1593]), .rdlo_out(a9_wr[1597]));
			radix2 #(.width(width)) rd_st8_1594  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1594]), .rdlo_in(a8_wr[1598]),  .coef_in(coef[512]), .rdup_out(a9_wr[1594]), .rdlo_out(a9_wr[1598]));
			radix2 #(.width(width)) rd_st8_1595  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1595]), .rdlo_in(a8_wr[1599]),  .coef_in(coef[768]), .rdup_out(a9_wr[1595]), .rdlo_out(a9_wr[1599]));
			radix2 #(.width(width)) rd_st8_1600  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1600]), .rdlo_in(a8_wr[1604]),  .coef_in(coef[0]), .rdup_out(a9_wr[1600]), .rdlo_out(a9_wr[1604]));
			radix2 #(.width(width)) rd_st8_1601  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1601]), .rdlo_in(a8_wr[1605]),  .coef_in(coef[256]), .rdup_out(a9_wr[1601]), .rdlo_out(a9_wr[1605]));
			radix2 #(.width(width)) rd_st8_1602  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1602]), .rdlo_in(a8_wr[1606]),  .coef_in(coef[512]), .rdup_out(a9_wr[1602]), .rdlo_out(a9_wr[1606]));
			radix2 #(.width(width)) rd_st8_1603  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1603]), .rdlo_in(a8_wr[1607]),  .coef_in(coef[768]), .rdup_out(a9_wr[1603]), .rdlo_out(a9_wr[1607]));
			radix2 #(.width(width)) rd_st8_1608  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1608]), .rdlo_in(a8_wr[1612]),  .coef_in(coef[0]), .rdup_out(a9_wr[1608]), .rdlo_out(a9_wr[1612]));
			radix2 #(.width(width)) rd_st8_1609  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1609]), .rdlo_in(a8_wr[1613]),  .coef_in(coef[256]), .rdup_out(a9_wr[1609]), .rdlo_out(a9_wr[1613]));
			radix2 #(.width(width)) rd_st8_1610  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1610]), .rdlo_in(a8_wr[1614]),  .coef_in(coef[512]), .rdup_out(a9_wr[1610]), .rdlo_out(a9_wr[1614]));
			radix2 #(.width(width)) rd_st8_1611  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1611]), .rdlo_in(a8_wr[1615]),  .coef_in(coef[768]), .rdup_out(a9_wr[1611]), .rdlo_out(a9_wr[1615]));
			radix2 #(.width(width)) rd_st8_1616  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1616]), .rdlo_in(a8_wr[1620]),  .coef_in(coef[0]), .rdup_out(a9_wr[1616]), .rdlo_out(a9_wr[1620]));
			radix2 #(.width(width)) rd_st8_1617  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1617]), .rdlo_in(a8_wr[1621]),  .coef_in(coef[256]), .rdup_out(a9_wr[1617]), .rdlo_out(a9_wr[1621]));
			radix2 #(.width(width)) rd_st8_1618  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1618]), .rdlo_in(a8_wr[1622]),  .coef_in(coef[512]), .rdup_out(a9_wr[1618]), .rdlo_out(a9_wr[1622]));
			radix2 #(.width(width)) rd_st8_1619  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1619]), .rdlo_in(a8_wr[1623]),  .coef_in(coef[768]), .rdup_out(a9_wr[1619]), .rdlo_out(a9_wr[1623]));
			radix2 #(.width(width)) rd_st8_1624  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1624]), .rdlo_in(a8_wr[1628]),  .coef_in(coef[0]), .rdup_out(a9_wr[1624]), .rdlo_out(a9_wr[1628]));
			radix2 #(.width(width)) rd_st8_1625  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1625]), .rdlo_in(a8_wr[1629]),  .coef_in(coef[256]), .rdup_out(a9_wr[1625]), .rdlo_out(a9_wr[1629]));
			radix2 #(.width(width)) rd_st8_1626  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1626]), .rdlo_in(a8_wr[1630]),  .coef_in(coef[512]), .rdup_out(a9_wr[1626]), .rdlo_out(a9_wr[1630]));
			radix2 #(.width(width)) rd_st8_1627  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1627]), .rdlo_in(a8_wr[1631]),  .coef_in(coef[768]), .rdup_out(a9_wr[1627]), .rdlo_out(a9_wr[1631]));
			radix2 #(.width(width)) rd_st8_1632  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1632]), .rdlo_in(a8_wr[1636]),  .coef_in(coef[0]), .rdup_out(a9_wr[1632]), .rdlo_out(a9_wr[1636]));
			radix2 #(.width(width)) rd_st8_1633  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1633]), .rdlo_in(a8_wr[1637]),  .coef_in(coef[256]), .rdup_out(a9_wr[1633]), .rdlo_out(a9_wr[1637]));
			radix2 #(.width(width)) rd_st8_1634  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1634]), .rdlo_in(a8_wr[1638]),  .coef_in(coef[512]), .rdup_out(a9_wr[1634]), .rdlo_out(a9_wr[1638]));
			radix2 #(.width(width)) rd_st8_1635  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1635]), .rdlo_in(a8_wr[1639]),  .coef_in(coef[768]), .rdup_out(a9_wr[1635]), .rdlo_out(a9_wr[1639]));
			radix2 #(.width(width)) rd_st8_1640  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1640]), .rdlo_in(a8_wr[1644]),  .coef_in(coef[0]), .rdup_out(a9_wr[1640]), .rdlo_out(a9_wr[1644]));
			radix2 #(.width(width)) rd_st8_1641  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1641]), .rdlo_in(a8_wr[1645]),  .coef_in(coef[256]), .rdup_out(a9_wr[1641]), .rdlo_out(a9_wr[1645]));
			radix2 #(.width(width)) rd_st8_1642  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1642]), .rdlo_in(a8_wr[1646]),  .coef_in(coef[512]), .rdup_out(a9_wr[1642]), .rdlo_out(a9_wr[1646]));
			radix2 #(.width(width)) rd_st8_1643  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1643]), .rdlo_in(a8_wr[1647]),  .coef_in(coef[768]), .rdup_out(a9_wr[1643]), .rdlo_out(a9_wr[1647]));
			radix2 #(.width(width)) rd_st8_1648  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1648]), .rdlo_in(a8_wr[1652]),  .coef_in(coef[0]), .rdup_out(a9_wr[1648]), .rdlo_out(a9_wr[1652]));
			radix2 #(.width(width)) rd_st8_1649  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1649]), .rdlo_in(a8_wr[1653]),  .coef_in(coef[256]), .rdup_out(a9_wr[1649]), .rdlo_out(a9_wr[1653]));
			radix2 #(.width(width)) rd_st8_1650  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1650]), .rdlo_in(a8_wr[1654]),  .coef_in(coef[512]), .rdup_out(a9_wr[1650]), .rdlo_out(a9_wr[1654]));
			radix2 #(.width(width)) rd_st8_1651  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1651]), .rdlo_in(a8_wr[1655]),  .coef_in(coef[768]), .rdup_out(a9_wr[1651]), .rdlo_out(a9_wr[1655]));
			radix2 #(.width(width)) rd_st8_1656  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1656]), .rdlo_in(a8_wr[1660]),  .coef_in(coef[0]), .rdup_out(a9_wr[1656]), .rdlo_out(a9_wr[1660]));
			radix2 #(.width(width)) rd_st8_1657  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1657]), .rdlo_in(a8_wr[1661]),  .coef_in(coef[256]), .rdup_out(a9_wr[1657]), .rdlo_out(a9_wr[1661]));
			radix2 #(.width(width)) rd_st8_1658  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1658]), .rdlo_in(a8_wr[1662]),  .coef_in(coef[512]), .rdup_out(a9_wr[1658]), .rdlo_out(a9_wr[1662]));
			radix2 #(.width(width)) rd_st8_1659  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1659]), .rdlo_in(a8_wr[1663]),  .coef_in(coef[768]), .rdup_out(a9_wr[1659]), .rdlo_out(a9_wr[1663]));
			radix2 #(.width(width)) rd_st8_1664  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1664]), .rdlo_in(a8_wr[1668]),  .coef_in(coef[0]), .rdup_out(a9_wr[1664]), .rdlo_out(a9_wr[1668]));
			radix2 #(.width(width)) rd_st8_1665  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1665]), .rdlo_in(a8_wr[1669]),  .coef_in(coef[256]), .rdup_out(a9_wr[1665]), .rdlo_out(a9_wr[1669]));
			radix2 #(.width(width)) rd_st8_1666  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1666]), .rdlo_in(a8_wr[1670]),  .coef_in(coef[512]), .rdup_out(a9_wr[1666]), .rdlo_out(a9_wr[1670]));
			radix2 #(.width(width)) rd_st8_1667  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1667]), .rdlo_in(a8_wr[1671]),  .coef_in(coef[768]), .rdup_out(a9_wr[1667]), .rdlo_out(a9_wr[1671]));
			radix2 #(.width(width)) rd_st8_1672  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1672]), .rdlo_in(a8_wr[1676]),  .coef_in(coef[0]), .rdup_out(a9_wr[1672]), .rdlo_out(a9_wr[1676]));
			radix2 #(.width(width)) rd_st8_1673  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1673]), .rdlo_in(a8_wr[1677]),  .coef_in(coef[256]), .rdup_out(a9_wr[1673]), .rdlo_out(a9_wr[1677]));
			radix2 #(.width(width)) rd_st8_1674  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1674]), .rdlo_in(a8_wr[1678]),  .coef_in(coef[512]), .rdup_out(a9_wr[1674]), .rdlo_out(a9_wr[1678]));
			radix2 #(.width(width)) rd_st8_1675  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1675]), .rdlo_in(a8_wr[1679]),  .coef_in(coef[768]), .rdup_out(a9_wr[1675]), .rdlo_out(a9_wr[1679]));
			radix2 #(.width(width)) rd_st8_1680  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1680]), .rdlo_in(a8_wr[1684]),  .coef_in(coef[0]), .rdup_out(a9_wr[1680]), .rdlo_out(a9_wr[1684]));
			radix2 #(.width(width)) rd_st8_1681  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1681]), .rdlo_in(a8_wr[1685]),  .coef_in(coef[256]), .rdup_out(a9_wr[1681]), .rdlo_out(a9_wr[1685]));
			radix2 #(.width(width)) rd_st8_1682  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1682]), .rdlo_in(a8_wr[1686]),  .coef_in(coef[512]), .rdup_out(a9_wr[1682]), .rdlo_out(a9_wr[1686]));
			radix2 #(.width(width)) rd_st8_1683  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1683]), .rdlo_in(a8_wr[1687]),  .coef_in(coef[768]), .rdup_out(a9_wr[1683]), .rdlo_out(a9_wr[1687]));
			radix2 #(.width(width)) rd_st8_1688  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1688]), .rdlo_in(a8_wr[1692]),  .coef_in(coef[0]), .rdup_out(a9_wr[1688]), .rdlo_out(a9_wr[1692]));
			radix2 #(.width(width)) rd_st8_1689  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1689]), .rdlo_in(a8_wr[1693]),  .coef_in(coef[256]), .rdup_out(a9_wr[1689]), .rdlo_out(a9_wr[1693]));
			radix2 #(.width(width)) rd_st8_1690  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1690]), .rdlo_in(a8_wr[1694]),  .coef_in(coef[512]), .rdup_out(a9_wr[1690]), .rdlo_out(a9_wr[1694]));
			radix2 #(.width(width)) rd_st8_1691  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1691]), .rdlo_in(a8_wr[1695]),  .coef_in(coef[768]), .rdup_out(a9_wr[1691]), .rdlo_out(a9_wr[1695]));
			radix2 #(.width(width)) rd_st8_1696  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1696]), .rdlo_in(a8_wr[1700]),  .coef_in(coef[0]), .rdup_out(a9_wr[1696]), .rdlo_out(a9_wr[1700]));
			radix2 #(.width(width)) rd_st8_1697  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1697]), .rdlo_in(a8_wr[1701]),  .coef_in(coef[256]), .rdup_out(a9_wr[1697]), .rdlo_out(a9_wr[1701]));
			radix2 #(.width(width)) rd_st8_1698  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1698]), .rdlo_in(a8_wr[1702]),  .coef_in(coef[512]), .rdup_out(a9_wr[1698]), .rdlo_out(a9_wr[1702]));
			radix2 #(.width(width)) rd_st8_1699  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1699]), .rdlo_in(a8_wr[1703]),  .coef_in(coef[768]), .rdup_out(a9_wr[1699]), .rdlo_out(a9_wr[1703]));
			radix2 #(.width(width)) rd_st8_1704  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1704]), .rdlo_in(a8_wr[1708]),  .coef_in(coef[0]), .rdup_out(a9_wr[1704]), .rdlo_out(a9_wr[1708]));
			radix2 #(.width(width)) rd_st8_1705  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1705]), .rdlo_in(a8_wr[1709]),  .coef_in(coef[256]), .rdup_out(a9_wr[1705]), .rdlo_out(a9_wr[1709]));
			radix2 #(.width(width)) rd_st8_1706  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1706]), .rdlo_in(a8_wr[1710]),  .coef_in(coef[512]), .rdup_out(a9_wr[1706]), .rdlo_out(a9_wr[1710]));
			radix2 #(.width(width)) rd_st8_1707  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1707]), .rdlo_in(a8_wr[1711]),  .coef_in(coef[768]), .rdup_out(a9_wr[1707]), .rdlo_out(a9_wr[1711]));
			radix2 #(.width(width)) rd_st8_1712  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1712]), .rdlo_in(a8_wr[1716]),  .coef_in(coef[0]), .rdup_out(a9_wr[1712]), .rdlo_out(a9_wr[1716]));
			radix2 #(.width(width)) rd_st8_1713  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1713]), .rdlo_in(a8_wr[1717]),  .coef_in(coef[256]), .rdup_out(a9_wr[1713]), .rdlo_out(a9_wr[1717]));
			radix2 #(.width(width)) rd_st8_1714  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1714]), .rdlo_in(a8_wr[1718]),  .coef_in(coef[512]), .rdup_out(a9_wr[1714]), .rdlo_out(a9_wr[1718]));
			radix2 #(.width(width)) rd_st8_1715  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1715]), .rdlo_in(a8_wr[1719]),  .coef_in(coef[768]), .rdup_out(a9_wr[1715]), .rdlo_out(a9_wr[1719]));
			radix2 #(.width(width)) rd_st8_1720  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1720]), .rdlo_in(a8_wr[1724]),  .coef_in(coef[0]), .rdup_out(a9_wr[1720]), .rdlo_out(a9_wr[1724]));
			radix2 #(.width(width)) rd_st8_1721  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1721]), .rdlo_in(a8_wr[1725]),  .coef_in(coef[256]), .rdup_out(a9_wr[1721]), .rdlo_out(a9_wr[1725]));
			radix2 #(.width(width)) rd_st8_1722  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1722]), .rdlo_in(a8_wr[1726]),  .coef_in(coef[512]), .rdup_out(a9_wr[1722]), .rdlo_out(a9_wr[1726]));
			radix2 #(.width(width)) rd_st8_1723  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1723]), .rdlo_in(a8_wr[1727]),  .coef_in(coef[768]), .rdup_out(a9_wr[1723]), .rdlo_out(a9_wr[1727]));
			radix2 #(.width(width)) rd_st8_1728  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1728]), .rdlo_in(a8_wr[1732]),  .coef_in(coef[0]), .rdup_out(a9_wr[1728]), .rdlo_out(a9_wr[1732]));
			radix2 #(.width(width)) rd_st8_1729  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1729]), .rdlo_in(a8_wr[1733]),  .coef_in(coef[256]), .rdup_out(a9_wr[1729]), .rdlo_out(a9_wr[1733]));
			radix2 #(.width(width)) rd_st8_1730  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1730]), .rdlo_in(a8_wr[1734]),  .coef_in(coef[512]), .rdup_out(a9_wr[1730]), .rdlo_out(a9_wr[1734]));
			radix2 #(.width(width)) rd_st8_1731  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1731]), .rdlo_in(a8_wr[1735]),  .coef_in(coef[768]), .rdup_out(a9_wr[1731]), .rdlo_out(a9_wr[1735]));
			radix2 #(.width(width)) rd_st8_1736  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1736]), .rdlo_in(a8_wr[1740]),  .coef_in(coef[0]), .rdup_out(a9_wr[1736]), .rdlo_out(a9_wr[1740]));
			radix2 #(.width(width)) rd_st8_1737  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1737]), .rdlo_in(a8_wr[1741]),  .coef_in(coef[256]), .rdup_out(a9_wr[1737]), .rdlo_out(a9_wr[1741]));
			radix2 #(.width(width)) rd_st8_1738  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1738]), .rdlo_in(a8_wr[1742]),  .coef_in(coef[512]), .rdup_out(a9_wr[1738]), .rdlo_out(a9_wr[1742]));
			radix2 #(.width(width)) rd_st8_1739  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1739]), .rdlo_in(a8_wr[1743]),  .coef_in(coef[768]), .rdup_out(a9_wr[1739]), .rdlo_out(a9_wr[1743]));
			radix2 #(.width(width)) rd_st8_1744  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1744]), .rdlo_in(a8_wr[1748]),  .coef_in(coef[0]), .rdup_out(a9_wr[1744]), .rdlo_out(a9_wr[1748]));
			radix2 #(.width(width)) rd_st8_1745  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1745]), .rdlo_in(a8_wr[1749]),  .coef_in(coef[256]), .rdup_out(a9_wr[1745]), .rdlo_out(a9_wr[1749]));
			radix2 #(.width(width)) rd_st8_1746  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1746]), .rdlo_in(a8_wr[1750]),  .coef_in(coef[512]), .rdup_out(a9_wr[1746]), .rdlo_out(a9_wr[1750]));
			radix2 #(.width(width)) rd_st8_1747  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1747]), .rdlo_in(a8_wr[1751]),  .coef_in(coef[768]), .rdup_out(a9_wr[1747]), .rdlo_out(a9_wr[1751]));
			radix2 #(.width(width)) rd_st8_1752  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1752]), .rdlo_in(a8_wr[1756]),  .coef_in(coef[0]), .rdup_out(a9_wr[1752]), .rdlo_out(a9_wr[1756]));
			radix2 #(.width(width)) rd_st8_1753  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1753]), .rdlo_in(a8_wr[1757]),  .coef_in(coef[256]), .rdup_out(a9_wr[1753]), .rdlo_out(a9_wr[1757]));
			radix2 #(.width(width)) rd_st8_1754  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1754]), .rdlo_in(a8_wr[1758]),  .coef_in(coef[512]), .rdup_out(a9_wr[1754]), .rdlo_out(a9_wr[1758]));
			radix2 #(.width(width)) rd_st8_1755  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1755]), .rdlo_in(a8_wr[1759]),  .coef_in(coef[768]), .rdup_out(a9_wr[1755]), .rdlo_out(a9_wr[1759]));
			radix2 #(.width(width)) rd_st8_1760  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1760]), .rdlo_in(a8_wr[1764]),  .coef_in(coef[0]), .rdup_out(a9_wr[1760]), .rdlo_out(a9_wr[1764]));
			radix2 #(.width(width)) rd_st8_1761  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1761]), .rdlo_in(a8_wr[1765]),  .coef_in(coef[256]), .rdup_out(a9_wr[1761]), .rdlo_out(a9_wr[1765]));
			radix2 #(.width(width)) rd_st8_1762  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1762]), .rdlo_in(a8_wr[1766]),  .coef_in(coef[512]), .rdup_out(a9_wr[1762]), .rdlo_out(a9_wr[1766]));
			radix2 #(.width(width)) rd_st8_1763  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1763]), .rdlo_in(a8_wr[1767]),  .coef_in(coef[768]), .rdup_out(a9_wr[1763]), .rdlo_out(a9_wr[1767]));
			radix2 #(.width(width)) rd_st8_1768  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1768]), .rdlo_in(a8_wr[1772]),  .coef_in(coef[0]), .rdup_out(a9_wr[1768]), .rdlo_out(a9_wr[1772]));
			radix2 #(.width(width)) rd_st8_1769  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1769]), .rdlo_in(a8_wr[1773]),  .coef_in(coef[256]), .rdup_out(a9_wr[1769]), .rdlo_out(a9_wr[1773]));
			radix2 #(.width(width)) rd_st8_1770  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1770]), .rdlo_in(a8_wr[1774]),  .coef_in(coef[512]), .rdup_out(a9_wr[1770]), .rdlo_out(a9_wr[1774]));
			radix2 #(.width(width)) rd_st8_1771  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1771]), .rdlo_in(a8_wr[1775]),  .coef_in(coef[768]), .rdup_out(a9_wr[1771]), .rdlo_out(a9_wr[1775]));
			radix2 #(.width(width)) rd_st8_1776  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1776]), .rdlo_in(a8_wr[1780]),  .coef_in(coef[0]), .rdup_out(a9_wr[1776]), .rdlo_out(a9_wr[1780]));
			radix2 #(.width(width)) rd_st8_1777  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1777]), .rdlo_in(a8_wr[1781]),  .coef_in(coef[256]), .rdup_out(a9_wr[1777]), .rdlo_out(a9_wr[1781]));
			radix2 #(.width(width)) rd_st8_1778  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1778]), .rdlo_in(a8_wr[1782]),  .coef_in(coef[512]), .rdup_out(a9_wr[1778]), .rdlo_out(a9_wr[1782]));
			radix2 #(.width(width)) rd_st8_1779  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1779]), .rdlo_in(a8_wr[1783]),  .coef_in(coef[768]), .rdup_out(a9_wr[1779]), .rdlo_out(a9_wr[1783]));
			radix2 #(.width(width)) rd_st8_1784  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1784]), .rdlo_in(a8_wr[1788]),  .coef_in(coef[0]), .rdup_out(a9_wr[1784]), .rdlo_out(a9_wr[1788]));
			radix2 #(.width(width)) rd_st8_1785  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1785]), .rdlo_in(a8_wr[1789]),  .coef_in(coef[256]), .rdup_out(a9_wr[1785]), .rdlo_out(a9_wr[1789]));
			radix2 #(.width(width)) rd_st8_1786  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1786]), .rdlo_in(a8_wr[1790]),  .coef_in(coef[512]), .rdup_out(a9_wr[1786]), .rdlo_out(a9_wr[1790]));
			radix2 #(.width(width)) rd_st8_1787  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1787]), .rdlo_in(a8_wr[1791]),  .coef_in(coef[768]), .rdup_out(a9_wr[1787]), .rdlo_out(a9_wr[1791]));
			radix2 #(.width(width)) rd_st8_1792  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1792]), .rdlo_in(a8_wr[1796]),  .coef_in(coef[0]), .rdup_out(a9_wr[1792]), .rdlo_out(a9_wr[1796]));
			radix2 #(.width(width)) rd_st8_1793  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1793]), .rdlo_in(a8_wr[1797]),  .coef_in(coef[256]), .rdup_out(a9_wr[1793]), .rdlo_out(a9_wr[1797]));
			radix2 #(.width(width)) rd_st8_1794  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1794]), .rdlo_in(a8_wr[1798]),  .coef_in(coef[512]), .rdup_out(a9_wr[1794]), .rdlo_out(a9_wr[1798]));
			radix2 #(.width(width)) rd_st8_1795  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1795]), .rdlo_in(a8_wr[1799]),  .coef_in(coef[768]), .rdup_out(a9_wr[1795]), .rdlo_out(a9_wr[1799]));
			radix2 #(.width(width)) rd_st8_1800  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1800]), .rdlo_in(a8_wr[1804]),  .coef_in(coef[0]), .rdup_out(a9_wr[1800]), .rdlo_out(a9_wr[1804]));
			radix2 #(.width(width)) rd_st8_1801  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1801]), .rdlo_in(a8_wr[1805]),  .coef_in(coef[256]), .rdup_out(a9_wr[1801]), .rdlo_out(a9_wr[1805]));
			radix2 #(.width(width)) rd_st8_1802  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1802]), .rdlo_in(a8_wr[1806]),  .coef_in(coef[512]), .rdup_out(a9_wr[1802]), .rdlo_out(a9_wr[1806]));
			radix2 #(.width(width)) rd_st8_1803  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1803]), .rdlo_in(a8_wr[1807]),  .coef_in(coef[768]), .rdup_out(a9_wr[1803]), .rdlo_out(a9_wr[1807]));
			radix2 #(.width(width)) rd_st8_1808  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1808]), .rdlo_in(a8_wr[1812]),  .coef_in(coef[0]), .rdup_out(a9_wr[1808]), .rdlo_out(a9_wr[1812]));
			radix2 #(.width(width)) rd_st8_1809  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1809]), .rdlo_in(a8_wr[1813]),  .coef_in(coef[256]), .rdup_out(a9_wr[1809]), .rdlo_out(a9_wr[1813]));
			radix2 #(.width(width)) rd_st8_1810  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1810]), .rdlo_in(a8_wr[1814]),  .coef_in(coef[512]), .rdup_out(a9_wr[1810]), .rdlo_out(a9_wr[1814]));
			radix2 #(.width(width)) rd_st8_1811  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1811]), .rdlo_in(a8_wr[1815]),  .coef_in(coef[768]), .rdup_out(a9_wr[1811]), .rdlo_out(a9_wr[1815]));
			radix2 #(.width(width)) rd_st8_1816  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1816]), .rdlo_in(a8_wr[1820]),  .coef_in(coef[0]), .rdup_out(a9_wr[1816]), .rdlo_out(a9_wr[1820]));
			radix2 #(.width(width)) rd_st8_1817  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1817]), .rdlo_in(a8_wr[1821]),  .coef_in(coef[256]), .rdup_out(a9_wr[1817]), .rdlo_out(a9_wr[1821]));
			radix2 #(.width(width)) rd_st8_1818  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1818]), .rdlo_in(a8_wr[1822]),  .coef_in(coef[512]), .rdup_out(a9_wr[1818]), .rdlo_out(a9_wr[1822]));
			radix2 #(.width(width)) rd_st8_1819  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1819]), .rdlo_in(a8_wr[1823]),  .coef_in(coef[768]), .rdup_out(a9_wr[1819]), .rdlo_out(a9_wr[1823]));
			radix2 #(.width(width)) rd_st8_1824  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1824]), .rdlo_in(a8_wr[1828]),  .coef_in(coef[0]), .rdup_out(a9_wr[1824]), .rdlo_out(a9_wr[1828]));
			radix2 #(.width(width)) rd_st8_1825  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1825]), .rdlo_in(a8_wr[1829]),  .coef_in(coef[256]), .rdup_out(a9_wr[1825]), .rdlo_out(a9_wr[1829]));
			radix2 #(.width(width)) rd_st8_1826  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1826]), .rdlo_in(a8_wr[1830]),  .coef_in(coef[512]), .rdup_out(a9_wr[1826]), .rdlo_out(a9_wr[1830]));
			radix2 #(.width(width)) rd_st8_1827  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1827]), .rdlo_in(a8_wr[1831]),  .coef_in(coef[768]), .rdup_out(a9_wr[1827]), .rdlo_out(a9_wr[1831]));
			radix2 #(.width(width)) rd_st8_1832  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1832]), .rdlo_in(a8_wr[1836]),  .coef_in(coef[0]), .rdup_out(a9_wr[1832]), .rdlo_out(a9_wr[1836]));
			radix2 #(.width(width)) rd_st8_1833  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1833]), .rdlo_in(a8_wr[1837]),  .coef_in(coef[256]), .rdup_out(a9_wr[1833]), .rdlo_out(a9_wr[1837]));
			radix2 #(.width(width)) rd_st8_1834  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1834]), .rdlo_in(a8_wr[1838]),  .coef_in(coef[512]), .rdup_out(a9_wr[1834]), .rdlo_out(a9_wr[1838]));
			radix2 #(.width(width)) rd_st8_1835  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1835]), .rdlo_in(a8_wr[1839]),  .coef_in(coef[768]), .rdup_out(a9_wr[1835]), .rdlo_out(a9_wr[1839]));
			radix2 #(.width(width)) rd_st8_1840  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1840]), .rdlo_in(a8_wr[1844]),  .coef_in(coef[0]), .rdup_out(a9_wr[1840]), .rdlo_out(a9_wr[1844]));
			radix2 #(.width(width)) rd_st8_1841  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1841]), .rdlo_in(a8_wr[1845]),  .coef_in(coef[256]), .rdup_out(a9_wr[1841]), .rdlo_out(a9_wr[1845]));
			radix2 #(.width(width)) rd_st8_1842  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1842]), .rdlo_in(a8_wr[1846]),  .coef_in(coef[512]), .rdup_out(a9_wr[1842]), .rdlo_out(a9_wr[1846]));
			radix2 #(.width(width)) rd_st8_1843  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1843]), .rdlo_in(a8_wr[1847]),  .coef_in(coef[768]), .rdup_out(a9_wr[1843]), .rdlo_out(a9_wr[1847]));
			radix2 #(.width(width)) rd_st8_1848  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1848]), .rdlo_in(a8_wr[1852]),  .coef_in(coef[0]), .rdup_out(a9_wr[1848]), .rdlo_out(a9_wr[1852]));
			radix2 #(.width(width)) rd_st8_1849  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1849]), .rdlo_in(a8_wr[1853]),  .coef_in(coef[256]), .rdup_out(a9_wr[1849]), .rdlo_out(a9_wr[1853]));
			radix2 #(.width(width)) rd_st8_1850  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1850]), .rdlo_in(a8_wr[1854]),  .coef_in(coef[512]), .rdup_out(a9_wr[1850]), .rdlo_out(a9_wr[1854]));
			radix2 #(.width(width)) rd_st8_1851  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1851]), .rdlo_in(a8_wr[1855]),  .coef_in(coef[768]), .rdup_out(a9_wr[1851]), .rdlo_out(a9_wr[1855]));
			radix2 #(.width(width)) rd_st8_1856  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1856]), .rdlo_in(a8_wr[1860]),  .coef_in(coef[0]), .rdup_out(a9_wr[1856]), .rdlo_out(a9_wr[1860]));
			radix2 #(.width(width)) rd_st8_1857  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1857]), .rdlo_in(a8_wr[1861]),  .coef_in(coef[256]), .rdup_out(a9_wr[1857]), .rdlo_out(a9_wr[1861]));
			radix2 #(.width(width)) rd_st8_1858  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1858]), .rdlo_in(a8_wr[1862]),  .coef_in(coef[512]), .rdup_out(a9_wr[1858]), .rdlo_out(a9_wr[1862]));
			radix2 #(.width(width)) rd_st8_1859  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1859]), .rdlo_in(a8_wr[1863]),  .coef_in(coef[768]), .rdup_out(a9_wr[1859]), .rdlo_out(a9_wr[1863]));
			radix2 #(.width(width)) rd_st8_1864  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1864]), .rdlo_in(a8_wr[1868]),  .coef_in(coef[0]), .rdup_out(a9_wr[1864]), .rdlo_out(a9_wr[1868]));
			radix2 #(.width(width)) rd_st8_1865  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1865]), .rdlo_in(a8_wr[1869]),  .coef_in(coef[256]), .rdup_out(a9_wr[1865]), .rdlo_out(a9_wr[1869]));
			radix2 #(.width(width)) rd_st8_1866  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1866]), .rdlo_in(a8_wr[1870]),  .coef_in(coef[512]), .rdup_out(a9_wr[1866]), .rdlo_out(a9_wr[1870]));
			radix2 #(.width(width)) rd_st8_1867  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1867]), .rdlo_in(a8_wr[1871]),  .coef_in(coef[768]), .rdup_out(a9_wr[1867]), .rdlo_out(a9_wr[1871]));
			radix2 #(.width(width)) rd_st8_1872  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1872]), .rdlo_in(a8_wr[1876]),  .coef_in(coef[0]), .rdup_out(a9_wr[1872]), .rdlo_out(a9_wr[1876]));
			radix2 #(.width(width)) rd_st8_1873  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1873]), .rdlo_in(a8_wr[1877]),  .coef_in(coef[256]), .rdup_out(a9_wr[1873]), .rdlo_out(a9_wr[1877]));
			radix2 #(.width(width)) rd_st8_1874  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1874]), .rdlo_in(a8_wr[1878]),  .coef_in(coef[512]), .rdup_out(a9_wr[1874]), .rdlo_out(a9_wr[1878]));
			radix2 #(.width(width)) rd_st8_1875  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1875]), .rdlo_in(a8_wr[1879]),  .coef_in(coef[768]), .rdup_out(a9_wr[1875]), .rdlo_out(a9_wr[1879]));
			radix2 #(.width(width)) rd_st8_1880  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1880]), .rdlo_in(a8_wr[1884]),  .coef_in(coef[0]), .rdup_out(a9_wr[1880]), .rdlo_out(a9_wr[1884]));
			radix2 #(.width(width)) rd_st8_1881  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1881]), .rdlo_in(a8_wr[1885]),  .coef_in(coef[256]), .rdup_out(a9_wr[1881]), .rdlo_out(a9_wr[1885]));
			radix2 #(.width(width)) rd_st8_1882  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1882]), .rdlo_in(a8_wr[1886]),  .coef_in(coef[512]), .rdup_out(a9_wr[1882]), .rdlo_out(a9_wr[1886]));
			radix2 #(.width(width)) rd_st8_1883  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1883]), .rdlo_in(a8_wr[1887]),  .coef_in(coef[768]), .rdup_out(a9_wr[1883]), .rdlo_out(a9_wr[1887]));
			radix2 #(.width(width)) rd_st8_1888  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1888]), .rdlo_in(a8_wr[1892]),  .coef_in(coef[0]), .rdup_out(a9_wr[1888]), .rdlo_out(a9_wr[1892]));
			radix2 #(.width(width)) rd_st8_1889  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1889]), .rdlo_in(a8_wr[1893]),  .coef_in(coef[256]), .rdup_out(a9_wr[1889]), .rdlo_out(a9_wr[1893]));
			radix2 #(.width(width)) rd_st8_1890  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1890]), .rdlo_in(a8_wr[1894]),  .coef_in(coef[512]), .rdup_out(a9_wr[1890]), .rdlo_out(a9_wr[1894]));
			radix2 #(.width(width)) rd_st8_1891  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1891]), .rdlo_in(a8_wr[1895]),  .coef_in(coef[768]), .rdup_out(a9_wr[1891]), .rdlo_out(a9_wr[1895]));
			radix2 #(.width(width)) rd_st8_1896  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1896]), .rdlo_in(a8_wr[1900]),  .coef_in(coef[0]), .rdup_out(a9_wr[1896]), .rdlo_out(a9_wr[1900]));
			radix2 #(.width(width)) rd_st8_1897  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1897]), .rdlo_in(a8_wr[1901]),  .coef_in(coef[256]), .rdup_out(a9_wr[1897]), .rdlo_out(a9_wr[1901]));
			radix2 #(.width(width)) rd_st8_1898  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1898]), .rdlo_in(a8_wr[1902]),  .coef_in(coef[512]), .rdup_out(a9_wr[1898]), .rdlo_out(a9_wr[1902]));
			radix2 #(.width(width)) rd_st8_1899  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1899]), .rdlo_in(a8_wr[1903]),  .coef_in(coef[768]), .rdup_out(a9_wr[1899]), .rdlo_out(a9_wr[1903]));
			radix2 #(.width(width)) rd_st8_1904  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1904]), .rdlo_in(a8_wr[1908]),  .coef_in(coef[0]), .rdup_out(a9_wr[1904]), .rdlo_out(a9_wr[1908]));
			radix2 #(.width(width)) rd_st8_1905  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1905]), .rdlo_in(a8_wr[1909]),  .coef_in(coef[256]), .rdup_out(a9_wr[1905]), .rdlo_out(a9_wr[1909]));
			radix2 #(.width(width)) rd_st8_1906  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1906]), .rdlo_in(a8_wr[1910]),  .coef_in(coef[512]), .rdup_out(a9_wr[1906]), .rdlo_out(a9_wr[1910]));
			radix2 #(.width(width)) rd_st8_1907  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1907]), .rdlo_in(a8_wr[1911]),  .coef_in(coef[768]), .rdup_out(a9_wr[1907]), .rdlo_out(a9_wr[1911]));
			radix2 #(.width(width)) rd_st8_1912  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1912]), .rdlo_in(a8_wr[1916]),  .coef_in(coef[0]), .rdup_out(a9_wr[1912]), .rdlo_out(a9_wr[1916]));
			radix2 #(.width(width)) rd_st8_1913  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1913]), .rdlo_in(a8_wr[1917]),  .coef_in(coef[256]), .rdup_out(a9_wr[1913]), .rdlo_out(a9_wr[1917]));
			radix2 #(.width(width)) rd_st8_1914  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1914]), .rdlo_in(a8_wr[1918]),  .coef_in(coef[512]), .rdup_out(a9_wr[1914]), .rdlo_out(a9_wr[1918]));
			radix2 #(.width(width)) rd_st8_1915  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1915]), .rdlo_in(a8_wr[1919]),  .coef_in(coef[768]), .rdup_out(a9_wr[1915]), .rdlo_out(a9_wr[1919]));
			radix2 #(.width(width)) rd_st8_1920  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1920]), .rdlo_in(a8_wr[1924]),  .coef_in(coef[0]), .rdup_out(a9_wr[1920]), .rdlo_out(a9_wr[1924]));
			radix2 #(.width(width)) rd_st8_1921  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1921]), .rdlo_in(a8_wr[1925]),  .coef_in(coef[256]), .rdup_out(a9_wr[1921]), .rdlo_out(a9_wr[1925]));
			radix2 #(.width(width)) rd_st8_1922  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1922]), .rdlo_in(a8_wr[1926]),  .coef_in(coef[512]), .rdup_out(a9_wr[1922]), .rdlo_out(a9_wr[1926]));
			radix2 #(.width(width)) rd_st8_1923  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1923]), .rdlo_in(a8_wr[1927]),  .coef_in(coef[768]), .rdup_out(a9_wr[1923]), .rdlo_out(a9_wr[1927]));
			radix2 #(.width(width)) rd_st8_1928  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1928]), .rdlo_in(a8_wr[1932]),  .coef_in(coef[0]), .rdup_out(a9_wr[1928]), .rdlo_out(a9_wr[1932]));
			radix2 #(.width(width)) rd_st8_1929  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1929]), .rdlo_in(a8_wr[1933]),  .coef_in(coef[256]), .rdup_out(a9_wr[1929]), .rdlo_out(a9_wr[1933]));
			radix2 #(.width(width)) rd_st8_1930  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1930]), .rdlo_in(a8_wr[1934]),  .coef_in(coef[512]), .rdup_out(a9_wr[1930]), .rdlo_out(a9_wr[1934]));
			radix2 #(.width(width)) rd_st8_1931  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1931]), .rdlo_in(a8_wr[1935]),  .coef_in(coef[768]), .rdup_out(a9_wr[1931]), .rdlo_out(a9_wr[1935]));
			radix2 #(.width(width)) rd_st8_1936  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1936]), .rdlo_in(a8_wr[1940]),  .coef_in(coef[0]), .rdup_out(a9_wr[1936]), .rdlo_out(a9_wr[1940]));
			radix2 #(.width(width)) rd_st8_1937  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1937]), .rdlo_in(a8_wr[1941]),  .coef_in(coef[256]), .rdup_out(a9_wr[1937]), .rdlo_out(a9_wr[1941]));
			radix2 #(.width(width)) rd_st8_1938  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1938]), .rdlo_in(a8_wr[1942]),  .coef_in(coef[512]), .rdup_out(a9_wr[1938]), .rdlo_out(a9_wr[1942]));
			radix2 #(.width(width)) rd_st8_1939  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1939]), .rdlo_in(a8_wr[1943]),  .coef_in(coef[768]), .rdup_out(a9_wr[1939]), .rdlo_out(a9_wr[1943]));
			radix2 #(.width(width)) rd_st8_1944  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1944]), .rdlo_in(a8_wr[1948]),  .coef_in(coef[0]), .rdup_out(a9_wr[1944]), .rdlo_out(a9_wr[1948]));
			radix2 #(.width(width)) rd_st8_1945  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1945]), .rdlo_in(a8_wr[1949]),  .coef_in(coef[256]), .rdup_out(a9_wr[1945]), .rdlo_out(a9_wr[1949]));
			radix2 #(.width(width)) rd_st8_1946  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1946]), .rdlo_in(a8_wr[1950]),  .coef_in(coef[512]), .rdup_out(a9_wr[1946]), .rdlo_out(a9_wr[1950]));
			radix2 #(.width(width)) rd_st8_1947  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1947]), .rdlo_in(a8_wr[1951]),  .coef_in(coef[768]), .rdup_out(a9_wr[1947]), .rdlo_out(a9_wr[1951]));
			radix2 #(.width(width)) rd_st8_1952  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1952]), .rdlo_in(a8_wr[1956]),  .coef_in(coef[0]), .rdup_out(a9_wr[1952]), .rdlo_out(a9_wr[1956]));
			radix2 #(.width(width)) rd_st8_1953  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1953]), .rdlo_in(a8_wr[1957]),  .coef_in(coef[256]), .rdup_out(a9_wr[1953]), .rdlo_out(a9_wr[1957]));
			radix2 #(.width(width)) rd_st8_1954  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1954]), .rdlo_in(a8_wr[1958]),  .coef_in(coef[512]), .rdup_out(a9_wr[1954]), .rdlo_out(a9_wr[1958]));
			radix2 #(.width(width)) rd_st8_1955  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1955]), .rdlo_in(a8_wr[1959]),  .coef_in(coef[768]), .rdup_out(a9_wr[1955]), .rdlo_out(a9_wr[1959]));
			radix2 #(.width(width)) rd_st8_1960  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1960]), .rdlo_in(a8_wr[1964]),  .coef_in(coef[0]), .rdup_out(a9_wr[1960]), .rdlo_out(a9_wr[1964]));
			radix2 #(.width(width)) rd_st8_1961  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1961]), .rdlo_in(a8_wr[1965]),  .coef_in(coef[256]), .rdup_out(a9_wr[1961]), .rdlo_out(a9_wr[1965]));
			radix2 #(.width(width)) rd_st8_1962  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1962]), .rdlo_in(a8_wr[1966]),  .coef_in(coef[512]), .rdup_out(a9_wr[1962]), .rdlo_out(a9_wr[1966]));
			radix2 #(.width(width)) rd_st8_1963  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1963]), .rdlo_in(a8_wr[1967]),  .coef_in(coef[768]), .rdup_out(a9_wr[1963]), .rdlo_out(a9_wr[1967]));
			radix2 #(.width(width)) rd_st8_1968  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1968]), .rdlo_in(a8_wr[1972]),  .coef_in(coef[0]), .rdup_out(a9_wr[1968]), .rdlo_out(a9_wr[1972]));
			radix2 #(.width(width)) rd_st8_1969  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1969]), .rdlo_in(a8_wr[1973]),  .coef_in(coef[256]), .rdup_out(a9_wr[1969]), .rdlo_out(a9_wr[1973]));
			radix2 #(.width(width)) rd_st8_1970  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1970]), .rdlo_in(a8_wr[1974]),  .coef_in(coef[512]), .rdup_out(a9_wr[1970]), .rdlo_out(a9_wr[1974]));
			radix2 #(.width(width)) rd_st8_1971  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1971]), .rdlo_in(a8_wr[1975]),  .coef_in(coef[768]), .rdup_out(a9_wr[1971]), .rdlo_out(a9_wr[1975]));
			radix2 #(.width(width)) rd_st8_1976  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1976]), .rdlo_in(a8_wr[1980]),  .coef_in(coef[0]), .rdup_out(a9_wr[1976]), .rdlo_out(a9_wr[1980]));
			radix2 #(.width(width)) rd_st8_1977  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1977]), .rdlo_in(a8_wr[1981]),  .coef_in(coef[256]), .rdup_out(a9_wr[1977]), .rdlo_out(a9_wr[1981]));
			radix2 #(.width(width)) rd_st8_1978  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1978]), .rdlo_in(a8_wr[1982]),  .coef_in(coef[512]), .rdup_out(a9_wr[1978]), .rdlo_out(a9_wr[1982]));
			radix2 #(.width(width)) rd_st8_1979  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1979]), .rdlo_in(a8_wr[1983]),  .coef_in(coef[768]), .rdup_out(a9_wr[1979]), .rdlo_out(a9_wr[1983]));
			radix2 #(.width(width)) rd_st8_1984  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1984]), .rdlo_in(a8_wr[1988]),  .coef_in(coef[0]), .rdup_out(a9_wr[1984]), .rdlo_out(a9_wr[1988]));
			radix2 #(.width(width)) rd_st8_1985  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1985]), .rdlo_in(a8_wr[1989]),  .coef_in(coef[256]), .rdup_out(a9_wr[1985]), .rdlo_out(a9_wr[1989]));
			radix2 #(.width(width)) rd_st8_1986  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1986]), .rdlo_in(a8_wr[1990]),  .coef_in(coef[512]), .rdup_out(a9_wr[1986]), .rdlo_out(a9_wr[1990]));
			radix2 #(.width(width)) rd_st8_1987  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1987]), .rdlo_in(a8_wr[1991]),  .coef_in(coef[768]), .rdup_out(a9_wr[1987]), .rdlo_out(a9_wr[1991]));
			radix2 #(.width(width)) rd_st8_1992  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1992]), .rdlo_in(a8_wr[1996]),  .coef_in(coef[0]), .rdup_out(a9_wr[1992]), .rdlo_out(a9_wr[1996]));
			radix2 #(.width(width)) rd_st8_1993  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1993]), .rdlo_in(a8_wr[1997]),  .coef_in(coef[256]), .rdup_out(a9_wr[1993]), .rdlo_out(a9_wr[1997]));
			radix2 #(.width(width)) rd_st8_1994  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1994]), .rdlo_in(a8_wr[1998]),  .coef_in(coef[512]), .rdup_out(a9_wr[1994]), .rdlo_out(a9_wr[1998]));
			radix2 #(.width(width)) rd_st8_1995  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[1995]), .rdlo_in(a8_wr[1999]),  .coef_in(coef[768]), .rdup_out(a9_wr[1995]), .rdlo_out(a9_wr[1999]));
			radix2 #(.width(width)) rd_st8_2000  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[2000]), .rdlo_in(a8_wr[2004]),  .coef_in(coef[0]), .rdup_out(a9_wr[2000]), .rdlo_out(a9_wr[2004]));
			radix2 #(.width(width)) rd_st8_2001  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[2001]), .rdlo_in(a8_wr[2005]),  .coef_in(coef[256]), .rdup_out(a9_wr[2001]), .rdlo_out(a9_wr[2005]));
			radix2 #(.width(width)) rd_st8_2002  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[2002]), .rdlo_in(a8_wr[2006]),  .coef_in(coef[512]), .rdup_out(a9_wr[2002]), .rdlo_out(a9_wr[2006]));
			radix2 #(.width(width)) rd_st8_2003  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[2003]), .rdlo_in(a8_wr[2007]),  .coef_in(coef[768]), .rdup_out(a9_wr[2003]), .rdlo_out(a9_wr[2007]));
			radix2 #(.width(width)) rd_st8_2008  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[2008]), .rdlo_in(a8_wr[2012]),  .coef_in(coef[0]), .rdup_out(a9_wr[2008]), .rdlo_out(a9_wr[2012]));
			radix2 #(.width(width)) rd_st8_2009  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[2009]), .rdlo_in(a8_wr[2013]),  .coef_in(coef[256]), .rdup_out(a9_wr[2009]), .rdlo_out(a9_wr[2013]));
			radix2 #(.width(width)) rd_st8_2010  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[2010]), .rdlo_in(a8_wr[2014]),  .coef_in(coef[512]), .rdup_out(a9_wr[2010]), .rdlo_out(a9_wr[2014]));
			radix2 #(.width(width)) rd_st8_2011  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[2011]), .rdlo_in(a8_wr[2015]),  .coef_in(coef[768]), .rdup_out(a9_wr[2011]), .rdlo_out(a9_wr[2015]));
			radix2 #(.width(width)) rd_st8_2016  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[2016]), .rdlo_in(a8_wr[2020]),  .coef_in(coef[0]), .rdup_out(a9_wr[2016]), .rdlo_out(a9_wr[2020]));
			radix2 #(.width(width)) rd_st8_2017  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[2017]), .rdlo_in(a8_wr[2021]),  .coef_in(coef[256]), .rdup_out(a9_wr[2017]), .rdlo_out(a9_wr[2021]));
			radix2 #(.width(width)) rd_st8_2018  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[2018]), .rdlo_in(a8_wr[2022]),  .coef_in(coef[512]), .rdup_out(a9_wr[2018]), .rdlo_out(a9_wr[2022]));
			radix2 #(.width(width)) rd_st8_2019  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[2019]), .rdlo_in(a8_wr[2023]),  .coef_in(coef[768]), .rdup_out(a9_wr[2019]), .rdlo_out(a9_wr[2023]));
			radix2 #(.width(width)) rd_st8_2024  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[2024]), .rdlo_in(a8_wr[2028]),  .coef_in(coef[0]), .rdup_out(a9_wr[2024]), .rdlo_out(a9_wr[2028]));
			radix2 #(.width(width)) rd_st8_2025  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[2025]), .rdlo_in(a8_wr[2029]),  .coef_in(coef[256]), .rdup_out(a9_wr[2025]), .rdlo_out(a9_wr[2029]));
			radix2 #(.width(width)) rd_st8_2026  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[2026]), .rdlo_in(a8_wr[2030]),  .coef_in(coef[512]), .rdup_out(a9_wr[2026]), .rdlo_out(a9_wr[2030]));
			radix2 #(.width(width)) rd_st8_2027  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[2027]), .rdlo_in(a8_wr[2031]),  .coef_in(coef[768]), .rdup_out(a9_wr[2027]), .rdlo_out(a9_wr[2031]));
			radix2 #(.width(width)) rd_st8_2032  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[2032]), .rdlo_in(a8_wr[2036]),  .coef_in(coef[0]), .rdup_out(a9_wr[2032]), .rdlo_out(a9_wr[2036]));
			radix2 #(.width(width)) rd_st8_2033  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[2033]), .rdlo_in(a8_wr[2037]),  .coef_in(coef[256]), .rdup_out(a9_wr[2033]), .rdlo_out(a9_wr[2037]));
			radix2 #(.width(width)) rd_st8_2034  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[2034]), .rdlo_in(a8_wr[2038]),  .coef_in(coef[512]), .rdup_out(a9_wr[2034]), .rdlo_out(a9_wr[2038]));
			radix2 #(.width(width)) rd_st8_2035  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[2035]), .rdlo_in(a8_wr[2039]),  .coef_in(coef[768]), .rdup_out(a9_wr[2035]), .rdlo_out(a9_wr[2039]));
			radix2 #(.width(width)) rd_st8_2040  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[2040]), .rdlo_in(a8_wr[2044]),  .coef_in(coef[0]), .rdup_out(a9_wr[2040]), .rdlo_out(a9_wr[2044]));
			radix2 #(.width(width)) rd_st8_2041  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[2041]), .rdlo_in(a8_wr[2045]),  .coef_in(coef[256]), .rdup_out(a9_wr[2041]), .rdlo_out(a9_wr[2045]));
			radix2 #(.width(width)) rd_st8_2042  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[2042]), .rdlo_in(a8_wr[2046]),  .coef_in(coef[512]), .rdup_out(a9_wr[2042]), .rdlo_out(a9_wr[2046]));
			radix2 #(.width(width)) rd_st8_2043  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a8_wr[2043]), .rdlo_in(a8_wr[2047]),  .coef_in(coef[768]), .rdup_out(a9_wr[2043]), .rdlo_out(a9_wr[2047]));

		//--- radix stage 9
			radix2 #(.width(width)) rd_st9_0   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[0]), .rdlo_in(a9_wr[2]),  .coef_in(coef[0]), .rdup_out(a10_wr[0]), .rdlo_out(a10_wr[2]));
			radix2 #(.width(width)) rd_st9_1   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1]), .rdlo_in(a9_wr[3]),  .coef_in(coef[512]), .rdup_out(a10_wr[1]), .rdlo_out(a10_wr[3]));
			radix2 #(.width(width)) rd_st9_4   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[4]), .rdlo_in(a9_wr[6]),  .coef_in(coef[0]), .rdup_out(a10_wr[4]), .rdlo_out(a10_wr[6]));
			radix2 #(.width(width)) rd_st9_5   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[5]), .rdlo_in(a9_wr[7]),  .coef_in(coef[512]), .rdup_out(a10_wr[5]), .rdlo_out(a10_wr[7]));
			radix2 #(.width(width)) rd_st9_8   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[8]), .rdlo_in(a9_wr[10]),  .coef_in(coef[0]), .rdup_out(a10_wr[8]), .rdlo_out(a10_wr[10]));
			radix2 #(.width(width)) rd_st9_9   (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[9]), .rdlo_in(a9_wr[11]),  .coef_in(coef[512]), .rdup_out(a10_wr[9]), .rdlo_out(a10_wr[11]));
			radix2 #(.width(width)) rd_st9_12  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[12]), .rdlo_in(a9_wr[14]),  .coef_in(coef[0]), .rdup_out(a10_wr[12]), .rdlo_out(a10_wr[14]));
			radix2 #(.width(width)) rd_st9_13  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[13]), .rdlo_in(a9_wr[15]),  .coef_in(coef[512]), .rdup_out(a10_wr[13]), .rdlo_out(a10_wr[15]));
			radix2 #(.width(width)) rd_st9_16  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[16]), .rdlo_in(a9_wr[18]),  .coef_in(coef[0]), .rdup_out(a10_wr[16]), .rdlo_out(a10_wr[18]));
			radix2 #(.width(width)) rd_st9_17  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[17]), .rdlo_in(a9_wr[19]),  .coef_in(coef[512]), .rdup_out(a10_wr[17]), .rdlo_out(a10_wr[19]));
			radix2 #(.width(width)) rd_st9_20  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[20]), .rdlo_in(a9_wr[22]),  .coef_in(coef[0]), .rdup_out(a10_wr[20]), .rdlo_out(a10_wr[22]));
			radix2 #(.width(width)) rd_st9_21  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[21]), .rdlo_in(a9_wr[23]),  .coef_in(coef[512]), .rdup_out(a10_wr[21]), .rdlo_out(a10_wr[23]));
			radix2 #(.width(width)) rd_st9_24  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[24]), .rdlo_in(a9_wr[26]),  .coef_in(coef[0]), .rdup_out(a10_wr[24]), .rdlo_out(a10_wr[26]));
			radix2 #(.width(width)) rd_st9_25  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[25]), .rdlo_in(a9_wr[27]),  .coef_in(coef[512]), .rdup_out(a10_wr[25]), .rdlo_out(a10_wr[27]));
			radix2 #(.width(width)) rd_st9_28  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[28]), .rdlo_in(a9_wr[30]),  .coef_in(coef[0]), .rdup_out(a10_wr[28]), .rdlo_out(a10_wr[30]));
			radix2 #(.width(width)) rd_st9_29  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[29]), .rdlo_in(a9_wr[31]),  .coef_in(coef[512]), .rdup_out(a10_wr[29]), .rdlo_out(a10_wr[31]));
			radix2 #(.width(width)) rd_st9_32  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[32]), .rdlo_in(a9_wr[34]),  .coef_in(coef[0]), .rdup_out(a10_wr[32]), .rdlo_out(a10_wr[34]));
			radix2 #(.width(width)) rd_st9_33  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[33]), .rdlo_in(a9_wr[35]),  .coef_in(coef[512]), .rdup_out(a10_wr[33]), .rdlo_out(a10_wr[35]));
			radix2 #(.width(width)) rd_st9_36  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[36]), .rdlo_in(a9_wr[38]),  .coef_in(coef[0]), .rdup_out(a10_wr[36]), .rdlo_out(a10_wr[38]));
			radix2 #(.width(width)) rd_st9_37  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[37]), .rdlo_in(a9_wr[39]),  .coef_in(coef[512]), .rdup_out(a10_wr[37]), .rdlo_out(a10_wr[39]));
			radix2 #(.width(width)) rd_st9_40  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[40]), .rdlo_in(a9_wr[42]),  .coef_in(coef[0]), .rdup_out(a10_wr[40]), .rdlo_out(a10_wr[42]));
			radix2 #(.width(width)) rd_st9_41  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[41]), .rdlo_in(a9_wr[43]),  .coef_in(coef[512]), .rdup_out(a10_wr[41]), .rdlo_out(a10_wr[43]));
			radix2 #(.width(width)) rd_st9_44  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[44]), .rdlo_in(a9_wr[46]),  .coef_in(coef[0]), .rdup_out(a10_wr[44]), .rdlo_out(a10_wr[46]));
			radix2 #(.width(width)) rd_st9_45  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[45]), .rdlo_in(a9_wr[47]),  .coef_in(coef[512]), .rdup_out(a10_wr[45]), .rdlo_out(a10_wr[47]));
			radix2 #(.width(width)) rd_st9_48  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[48]), .rdlo_in(a9_wr[50]),  .coef_in(coef[0]), .rdup_out(a10_wr[48]), .rdlo_out(a10_wr[50]));
			radix2 #(.width(width)) rd_st9_49  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[49]), .rdlo_in(a9_wr[51]),  .coef_in(coef[512]), .rdup_out(a10_wr[49]), .rdlo_out(a10_wr[51]));
			radix2 #(.width(width)) rd_st9_52  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[52]), .rdlo_in(a9_wr[54]),  .coef_in(coef[0]), .rdup_out(a10_wr[52]), .rdlo_out(a10_wr[54]));
			radix2 #(.width(width)) rd_st9_53  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[53]), .rdlo_in(a9_wr[55]),  .coef_in(coef[512]), .rdup_out(a10_wr[53]), .rdlo_out(a10_wr[55]));
			radix2 #(.width(width)) rd_st9_56  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[56]), .rdlo_in(a9_wr[58]),  .coef_in(coef[0]), .rdup_out(a10_wr[56]), .rdlo_out(a10_wr[58]));
			radix2 #(.width(width)) rd_st9_57  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[57]), .rdlo_in(a9_wr[59]),  .coef_in(coef[512]), .rdup_out(a10_wr[57]), .rdlo_out(a10_wr[59]));
			radix2 #(.width(width)) rd_st9_60  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[60]), .rdlo_in(a9_wr[62]),  .coef_in(coef[0]), .rdup_out(a10_wr[60]), .rdlo_out(a10_wr[62]));
			radix2 #(.width(width)) rd_st9_61  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[61]), .rdlo_in(a9_wr[63]),  .coef_in(coef[512]), .rdup_out(a10_wr[61]), .rdlo_out(a10_wr[63]));
			radix2 #(.width(width)) rd_st9_64  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[64]), .rdlo_in(a9_wr[66]),  .coef_in(coef[0]), .rdup_out(a10_wr[64]), .rdlo_out(a10_wr[66]));
			radix2 #(.width(width)) rd_st9_65  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[65]), .rdlo_in(a9_wr[67]),  .coef_in(coef[512]), .rdup_out(a10_wr[65]), .rdlo_out(a10_wr[67]));
			radix2 #(.width(width)) rd_st9_68  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[68]), .rdlo_in(a9_wr[70]),  .coef_in(coef[0]), .rdup_out(a10_wr[68]), .rdlo_out(a10_wr[70]));
			radix2 #(.width(width)) rd_st9_69  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[69]), .rdlo_in(a9_wr[71]),  .coef_in(coef[512]), .rdup_out(a10_wr[69]), .rdlo_out(a10_wr[71]));
			radix2 #(.width(width)) rd_st9_72  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[72]), .rdlo_in(a9_wr[74]),  .coef_in(coef[0]), .rdup_out(a10_wr[72]), .rdlo_out(a10_wr[74]));
			radix2 #(.width(width)) rd_st9_73  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[73]), .rdlo_in(a9_wr[75]),  .coef_in(coef[512]), .rdup_out(a10_wr[73]), .rdlo_out(a10_wr[75]));
			radix2 #(.width(width)) rd_st9_76  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[76]), .rdlo_in(a9_wr[78]),  .coef_in(coef[0]), .rdup_out(a10_wr[76]), .rdlo_out(a10_wr[78]));
			radix2 #(.width(width)) rd_st9_77  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[77]), .rdlo_in(a9_wr[79]),  .coef_in(coef[512]), .rdup_out(a10_wr[77]), .rdlo_out(a10_wr[79]));
			radix2 #(.width(width)) rd_st9_80  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[80]), .rdlo_in(a9_wr[82]),  .coef_in(coef[0]), .rdup_out(a10_wr[80]), .rdlo_out(a10_wr[82]));
			radix2 #(.width(width)) rd_st9_81  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[81]), .rdlo_in(a9_wr[83]),  .coef_in(coef[512]), .rdup_out(a10_wr[81]), .rdlo_out(a10_wr[83]));
			radix2 #(.width(width)) rd_st9_84  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[84]), .rdlo_in(a9_wr[86]),  .coef_in(coef[0]), .rdup_out(a10_wr[84]), .rdlo_out(a10_wr[86]));
			radix2 #(.width(width)) rd_st9_85  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[85]), .rdlo_in(a9_wr[87]),  .coef_in(coef[512]), .rdup_out(a10_wr[85]), .rdlo_out(a10_wr[87]));
			radix2 #(.width(width)) rd_st9_88  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[88]), .rdlo_in(a9_wr[90]),  .coef_in(coef[0]), .rdup_out(a10_wr[88]), .rdlo_out(a10_wr[90]));
			radix2 #(.width(width)) rd_st9_89  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[89]), .rdlo_in(a9_wr[91]),  .coef_in(coef[512]), .rdup_out(a10_wr[89]), .rdlo_out(a10_wr[91]));
			radix2 #(.width(width)) rd_st9_92  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[92]), .rdlo_in(a9_wr[94]),  .coef_in(coef[0]), .rdup_out(a10_wr[92]), .rdlo_out(a10_wr[94]));
			radix2 #(.width(width)) rd_st9_93  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[93]), .rdlo_in(a9_wr[95]),  .coef_in(coef[512]), .rdup_out(a10_wr[93]), .rdlo_out(a10_wr[95]));
			radix2 #(.width(width)) rd_st9_96  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[96]), .rdlo_in(a9_wr[98]),  .coef_in(coef[0]), .rdup_out(a10_wr[96]), .rdlo_out(a10_wr[98]));
			radix2 #(.width(width)) rd_st9_97  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[97]), .rdlo_in(a9_wr[99]),  .coef_in(coef[512]), .rdup_out(a10_wr[97]), .rdlo_out(a10_wr[99]));
			radix2 #(.width(width)) rd_st9_100  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[100]), .rdlo_in(a9_wr[102]),  .coef_in(coef[0]), .rdup_out(a10_wr[100]), .rdlo_out(a10_wr[102]));
			radix2 #(.width(width)) rd_st9_101  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[101]), .rdlo_in(a9_wr[103]),  .coef_in(coef[512]), .rdup_out(a10_wr[101]), .rdlo_out(a10_wr[103]));
			radix2 #(.width(width)) rd_st9_104  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[104]), .rdlo_in(a9_wr[106]),  .coef_in(coef[0]), .rdup_out(a10_wr[104]), .rdlo_out(a10_wr[106]));
			radix2 #(.width(width)) rd_st9_105  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[105]), .rdlo_in(a9_wr[107]),  .coef_in(coef[512]), .rdup_out(a10_wr[105]), .rdlo_out(a10_wr[107]));
			radix2 #(.width(width)) rd_st9_108  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[108]), .rdlo_in(a9_wr[110]),  .coef_in(coef[0]), .rdup_out(a10_wr[108]), .rdlo_out(a10_wr[110]));
			radix2 #(.width(width)) rd_st9_109  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[109]), .rdlo_in(a9_wr[111]),  .coef_in(coef[512]), .rdup_out(a10_wr[109]), .rdlo_out(a10_wr[111]));
			radix2 #(.width(width)) rd_st9_112  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[112]), .rdlo_in(a9_wr[114]),  .coef_in(coef[0]), .rdup_out(a10_wr[112]), .rdlo_out(a10_wr[114]));
			radix2 #(.width(width)) rd_st9_113  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[113]), .rdlo_in(a9_wr[115]),  .coef_in(coef[512]), .rdup_out(a10_wr[113]), .rdlo_out(a10_wr[115]));
			radix2 #(.width(width)) rd_st9_116  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[116]), .rdlo_in(a9_wr[118]),  .coef_in(coef[0]), .rdup_out(a10_wr[116]), .rdlo_out(a10_wr[118]));
			radix2 #(.width(width)) rd_st9_117  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[117]), .rdlo_in(a9_wr[119]),  .coef_in(coef[512]), .rdup_out(a10_wr[117]), .rdlo_out(a10_wr[119]));
			radix2 #(.width(width)) rd_st9_120  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[120]), .rdlo_in(a9_wr[122]),  .coef_in(coef[0]), .rdup_out(a10_wr[120]), .rdlo_out(a10_wr[122]));
			radix2 #(.width(width)) rd_st9_121  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[121]), .rdlo_in(a9_wr[123]),  .coef_in(coef[512]), .rdup_out(a10_wr[121]), .rdlo_out(a10_wr[123]));
			radix2 #(.width(width)) rd_st9_124  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[124]), .rdlo_in(a9_wr[126]),  .coef_in(coef[0]), .rdup_out(a10_wr[124]), .rdlo_out(a10_wr[126]));
			radix2 #(.width(width)) rd_st9_125  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[125]), .rdlo_in(a9_wr[127]),  .coef_in(coef[512]), .rdup_out(a10_wr[125]), .rdlo_out(a10_wr[127]));
			radix2 #(.width(width)) rd_st9_128  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[128]), .rdlo_in(a9_wr[130]),  .coef_in(coef[0]), .rdup_out(a10_wr[128]), .rdlo_out(a10_wr[130]));
			radix2 #(.width(width)) rd_st9_129  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[129]), .rdlo_in(a9_wr[131]),  .coef_in(coef[512]), .rdup_out(a10_wr[129]), .rdlo_out(a10_wr[131]));
			radix2 #(.width(width)) rd_st9_132  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[132]), .rdlo_in(a9_wr[134]),  .coef_in(coef[0]), .rdup_out(a10_wr[132]), .rdlo_out(a10_wr[134]));
			radix2 #(.width(width)) rd_st9_133  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[133]), .rdlo_in(a9_wr[135]),  .coef_in(coef[512]), .rdup_out(a10_wr[133]), .rdlo_out(a10_wr[135]));
			radix2 #(.width(width)) rd_st9_136  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[136]), .rdlo_in(a9_wr[138]),  .coef_in(coef[0]), .rdup_out(a10_wr[136]), .rdlo_out(a10_wr[138]));
			radix2 #(.width(width)) rd_st9_137  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[137]), .rdlo_in(a9_wr[139]),  .coef_in(coef[512]), .rdup_out(a10_wr[137]), .rdlo_out(a10_wr[139]));
			radix2 #(.width(width)) rd_st9_140  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[140]), .rdlo_in(a9_wr[142]),  .coef_in(coef[0]), .rdup_out(a10_wr[140]), .rdlo_out(a10_wr[142]));
			radix2 #(.width(width)) rd_st9_141  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[141]), .rdlo_in(a9_wr[143]),  .coef_in(coef[512]), .rdup_out(a10_wr[141]), .rdlo_out(a10_wr[143]));
			radix2 #(.width(width)) rd_st9_144  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[144]), .rdlo_in(a9_wr[146]),  .coef_in(coef[0]), .rdup_out(a10_wr[144]), .rdlo_out(a10_wr[146]));
			radix2 #(.width(width)) rd_st9_145  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[145]), .rdlo_in(a9_wr[147]),  .coef_in(coef[512]), .rdup_out(a10_wr[145]), .rdlo_out(a10_wr[147]));
			radix2 #(.width(width)) rd_st9_148  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[148]), .rdlo_in(a9_wr[150]),  .coef_in(coef[0]), .rdup_out(a10_wr[148]), .rdlo_out(a10_wr[150]));
			radix2 #(.width(width)) rd_st9_149  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[149]), .rdlo_in(a9_wr[151]),  .coef_in(coef[512]), .rdup_out(a10_wr[149]), .rdlo_out(a10_wr[151]));
			radix2 #(.width(width)) rd_st9_152  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[152]), .rdlo_in(a9_wr[154]),  .coef_in(coef[0]), .rdup_out(a10_wr[152]), .rdlo_out(a10_wr[154]));
			radix2 #(.width(width)) rd_st9_153  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[153]), .rdlo_in(a9_wr[155]),  .coef_in(coef[512]), .rdup_out(a10_wr[153]), .rdlo_out(a10_wr[155]));
			radix2 #(.width(width)) rd_st9_156  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[156]), .rdlo_in(a9_wr[158]),  .coef_in(coef[0]), .rdup_out(a10_wr[156]), .rdlo_out(a10_wr[158]));
			radix2 #(.width(width)) rd_st9_157  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[157]), .rdlo_in(a9_wr[159]),  .coef_in(coef[512]), .rdup_out(a10_wr[157]), .rdlo_out(a10_wr[159]));
			radix2 #(.width(width)) rd_st9_160  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[160]), .rdlo_in(a9_wr[162]),  .coef_in(coef[0]), .rdup_out(a10_wr[160]), .rdlo_out(a10_wr[162]));
			radix2 #(.width(width)) rd_st9_161  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[161]), .rdlo_in(a9_wr[163]),  .coef_in(coef[512]), .rdup_out(a10_wr[161]), .rdlo_out(a10_wr[163]));
			radix2 #(.width(width)) rd_st9_164  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[164]), .rdlo_in(a9_wr[166]),  .coef_in(coef[0]), .rdup_out(a10_wr[164]), .rdlo_out(a10_wr[166]));
			radix2 #(.width(width)) rd_st9_165  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[165]), .rdlo_in(a9_wr[167]),  .coef_in(coef[512]), .rdup_out(a10_wr[165]), .rdlo_out(a10_wr[167]));
			radix2 #(.width(width)) rd_st9_168  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[168]), .rdlo_in(a9_wr[170]),  .coef_in(coef[0]), .rdup_out(a10_wr[168]), .rdlo_out(a10_wr[170]));
			radix2 #(.width(width)) rd_st9_169  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[169]), .rdlo_in(a9_wr[171]),  .coef_in(coef[512]), .rdup_out(a10_wr[169]), .rdlo_out(a10_wr[171]));
			radix2 #(.width(width)) rd_st9_172  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[172]), .rdlo_in(a9_wr[174]),  .coef_in(coef[0]), .rdup_out(a10_wr[172]), .rdlo_out(a10_wr[174]));
			radix2 #(.width(width)) rd_st9_173  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[173]), .rdlo_in(a9_wr[175]),  .coef_in(coef[512]), .rdup_out(a10_wr[173]), .rdlo_out(a10_wr[175]));
			radix2 #(.width(width)) rd_st9_176  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[176]), .rdlo_in(a9_wr[178]),  .coef_in(coef[0]), .rdup_out(a10_wr[176]), .rdlo_out(a10_wr[178]));
			radix2 #(.width(width)) rd_st9_177  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[177]), .rdlo_in(a9_wr[179]),  .coef_in(coef[512]), .rdup_out(a10_wr[177]), .rdlo_out(a10_wr[179]));
			radix2 #(.width(width)) rd_st9_180  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[180]), .rdlo_in(a9_wr[182]),  .coef_in(coef[0]), .rdup_out(a10_wr[180]), .rdlo_out(a10_wr[182]));
			radix2 #(.width(width)) rd_st9_181  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[181]), .rdlo_in(a9_wr[183]),  .coef_in(coef[512]), .rdup_out(a10_wr[181]), .rdlo_out(a10_wr[183]));
			radix2 #(.width(width)) rd_st9_184  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[184]), .rdlo_in(a9_wr[186]),  .coef_in(coef[0]), .rdup_out(a10_wr[184]), .rdlo_out(a10_wr[186]));
			radix2 #(.width(width)) rd_st9_185  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[185]), .rdlo_in(a9_wr[187]),  .coef_in(coef[512]), .rdup_out(a10_wr[185]), .rdlo_out(a10_wr[187]));
			radix2 #(.width(width)) rd_st9_188  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[188]), .rdlo_in(a9_wr[190]),  .coef_in(coef[0]), .rdup_out(a10_wr[188]), .rdlo_out(a10_wr[190]));
			radix2 #(.width(width)) rd_st9_189  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[189]), .rdlo_in(a9_wr[191]),  .coef_in(coef[512]), .rdup_out(a10_wr[189]), .rdlo_out(a10_wr[191]));
			radix2 #(.width(width)) rd_st9_192  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[192]), .rdlo_in(a9_wr[194]),  .coef_in(coef[0]), .rdup_out(a10_wr[192]), .rdlo_out(a10_wr[194]));
			radix2 #(.width(width)) rd_st9_193  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[193]), .rdlo_in(a9_wr[195]),  .coef_in(coef[512]), .rdup_out(a10_wr[193]), .rdlo_out(a10_wr[195]));
			radix2 #(.width(width)) rd_st9_196  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[196]), .rdlo_in(a9_wr[198]),  .coef_in(coef[0]), .rdup_out(a10_wr[196]), .rdlo_out(a10_wr[198]));
			radix2 #(.width(width)) rd_st9_197  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[197]), .rdlo_in(a9_wr[199]),  .coef_in(coef[512]), .rdup_out(a10_wr[197]), .rdlo_out(a10_wr[199]));
			radix2 #(.width(width)) rd_st9_200  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[200]), .rdlo_in(a9_wr[202]),  .coef_in(coef[0]), .rdup_out(a10_wr[200]), .rdlo_out(a10_wr[202]));
			radix2 #(.width(width)) rd_st9_201  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[201]), .rdlo_in(a9_wr[203]),  .coef_in(coef[512]), .rdup_out(a10_wr[201]), .rdlo_out(a10_wr[203]));
			radix2 #(.width(width)) rd_st9_204  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[204]), .rdlo_in(a9_wr[206]),  .coef_in(coef[0]), .rdup_out(a10_wr[204]), .rdlo_out(a10_wr[206]));
			radix2 #(.width(width)) rd_st9_205  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[205]), .rdlo_in(a9_wr[207]),  .coef_in(coef[512]), .rdup_out(a10_wr[205]), .rdlo_out(a10_wr[207]));
			radix2 #(.width(width)) rd_st9_208  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[208]), .rdlo_in(a9_wr[210]),  .coef_in(coef[0]), .rdup_out(a10_wr[208]), .rdlo_out(a10_wr[210]));
			radix2 #(.width(width)) rd_st9_209  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[209]), .rdlo_in(a9_wr[211]),  .coef_in(coef[512]), .rdup_out(a10_wr[209]), .rdlo_out(a10_wr[211]));
			radix2 #(.width(width)) rd_st9_212  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[212]), .rdlo_in(a9_wr[214]),  .coef_in(coef[0]), .rdup_out(a10_wr[212]), .rdlo_out(a10_wr[214]));
			radix2 #(.width(width)) rd_st9_213  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[213]), .rdlo_in(a9_wr[215]),  .coef_in(coef[512]), .rdup_out(a10_wr[213]), .rdlo_out(a10_wr[215]));
			radix2 #(.width(width)) rd_st9_216  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[216]), .rdlo_in(a9_wr[218]),  .coef_in(coef[0]), .rdup_out(a10_wr[216]), .rdlo_out(a10_wr[218]));
			radix2 #(.width(width)) rd_st9_217  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[217]), .rdlo_in(a9_wr[219]),  .coef_in(coef[512]), .rdup_out(a10_wr[217]), .rdlo_out(a10_wr[219]));
			radix2 #(.width(width)) rd_st9_220  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[220]), .rdlo_in(a9_wr[222]),  .coef_in(coef[0]), .rdup_out(a10_wr[220]), .rdlo_out(a10_wr[222]));
			radix2 #(.width(width)) rd_st9_221  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[221]), .rdlo_in(a9_wr[223]),  .coef_in(coef[512]), .rdup_out(a10_wr[221]), .rdlo_out(a10_wr[223]));
			radix2 #(.width(width)) rd_st9_224  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[224]), .rdlo_in(a9_wr[226]),  .coef_in(coef[0]), .rdup_out(a10_wr[224]), .rdlo_out(a10_wr[226]));
			radix2 #(.width(width)) rd_st9_225  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[225]), .rdlo_in(a9_wr[227]),  .coef_in(coef[512]), .rdup_out(a10_wr[225]), .rdlo_out(a10_wr[227]));
			radix2 #(.width(width)) rd_st9_228  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[228]), .rdlo_in(a9_wr[230]),  .coef_in(coef[0]), .rdup_out(a10_wr[228]), .rdlo_out(a10_wr[230]));
			radix2 #(.width(width)) rd_st9_229  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[229]), .rdlo_in(a9_wr[231]),  .coef_in(coef[512]), .rdup_out(a10_wr[229]), .rdlo_out(a10_wr[231]));
			radix2 #(.width(width)) rd_st9_232  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[232]), .rdlo_in(a9_wr[234]),  .coef_in(coef[0]), .rdup_out(a10_wr[232]), .rdlo_out(a10_wr[234]));
			radix2 #(.width(width)) rd_st9_233  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[233]), .rdlo_in(a9_wr[235]),  .coef_in(coef[512]), .rdup_out(a10_wr[233]), .rdlo_out(a10_wr[235]));
			radix2 #(.width(width)) rd_st9_236  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[236]), .rdlo_in(a9_wr[238]),  .coef_in(coef[0]), .rdup_out(a10_wr[236]), .rdlo_out(a10_wr[238]));
			radix2 #(.width(width)) rd_st9_237  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[237]), .rdlo_in(a9_wr[239]),  .coef_in(coef[512]), .rdup_out(a10_wr[237]), .rdlo_out(a10_wr[239]));
			radix2 #(.width(width)) rd_st9_240  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[240]), .rdlo_in(a9_wr[242]),  .coef_in(coef[0]), .rdup_out(a10_wr[240]), .rdlo_out(a10_wr[242]));
			radix2 #(.width(width)) rd_st9_241  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[241]), .rdlo_in(a9_wr[243]),  .coef_in(coef[512]), .rdup_out(a10_wr[241]), .rdlo_out(a10_wr[243]));
			radix2 #(.width(width)) rd_st9_244  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[244]), .rdlo_in(a9_wr[246]),  .coef_in(coef[0]), .rdup_out(a10_wr[244]), .rdlo_out(a10_wr[246]));
			radix2 #(.width(width)) rd_st9_245  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[245]), .rdlo_in(a9_wr[247]),  .coef_in(coef[512]), .rdup_out(a10_wr[245]), .rdlo_out(a10_wr[247]));
			radix2 #(.width(width)) rd_st9_248  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[248]), .rdlo_in(a9_wr[250]),  .coef_in(coef[0]), .rdup_out(a10_wr[248]), .rdlo_out(a10_wr[250]));
			radix2 #(.width(width)) rd_st9_249  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[249]), .rdlo_in(a9_wr[251]),  .coef_in(coef[512]), .rdup_out(a10_wr[249]), .rdlo_out(a10_wr[251]));
			radix2 #(.width(width)) rd_st9_252  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[252]), .rdlo_in(a9_wr[254]),  .coef_in(coef[0]), .rdup_out(a10_wr[252]), .rdlo_out(a10_wr[254]));
			radix2 #(.width(width)) rd_st9_253  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[253]), .rdlo_in(a9_wr[255]),  .coef_in(coef[512]), .rdup_out(a10_wr[253]), .rdlo_out(a10_wr[255]));
			radix2 #(.width(width)) rd_st9_256  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[256]), .rdlo_in(a9_wr[258]),  .coef_in(coef[0]), .rdup_out(a10_wr[256]), .rdlo_out(a10_wr[258]));
			radix2 #(.width(width)) rd_st9_257  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[257]), .rdlo_in(a9_wr[259]),  .coef_in(coef[512]), .rdup_out(a10_wr[257]), .rdlo_out(a10_wr[259]));
			radix2 #(.width(width)) rd_st9_260  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[260]), .rdlo_in(a9_wr[262]),  .coef_in(coef[0]), .rdup_out(a10_wr[260]), .rdlo_out(a10_wr[262]));
			radix2 #(.width(width)) rd_st9_261  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[261]), .rdlo_in(a9_wr[263]),  .coef_in(coef[512]), .rdup_out(a10_wr[261]), .rdlo_out(a10_wr[263]));
			radix2 #(.width(width)) rd_st9_264  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[264]), .rdlo_in(a9_wr[266]),  .coef_in(coef[0]), .rdup_out(a10_wr[264]), .rdlo_out(a10_wr[266]));
			radix2 #(.width(width)) rd_st9_265  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[265]), .rdlo_in(a9_wr[267]),  .coef_in(coef[512]), .rdup_out(a10_wr[265]), .rdlo_out(a10_wr[267]));
			radix2 #(.width(width)) rd_st9_268  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[268]), .rdlo_in(a9_wr[270]),  .coef_in(coef[0]), .rdup_out(a10_wr[268]), .rdlo_out(a10_wr[270]));
			radix2 #(.width(width)) rd_st9_269  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[269]), .rdlo_in(a9_wr[271]),  .coef_in(coef[512]), .rdup_out(a10_wr[269]), .rdlo_out(a10_wr[271]));
			radix2 #(.width(width)) rd_st9_272  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[272]), .rdlo_in(a9_wr[274]),  .coef_in(coef[0]), .rdup_out(a10_wr[272]), .rdlo_out(a10_wr[274]));
			radix2 #(.width(width)) rd_st9_273  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[273]), .rdlo_in(a9_wr[275]),  .coef_in(coef[512]), .rdup_out(a10_wr[273]), .rdlo_out(a10_wr[275]));
			radix2 #(.width(width)) rd_st9_276  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[276]), .rdlo_in(a9_wr[278]),  .coef_in(coef[0]), .rdup_out(a10_wr[276]), .rdlo_out(a10_wr[278]));
			radix2 #(.width(width)) rd_st9_277  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[277]), .rdlo_in(a9_wr[279]),  .coef_in(coef[512]), .rdup_out(a10_wr[277]), .rdlo_out(a10_wr[279]));
			radix2 #(.width(width)) rd_st9_280  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[280]), .rdlo_in(a9_wr[282]),  .coef_in(coef[0]), .rdup_out(a10_wr[280]), .rdlo_out(a10_wr[282]));
			radix2 #(.width(width)) rd_st9_281  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[281]), .rdlo_in(a9_wr[283]),  .coef_in(coef[512]), .rdup_out(a10_wr[281]), .rdlo_out(a10_wr[283]));
			radix2 #(.width(width)) rd_st9_284  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[284]), .rdlo_in(a9_wr[286]),  .coef_in(coef[0]), .rdup_out(a10_wr[284]), .rdlo_out(a10_wr[286]));
			radix2 #(.width(width)) rd_st9_285  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[285]), .rdlo_in(a9_wr[287]),  .coef_in(coef[512]), .rdup_out(a10_wr[285]), .rdlo_out(a10_wr[287]));
			radix2 #(.width(width)) rd_st9_288  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[288]), .rdlo_in(a9_wr[290]),  .coef_in(coef[0]), .rdup_out(a10_wr[288]), .rdlo_out(a10_wr[290]));
			radix2 #(.width(width)) rd_st9_289  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[289]), .rdlo_in(a9_wr[291]),  .coef_in(coef[512]), .rdup_out(a10_wr[289]), .rdlo_out(a10_wr[291]));
			radix2 #(.width(width)) rd_st9_292  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[292]), .rdlo_in(a9_wr[294]),  .coef_in(coef[0]), .rdup_out(a10_wr[292]), .rdlo_out(a10_wr[294]));
			radix2 #(.width(width)) rd_st9_293  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[293]), .rdlo_in(a9_wr[295]),  .coef_in(coef[512]), .rdup_out(a10_wr[293]), .rdlo_out(a10_wr[295]));
			radix2 #(.width(width)) rd_st9_296  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[296]), .rdlo_in(a9_wr[298]),  .coef_in(coef[0]), .rdup_out(a10_wr[296]), .rdlo_out(a10_wr[298]));
			radix2 #(.width(width)) rd_st9_297  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[297]), .rdlo_in(a9_wr[299]),  .coef_in(coef[512]), .rdup_out(a10_wr[297]), .rdlo_out(a10_wr[299]));
			radix2 #(.width(width)) rd_st9_300  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[300]), .rdlo_in(a9_wr[302]),  .coef_in(coef[0]), .rdup_out(a10_wr[300]), .rdlo_out(a10_wr[302]));
			radix2 #(.width(width)) rd_st9_301  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[301]), .rdlo_in(a9_wr[303]),  .coef_in(coef[512]), .rdup_out(a10_wr[301]), .rdlo_out(a10_wr[303]));
			radix2 #(.width(width)) rd_st9_304  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[304]), .rdlo_in(a9_wr[306]),  .coef_in(coef[0]), .rdup_out(a10_wr[304]), .rdlo_out(a10_wr[306]));
			radix2 #(.width(width)) rd_st9_305  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[305]), .rdlo_in(a9_wr[307]),  .coef_in(coef[512]), .rdup_out(a10_wr[305]), .rdlo_out(a10_wr[307]));
			radix2 #(.width(width)) rd_st9_308  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[308]), .rdlo_in(a9_wr[310]),  .coef_in(coef[0]), .rdup_out(a10_wr[308]), .rdlo_out(a10_wr[310]));
			radix2 #(.width(width)) rd_st9_309  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[309]), .rdlo_in(a9_wr[311]),  .coef_in(coef[512]), .rdup_out(a10_wr[309]), .rdlo_out(a10_wr[311]));
			radix2 #(.width(width)) rd_st9_312  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[312]), .rdlo_in(a9_wr[314]),  .coef_in(coef[0]), .rdup_out(a10_wr[312]), .rdlo_out(a10_wr[314]));
			radix2 #(.width(width)) rd_st9_313  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[313]), .rdlo_in(a9_wr[315]),  .coef_in(coef[512]), .rdup_out(a10_wr[313]), .rdlo_out(a10_wr[315]));
			radix2 #(.width(width)) rd_st9_316  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[316]), .rdlo_in(a9_wr[318]),  .coef_in(coef[0]), .rdup_out(a10_wr[316]), .rdlo_out(a10_wr[318]));
			radix2 #(.width(width)) rd_st9_317  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[317]), .rdlo_in(a9_wr[319]),  .coef_in(coef[512]), .rdup_out(a10_wr[317]), .rdlo_out(a10_wr[319]));
			radix2 #(.width(width)) rd_st9_320  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[320]), .rdlo_in(a9_wr[322]),  .coef_in(coef[0]), .rdup_out(a10_wr[320]), .rdlo_out(a10_wr[322]));
			radix2 #(.width(width)) rd_st9_321  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[321]), .rdlo_in(a9_wr[323]),  .coef_in(coef[512]), .rdup_out(a10_wr[321]), .rdlo_out(a10_wr[323]));
			radix2 #(.width(width)) rd_st9_324  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[324]), .rdlo_in(a9_wr[326]),  .coef_in(coef[0]), .rdup_out(a10_wr[324]), .rdlo_out(a10_wr[326]));
			radix2 #(.width(width)) rd_st9_325  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[325]), .rdlo_in(a9_wr[327]),  .coef_in(coef[512]), .rdup_out(a10_wr[325]), .rdlo_out(a10_wr[327]));
			radix2 #(.width(width)) rd_st9_328  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[328]), .rdlo_in(a9_wr[330]),  .coef_in(coef[0]), .rdup_out(a10_wr[328]), .rdlo_out(a10_wr[330]));
			radix2 #(.width(width)) rd_st9_329  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[329]), .rdlo_in(a9_wr[331]),  .coef_in(coef[512]), .rdup_out(a10_wr[329]), .rdlo_out(a10_wr[331]));
			radix2 #(.width(width)) rd_st9_332  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[332]), .rdlo_in(a9_wr[334]),  .coef_in(coef[0]), .rdup_out(a10_wr[332]), .rdlo_out(a10_wr[334]));
			radix2 #(.width(width)) rd_st9_333  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[333]), .rdlo_in(a9_wr[335]),  .coef_in(coef[512]), .rdup_out(a10_wr[333]), .rdlo_out(a10_wr[335]));
			radix2 #(.width(width)) rd_st9_336  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[336]), .rdlo_in(a9_wr[338]),  .coef_in(coef[0]), .rdup_out(a10_wr[336]), .rdlo_out(a10_wr[338]));
			radix2 #(.width(width)) rd_st9_337  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[337]), .rdlo_in(a9_wr[339]),  .coef_in(coef[512]), .rdup_out(a10_wr[337]), .rdlo_out(a10_wr[339]));
			radix2 #(.width(width)) rd_st9_340  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[340]), .rdlo_in(a9_wr[342]),  .coef_in(coef[0]), .rdup_out(a10_wr[340]), .rdlo_out(a10_wr[342]));
			radix2 #(.width(width)) rd_st9_341  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[341]), .rdlo_in(a9_wr[343]),  .coef_in(coef[512]), .rdup_out(a10_wr[341]), .rdlo_out(a10_wr[343]));
			radix2 #(.width(width)) rd_st9_344  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[344]), .rdlo_in(a9_wr[346]),  .coef_in(coef[0]), .rdup_out(a10_wr[344]), .rdlo_out(a10_wr[346]));
			radix2 #(.width(width)) rd_st9_345  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[345]), .rdlo_in(a9_wr[347]),  .coef_in(coef[512]), .rdup_out(a10_wr[345]), .rdlo_out(a10_wr[347]));
			radix2 #(.width(width)) rd_st9_348  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[348]), .rdlo_in(a9_wr[350]),  .coef_in(coef[0]), .rdup_out(a10_wr[348]), .rdlo_out(a10_wr[350]));
			radix2 #(.width(width)) rd_st9_349  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[349]), .rdlo_in(a9_wr[351]),  .coef_in(coef[512]), .rdup_out(a10_wr[349]), .rdlo_out(a10_wr[351]));
			radix2 #(.width(width)) rd_st9_352  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[352]), .rdlo_in(a9_wr[354]),  .coef_in(coef[0]), .rdup_out(a10_wr[352]), .rdlo_out(a10_wr[354]));
			radix2 #(.width(width)) rd_st9_353  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[353]), .rdlo_in(a9_wr[355]),  .coef_in(coef[512]), .rdup_out(a10_wr[353]), .rdlo_out(a10_wr[355]));
			radix2 #(.width(width)) rd_st9_356  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[356]), .rdlo_in(a9_wr[358]),  .coef_in(coef[0]), .rdup_out(a10_wr[356]), .rdlo_out(a10_wr[358]));
			radix2 #(.width(width)) rd_st9_357  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[357]), .rdlo_in(a9_wr[359]),  .coef_in(coef[512]), .rdup_out(a10_wr[357]), .rdlo_out(a10_wr[359]));
			radix2 #(.width(width)) rd_st9_360  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[360]), .rdlo_in(a9_wr[362]),  .coef_in(coef[0]), .rdup_out(a10_wr[360]), .rdlo_out(a10_wr[362]));
			radix2 #(.width(width)) rd_st9_361  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[361]), .rdlo_in(a9_wr[363]),  .coef_in(coef[512]), .rdup_out(a10_wr[361]), .rdlo_out(a10_wr[363]));
			radix2 #(.width(width)) rd_st9_364  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[364]), .rdlo_in(a9_wr[366]),  .coef_in(coef[0]), .rdup_out(a10_wr[364]), .rdlo_out(a10_wr[366]));
			radix2 #(.width(width)) rd_st9_365  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[365]), .rdlo_in(a9_wr[367]),  .coef_in(coef[512]), .rdup_out(a10_wr[365]), .rdlo_out(a10_wr[367]));
			radix2 #(.width(width)) rd_st9_368  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[368]), .rdlo_in(a9_wr[370]),  .coef_in(coef[0]), .rdup_out(a10_wr[368]), .rdlo_out(a10_wr[370]));
			radix2 #(.width(width)) rd_st9_369  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[369]), .rdlo_in(a9_wr[371]),  .coef_in(coef[512]), .rdup_out(a10_wr[369]), .rdlo_out(a10_wr[371]));
			radix2 #(.width(width)) rd_st9_372  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[372]), .rdlo_in(a9_wr[374]),  .coef_in(coef[0]), .rdup_out(a10_wr[372]), .rdlo_out(a10_wr[374]));
			radix2 #(.width(width)) rd_st9_373  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[373]), .rdlo_in(a9_wr[375]),  .coef_in(coef[512]), .rdup_out(a10_wr[373]), .rdlo_out(a10_wr[375]));
			radix2 #(.width(width)) rd_st9_376  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[376]), .rdlo_in(a9_wr[378]),  .coef_in(coef[0]), .rdup_out(a10_wr[376]), .rdlo_out(a10_wr[378]));
			radix2 #(.width(width)) rd_st9_377  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[377]), .rdlo_in(a9_wr[379]),  .coef_in(coef[512]), .rdup_out(a10_wr[377]), .rdlo_out(a10_wr[379]));
			radix2 #(.width(width)) rd_st9_380  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[380]), .rdlo_in(a9_wr[382]),  .coef_in(coef[0]), .rdup_out(a10_wr[380]), .rdlo_out(a10_wr[382]));
			radix2 #(.width(width)) rd_st9_381  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[381]), .rdlo_in(a9_wr[383]),  .coef_in(coef[512]), .rdup_out(a10_wr[381]), .rdlo_out(a10_wr[383]));
			radix2 #(.width(width)) rd_st9_384  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[384]), .rdlo_in(a9_wr[386]),  .coef_in(coef[0]), .rdup_out(a10_wr[384]), .rdlo_out(a10_wr[386]));
			radix2 #(.width(width)) rd_st9_385  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[385]), .rdlo_in(a9_wr[387]),  .coef_in(coef[512]), .rdup_out(a10_wr[385]), .rdlo_out(a10_wr[387]));
			radix2 #(.width(width)) rd_st9_388  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[388]), .rdlo_in(a9_wr[390]),  .coef_in(coef[0]), .rdup_out(a10_wr[388]), .rdlo_out(a10_wr[390]));
			radix2 #(.width(width)) rd_st9_389  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[389]), .rdlo_in(a9_wr[391]),  .coef_in(coef[512]), .rdup_out(a10_wr[389]), .rdlo_out(a10_wr[391]));
			radix2 #(.width(width)) rd_st9_392  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[392]), .rdlo_in(a9_wr[394]),  .coef_in(coef[0]), .rdup_out(a10_wr[392]), .rdlo_out(a10_wr[394]));
			radix2 #(.width(width)) rd_st9_393  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[393]), .rdlo_in(a9_wr[395]),  .coef_in(coef[512]), .rdup_out(a10_wr[393]), .rdlo_out(a10_wr[395]));
			radix2 #(.width(width)) rd_st9_396  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[396]), .rdlo_in(a9_wr[398]),  .coef_in(coef[0]), .rdup_out(a10_wr[396]), .rdlo_out(a10_wr[398]));
			radix2 #(.width(width)) rd_st9_397  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[397]), .rdlo_in(a9_wr[399]),  .coef_in(coef[512]), .rdup_out(a10_wr[397]), .rdlo_out(a10_wr[399]));
			radix2 #(.width(width)) rd_st9_400  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[400]), .rdlo_in(a9_wr[402]),  .coef_in(coef[0]), .rdup_out(a10_wr[400]), .rdlo_out(a10_wr[402]));
			radix2 #(.width(width)) rd_st9_401  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[401]), .rdlo_in(a9_wr[403]),  .coef_in(coef[512]), .rdup_out(a10_wr[401]), .rdlo_out(a10_wr[403]));
			radix2 #(.width(width)) rd_st9_404  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[404]), .rdlo_in(a9_wr[406]),  .coef_in(coef[0]), .rdup_out(a10_wr[404]), .rdlo_out(a10_wr[406]));
			radix2 #(.width(width)) rd_st9_405  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[405]), .rdlo_in(a9_wr[407]),  .coef_in(coef[512]), .rdup_out(a10_wr[405]), .rdlo_out(a10_wr[407]));
			radix2 #(.width(width)) rd_st9_408  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[408]), .rdlo_in(a9_wr[410]),  .coef_in(coef[0]), .rdup_out(a10_wr[408]), .rdlo_out(a10_wr[410]));
			radix2 #(.width(width)) rd_st9_409  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[409]), .rdlo_in(a9_wr[411]),  .coef_in(coef[512]), .rdup_out(a10_wr[409]), .rdlo_out(a10_wr[411]));
			radix2 #(.width(width)) rd_st9_412  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[412]), .rdlo_in(a9_wr[414]),  .coef_in(coef[0]), .rdup_out(a10_wr[412]), .rdlo_out(a10_wr[414]));
			radix2 #(.width(width)) rd_st9_413  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[413]), .rdlo_in(a9_wr[415]),  .coef_in(coef[512]), .rdup_out(a10_wr[413]), .rdlo_out(a10_wr[415]));
			radix2 #(.width(width)) rd_st9_416  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[416]), .rdlo_in(a9_wr[418]),  .coef_in(coef[0]), .rdup_out(a10_wr[416]), .rdlo_out(a10_wr[418]));
			radix2 #(.width(width)) rd_st9_417  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[417]), .rdlo_in(a9_wr[419]),  .coef_in(coef[512]), .rdup_out(a10_wr[417]), .rdlo_out(a10_wr[419]));
			radix2 #(.width(width)) rd_st9_420  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[420]), .rdlo_in(a9_wr[422]),  .coef_in(coef[0]), .rdup_out(a10_wr[420]), .rdlo_out(a10_wr[422]));
			radix2 #(.width(width)) rd_st9_421  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[421]), .rdlo_in(a9_wr[423]),  .coef_in(coef[512]), .rdup_out(a10_wr[421]), .rdlo_out(a10_wr[423]));
			radix2 #(.width(width)) rd_st9_424  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[424]), .rdlo_in(a9_wr[426]),  .coef_in(coef[0]), .rdup_out(a10_wr[424]), .rdlo_out(a10_wr[426]));
			radix2 #(.width(width)) rd_st9_425  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[425]), .rdlo_in(a9_wr[427]),  .coef_in(coef[512]), .rdup_out(a10_wr[425]), .rdlo_out(a10_wr[427]));
			radix2 #(.width(width)) rd_st9_428  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[428]), .rdlo_in(a9_wr[430]),  .coef_in(coef[0]), .rdup_out(a10_wr[428]), .rdlo_out(a10_wr[430]));
			radix2 #(.width(width)) rd_st9_429  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[429]), .rdlo_in(a9_wr[431]),  .coef_in(coef[512]), .rdup_out(a10_wr[429]), .rdlo_out(a10_wr[431]));
			radix2 #(.width(width)) rd_st9_432  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[432]), .rdlo_in(a9_wr[434]),  .coef_in(coef[0]), .rdup_out(a10_wr[432]), .rdlo_out(a10_wr[434]));
			radix2 #(.width(width)) rd_st9_433  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[433]), .rdlo_in(a9_wr[435]),  .coef_in(coef[512]), .rdup_out(a10_wr[433]), .rdlo_out(a10_wr[435]));
			radix2 #(.width(width)) rd_st9_436  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[436]), .rdlo_in(a9_wr[438]),  .coef_in(coef[0]), .rdup_out(a10_wr[436]), .rdlo_out(a10_wr[438]));
			radix2 #(.width(width)) rd_st9_437  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[437]), .rdlo_in(a9_wr[439]),  .coef_in(coef[512]), .rdup_out(a10_wr[437]), .rdlo_out(a10_wr[439]));
			radix2 #(.width(width)) rd_st9_440  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[440]), .rdlo_in(a9_wr[442]),  .coef_in(coef[0]), .rdup_out(a10_wr[440]), .rdlo_out(a10_wr[442]));
			radix2 #(.width(width)) rd_st9_441  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[441]), .rdlo_in(a9_wr[443]),  .coef_in(coef[512]), .rdup_out(a10_wr[441]), .rdlo_out(a10_wr[443]));
			radix2 #(.width(width)) rd_st9_444  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[444]), .rdlo_in(a9_wr[446]),  .coef_in(coef[0]), .rdup_out(a10_wr[444]), .rdlo_out(a10_wr[446]));
			radix2 #(.width(width)) rd_st9_445  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[445]), .rdlo_in(a9_wr[447]),  .coef_in(coef[512]), .rdup_out(a10_wr[445]), .rdlo_out(a10_wr[447]));
			radix2 #(.width(width)) rd_st9_448  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[448]), .rdlo_in(a9_wr[450]),  .coef_in(coef[0]), .rdup_out(a10_wr[448]), .rdlo_out(a10_wr[450]));
			radix2 #(.width(width)) rd_st9_449  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[449]), .rdlo_in(a9_wr[451]),  .coef_in(coef[512]), .rdup_out(a10_wr[449]), .rdlo_out(a10_wr[451]));
			radix2 #(.width(width)) rd_st9_452  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[452]), .rdlo_in(a9_wr[454]),  .coef_in(coef[0]), .rdup_out(a10_wr[452]), .rdlo_out(a10_wr[454]));
			radix2 #(.width(width)) rd_st9_453  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[453]), .rdlo_in(a9_wr[455]),  .coef_in(coef[512]), .rdup_out(a10_wr[453]), .rdlo_out(a10_wr[455]));
			radix2 #(.width(width)) rd_st9_456  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[456]), .rdlo_in(a9_wr[458]),  .coef_in(coef[0]), .rdup_out(a10_wr[456]), .rdlo_out(a10_wr[458]));
			radix2 #(.width(width)) rd_st9_457  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[457]), .rdlo_in(a9_wr[459]),  .coef_in(coef[512]), .rdup_out(a10_wr[457]), .rdlo_out(a10_wr[459]));
			radix2 #(.width(width)) rd_st9_460  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[460]), .rdlo_in(a9_wr[462]),  .coef_in(coef[0]), .rdup_out(a10_wr[460]), .rdlo_out(a10_wr[462]));
			radix2 #(.width(width)) rd_st9_461  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[461]), .rdlo_in(a9_wr[463]),  .coef_in(coef[512]), .rdup_out(a10_wr[461]), .rdlo_out(a10_wr[463]));
			radix2 #(.width(width)) rd_st9_464  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[464]), .rdlo_in(a9_wr[466]),  .coef_in(coef[0]), .rdup_out(a10_wr[464]), .rdlo_out(a10_wr[466]));
			radix2 #(.width(width)) rd_st9_465  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[465]), .rdlo_in(a9_wr[467]),  .coef_in(coef[512]), .rdup_out(a10_wr[465]), .rdlo_out(a10_wr[467]));
			radix2 #(.width(width)) rd_st9_468  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[468]), .rdlo_in(a9_wr[470]),  .coef_in(coef[0]), .rdup_out(a10_wr[468]), .rdlo_out(a10_wr[470]));
			radix2 #(.width(width)) rd_st9_469  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[469]), .rdlo_in(a9_wr[471]),  .coef_in(coef[512]), .rdup_out(a10_wr[469]), .rdlo_out(a10_wr[471]));
			radix2 #(.width(width)) rd_st9_472  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[472]), .rdlo_in(a9_wr[474]),  .coef_in(coef[0]), .rdup_out(a10_wr[472]), .rdlo_out(a10_wr[474]));
			radix2 #(.width(width)) rd_st9_473  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[473]), .rdlo_in(a9_wr[475]),  .coef_in(coef[512]), .rdup_out(a10_wr[473]), .rdlo_out(a10_wr[475]));
			radix2 #(.width(width)) rd_st9_476  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[476]), .rdlo_in(a9_wr[478]),  .coef_in(coef[0]), .rdup_out(a10_wr[476]), .rdlo_out(a10_wr[478]));
			radix2 #(.width(width)) rd_st9_477  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[477]), .rdlo_in(a9_wr[479]),  .coef_in(coef[512]), .rdup_out(a10_wr[477]), .rdlo_out(a10_wr[479]));
			radix2 #(.width(width)) rd_st9_480  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[480]), .rdlo_in(a9_wr[482]),  .coef_in(coef[0]), .rdup_out(a10_wr[480]), .rdlo_out(a10_wr[482]));
			radix2 #(.width(width)) rd_st9_481  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[481]), .rdlo_in(a9_wr[483]),  .coef_in(coef[512]), .rdup_out(a10_wr[481]), .rdlo_out(a10_wr[483]));
			radix2 #(.width(width)) rd_st9_484  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[484]), .rdlo_in(a9_wr[486]),  .coef_in(coef[0]), .rdup_out(a10_wr[484]), .rdlo_out(a10_wr[486]));
			radix2 #(.width(width)) rd_st9_485  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[485]), .rdlo_in(a9_wr[487]),  .coef_in(coef[512]), .rdup_out(a10_wr[485]), .rdlo_out(a10_wr[487]));
			radix2 #(.width(width)) rd_st9_488  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[488]), .rdlo_in(a9_wr[490]),  .coef_in(coef[0]), .rdup_out(a10_wr[488]), .rdlo_out(a10_wr[490]));
			radix2 #(.width(width)) rd_st9_489  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[489]), .rdlo_in(a9_wr[491]),  .coef_in(coef[512]), .rdup_out(a10_wr[489]), .rdlo_out(a10_wr[491]));
			radix2 #(.width(width)) rd_st9_492  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[492]), .rdlo_in(a9_wr[494]),  .coef_in(coef[0]), .rdup_out(a10_wr[492]), .rdlo_out(a10_wr[494]));
			radix2 #(.width(width)) rd_st9_493  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[493]), .rdlo_in(a9_wr[495]),  .coef_in(coef[512]), .rdup_out(a10_wr[493]), .rdlo_out(a10_wr[495]));
			radix2 #(.width(width)) rd_st9_496  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[496]), .rdlo_in(a9_wr[498]),  .coef_in(coef[0]), .rdup_out(a10_wr[496]), .rdlo_out(a10_wr[498]));
			radix2 #(.width(width)) rd_st9_497  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[497]), .rdlo_in(a9_wr[499]),  .coef_in(coef[512]), .rdup_out(a10_wr[497]), .rdlo_out(a10_wr[499]));
			radix2 #(.width(width)) rd_st9_500  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[500]), .rdlo_in(a9_wr[502]),  .coef_in(coef[0]), .rdup_out(a10_wr[500]), .rdlo_out(a10_wr[502]));
			radix2 #(.width(width)) rd_st9_501  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[501]), .rdlo_in(a9_wr[503]),  .coef_in(coef[512]), .rdup_out(a10_wr[501]), .rdlo_out(a10_wr[503]));
			radix2 #(.width(width)) rd_st9_504  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[504]), .rdlo_in(a9_wr[506]),  .coef_in(coef[0]), .rdup_out(a10_wr[504]), .rdlo_out(a10_wr[506]));
			radix2 #(.width(width)) rd_st9_505  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[505]), .rdlo_in(a9_wr[507]),  .coef_in(coef[512]), .rdup_out(a10_wr[505]), .rdlo_out(a10_wr[507]));
			radix2 #(.width(width)) rd_st9_508  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[508]), .rdlo_in(a9_wr[510]),  .coef_in(coef[0]), .rdup_out(a10_wr[508]), .rdlo_out(a10_wr[510]));
			radix2 #(.width(width)) rd_st9_509  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[509]), .rdlo_in(a9_wr[511]),  .coef_in(coef[512]), .rdup_out(a10_wr[509]), .rdlo_out(a10_wr[511]));
			radix2 #(.width(width)) rd_st9_512  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[512]), .rdlo_in(a9_wr[514]),  .coef_in(coef[0]), .rdup_out(a10_wr[512]), .rdlo_out(a10_wr[514]));
			radix2 #(.width(width)) rd_st9_513  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[513]), .rdlo_in(a9_wr[515]),  .coef_in(coef[512]), .rdup_out(a10_wr[513]), .rdlo_out(a10_wr[515]));
			radix2 #(.width(width)) rd_st9_516  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[516]), .rdlo_in(a9_wr[518]),  .coef_in(coef[0]), .rdup_out(a10_wr[516]), .rdlo_out(a10_wr[518]));
			radix2 #(.width(width)) rd_st9_517  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[517]), .rdlo_in(a9_wr[519]),  .coef_in(coef[512]), .rdup_out(a10_wr[517]), .rdlo_out(a10_wr[519]));
			radix2 #(.width(width)) rd_st9_520  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[520]), .rdlo_in(a9_wr[522]),  .coef_in(coef[0]), .rdup_out(a10_wr[520]), .rdlo_out(a10_wr[522]));
			radix2 #(.width(width)) rd_st9_521  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[521]), .rdlo_in(a9_wr[523]),  .coef_in(coef[512]), .rdup_out(a10_wr[521]), .rdlo_out(a10_wr[523]));
			radix2 #(.width(width)) rd_st9_524  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[524]), .rdlo_in(a9_wr[526]),  .coef_in(coef[0]), .rdup_out(a10_wr[524]), .rdlo_out(a10_wr[526]));
			radix2 #(.width(width)) rd_st9_525  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[525]), .rdlo_in(a9_wr[527]),  .coef_in(coef[512]), .rdup_out(a10_wr[525]), .rdlo_out(a10_wr[527]));
			radix2 #(.width(width)) rd_st9_528  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[528]), .rdlo_in(a9_wr[530]),  .coef_in(coef[0]), .rdup_out(a10_wr[528]), .rdlo_out(a10_wr[530]));
			radix2 #(.width(width)) rd_st9_529  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[529]), .rdlo_in(a9_wr[531]),  .coef_in(coef[512]), .rdup_out(a10_wr[529]), .rdlo_out(a10_wr[531]));
			radix2 #(.width(width)) rd_st9_532  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[532]), .rdlo_in(a9_wr[534]),  .coef_in(coef[0]), .rdup_out(a10_wr[532]), .rdlo_out(a10_wr[534]));
			radix2 #(.width(width)) rd_st9_533  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[533]), .rdlo_in(a9_wr[535]),  .coef_in(coef[512]), .rdup_out(a10_wr[533]), .rdlo_out(a10_wr[535]));
			radix2 #(.width(width)) rd_st9_536  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[536]), .rdlo_in(a9_wr[538]),  .coef_in(coef[0]), .rdup_out(a10_wr[536]), .rdlo_out(a10_wr[538]));
			radix2 #(.width(width)) rd_st9_537  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[537]), .rdlo_in(a9_wr[539]),  .coef_in(coef[512]), .rdup_out(a10_wr[537]), .rdlo_out(a10_wr[539]));
			radix2 #(.width(width)) rd_st9_540  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[540]), .rdlo_in(a9_wr[542]),  .coef_in(coef[0]), .rdup_out(a10_wr[540]), .rdlo_out(a10_wr[542]));
			radix2 #(.width(width)) rd_st9_541  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[541]), .rdlo_in(a9_wr[543]),  .coef_in(coef[512]), .rdup_out(a10_wr[541]), .rdlo_out(a10_wr[543]));
			radix2 #(.width(width)) rd_st9_544  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[544]), .rdlo_in(a9_wr[546]),  .coef_in(coef[0]), .rdup_out(a10_wr[544]), .rdlo_out(a10_wr[546]));
			radix2 #(.width(width)) rd_st9_545  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[545]), .rdlo_in(a9_wr[547]),  .coef_in(coef[512]), .rdup_out(a10_wr[545]), .rdlo_out(a10_wr[547]));
			radix2 #(.width(width)) rd_st9_548  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[548]), .rdlo_in(a9_wr[550]),  .coef_in(coef[0]), .rdup_out(a10_wr[548]), .rdlo_out(a10_wr[550]));
			radix2 #(.width(width)) rd_st9_549  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[549]), .rdlo_in(a9_wr[551]),  .coef_in(coef[512]), .rdup_out(a10_wr[549]), .rdlo_out(a10_wr[551]));
			radix2 #(.width(width)) rd_st9_552  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[552]), .rdlo_in(a9_wr[554]),  .coef_in(coef[0]), .rdup_out(a10_wr[552]), .rdlo_out(a10_wr[554]));
			radix2 #(.width(width)) rd_st9_553  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[553]), .rdlo_in(a9_wr[555]),  .coef_in(coef[512]), .rdup_out(a10_wr[553]), .rdlo_out(a10_wr[555]));
			radix2 #(.width(width)) rd_st9_556  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[556]), .rdlo_in(a9_wr[558]),  .coef_in(coef[0]), .rdup_out(a10_wr[556]), .rdlo_out(a10_wr[558]));
			radix2 #(.width(width)) rd_st9_557  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[557]), .rdlo_in(a9_wr[559]),  .coef_in(coef[512]), .rdup_out(a10_wr[557]), .rdlo_out(a10_wr[559]));
			radix2 #(.width(width)) rd_st9_560  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[560]), .rdlo_in(a9_wr[562]),  .coef_in(coef[0]), .rdup_out(a10_wr[560]), .rdlo_out(a10_wr[562]));
			radix2 #(.width(width)) rd_st9_561  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[561]), .rdlo_in(a9_wr[563]),  .coef_in(coef[512]), .rdup_out(a10_wr[561]), .rdlo_out(a10_wr[563]));
			radix2 #(.width(width)) rd_st9_564  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[564]), .rdlo_in(a9_wr[566]),  .coef_in(coef[0]), .rdup_out(a10_wr[564]), .rdlo_out(a10_wr[566]));
			radix2 #(.width(width)) rd_st9_565  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[565]), .rdlo_in(a9_wr[567]),  .coef_in(coef[512]), .rdup_out(a10_wr[565]), .rdlo_out(a10_wr[567]));
			radix2 #(.width(width)) rd_st9_568  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[568]), .rdlo_in(a9_wr[570]),  .coef_in(coef[0]), .rdup_out(a10_wr[568]), .rdlo_out(a10_wr[570]));
			radix2 #(.width(width)) rd_st9_569  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[569]), .rdlo_in(a9_wr[571]),  .coef_in(coef[512]), .rdup_out(a10_wr[569]), .rdlo_out(a10_wr[571]));
			radix2 #(.width(width)) rd_st9_572  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[572]), .rdlo_in(a9_wr[574]),  .coef_in(coef[0]), .rdup_out(a10_wr[572]), .rdlo_out(a10_wr[574]));
			radix2 #(.width(width)) rd_st9_573  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[573]), .rdlo_in(a9_wr[575]),  .coef_in(coef[512]), .rdup_out(a10_wr[573]), .rdlo_out(a10_wr[575]));
			radix2 #(.width(width)) rd_st9_576  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[576]), .rdlo_in(a9_wr[578]),  .coef_in(coef[0]), .rdup_out(a10_wr[576]), .rdlo_out(a10_wr[578]));
			radix2 #(.width(width)) rd_st9_577  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[577]), .rdlo_in(a9_wr[579]),  .coef_in(coef[512]), .rdup_out(a10_wr[577]), .rdlo_out(a10_wr[579]));
			radix2 #(.width(width)) rd_st9_580  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[580]), .rdlo_in(a9_wr[582]),  .coef_in(coef[0]), .rdup_out(a10_wr[580]), .rdlo_out(a10_wr[582]));
			radix2 #(.width(width)) rd_st9_581  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[581]), .rdlo_in(a9_wr[583]),  .coef_in(coef[512]), .rdup_out(a10_wr[581]), .rdlo_out(a10_wr[583]));
			radix2 #(.width(width)) rd_st9_584  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[584]), .rdlo_in(a9_wr[586]),  .coef_in(coef[0]), .rdup_out(a10_wr[584]), .rdlo_out(a10_wr[586]));
			radix2 #(.width(width)) rd_st9_585  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[585]), .rdlo_in(a9_wr[587]),  .coef_in(coef[512]), .rdup_out(a10_wr[585]), .rdlo_out(a10_wr[587]));
			radix2 #(.width(width)) rd_st9_588  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[588]), .rdlo_in(a9_wr[590]),  .coef_in(coef[0]), .rdup_out(a10_wr[588]), .rdlo_out(a10_wr[590]));
			radix2 #(.width(width)) rd_st9_589  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[589]), .rdlo_in(a9_wr[591]),  .coef_in(coef[512]), .rdup_out(a10_wr[589]), .rdlo_out(a10_wr[591]));
			radix2 #(.width(width)) rd_st9_592  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[592]), .rdlo_in(a9_wr[594]),  .coef_in(coef[0]), .rdup_out(a10_wr[592]), .rdlo_out(a10_wr[594]));
			radix2 #(.width(width)) rd_st9_593  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[593]), .rdlo_in(a9_wr[595]),  .coef_in(coef[512]), .rdup_out(a10_wr[593]), .rdlo_out(a10_wr[595]));
			radix2 #(.width(width)) rd_st9_596  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[596]), .rdlo_in(a9_wr[598]),  .coef_in(coef[0]), .rdup_out(a10_wr[596]), .rdlo_out(a10_wr[598]));
			radix2 #(.width(width)) rd_st9_597  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[597]), .rdlo_in(a9_wr[599]),  .coef_in(coef[512]), .rdup_out(a10_wr[597]), .rdlo_out(a10_wr[599]));
			radix2 #(.width(width)) rd_st9_600  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[600]), .rdlo_in(a9_wr[602]),  .coef_in(coef[0]), .rdup_out(a10_wr[600]), .rdlo_out(a10_wr[602]));
			radix2 #(.width(width)) rd_st9_601  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[601]), .rdlo_in(a9_wr[603]),  .coef_in(coef[512]), .rdup_out(a10_wr[601]), .rdlo_out(a10_wr[603]));
			radix2 #(.width(width)) rd_st9_604  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[604]), .rdlo_in(a9_wr[606]),  .coef_in(coef[0]), .rdup_out(a10_wr[604]), .rdlo_out(a10_wr[606]));
			radix2 #(.width(width)) rd_st9_605  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[605]), .rdlo_in(a9_wr[607]),  .coef_in(coef[512]), .rdup_out(a10_wr[605]), .rdlo_out(a10_wr[607]));
			radix2 #(.width(width)) rd_st9_608  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[608]), .rdlo_in(a9_wr[610]),  .coef_in(coef[0]), .rdup_out(a10_wr[608]), .rdlo_out(a10_wr[610]));
			radix2 #(.width(width)) rd_st9_609  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[609]), .rdlo_in(a9_wr[611]),  .coef_in(coef[512]), .rdup_out(a10_wr[609]), .rdlo_out(a10_wr[611]));
			radix2 #(.width(width)) rd_st9_612  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[612]), .rdlo_in(a9_wr[614]),  .coef_in(coef[0]), .rdup_out(a10_wr[612]), .rdlo_out(a10_wr[614]));
			radix2 #(.width(width)) rd_st9_613  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[613]), .rdlo_in(a9_wr[615]),  .coef_in(coef[512]), .rdup_out(a10_wr[613]), .rdlo_out(a10_wr[615]));
			radix2 #(.width(width)) rd_st9_616  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[616]), .rdlo_in(a9_wr[618]),  .coef_in(coef[0]), .rdup_out(a10_wr[616]), .rdlo_out(a10_wr[618]));
			radix2 #(.width(width)) rd_st9_617  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[617]), .rdlo_in(a9_wr[619]),  .coef_in(coef[512]), .rdup_out(a10_wr[617]), .rdlo_out(a10_wr[619]));
			radix2 #(.width(width)) rd_st9_620  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[620]), .rdlo_in(a9_wr[622]),  .coef_in(coef[0]), .rdup_out(a10_wr[620]), .rdlo_out(a10_wr[622]));
			radix2 #(.width(width)) rd_st9_621  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[621]), .rdlo_in(a9_wr[623]),  .coef_in(coef[512]), .rdup_out(a10_wr[621]), .rdlo_out(a10_wr[623]));
			radix2 #(.width(width)) rd_st9_624  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[624]), .rdlo_in(a9_wr[626]),  .coef_in(coef[0]), .rdup_out(a10_wr[624]), .rdlo_out(a10_wr[626]));
			radix2 #(.width(width)) rd_st9_625  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[625]), .rdlo_in(a9_wr[627]),  .coef_in(coef[512]), .rdup_out(a10_wr[625]), .rdlo_out(a10_wr[627]));
			radix2 #(.width(width)) rd_st9_628  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[628]), .rdlo_in(a9_wr[630]),  .coef_in(coef[0]), .rdup_out(a10_wr[628]), .rdlo_out(a10_wr[630]));
			radix2 #(.width(width)) rd_st9_629  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[629]), .rdlo_in(a9_wr[631]),  .coef_in(coef[512]), .rdup_out(a10_wr[629]), .rdlo_out(a10_wr[631]));
			radix2 #(.width(width)) rd_st9_632  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[632]), .rdlo_in(a9_wr[634]),  .coef_in(coef[0]), .rdup_out(a10_wr[632]), .rdlo_out(a10_wr[634]));
			radix2 #(.width(width)) rd_st9_633  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[633]), .rdlo_in(a9_wr[635]),  .coef_in(coef[512]), .rdup_out(a10_wr[633]), .rdlo_out(a10_wr[635]));
			radix2 #(.width(width)) rd_st9_636  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[636]), .rdlo_in(a9_wr[638]),  .coef_in(coef[0]), .rdup_out(a10_wr[636]), .rdlo_out(a10_wr[638]));
			radix2 #(.width(width)) rd_st9_637  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[637]), .rdlo_in(a9_wr[639]),  .coef_in(coef[512]), .rdup_out(a10_wr[637]), .rdlo_out(a10_wr[639]));
			radix2 #(.width(width)) rd_st9_640  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[640]), .rdlo_in(a9_wr[642]),  .coef_in(coef[0]), .rdup_out(a10_wr[640]), .rdlo_out(a10_wr[642]));
			radix2 #(.width(width)) rd_st9_641  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[641]), .rdlo_in(a9_wr[643]),  .coef_in(coef[512]), .rdup_out(a10_wr[641]), .rdlo_out(a10_wr[643]));
			radix2 #(.width(width)) rd_st9_644  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[644]), .rdlo_in(a9_wr[646]),  .coef_in(coef[0]), .rdup_out(a10_wr[644]), .rdlo_out(a10_wr[646]));
			radix2 #(.width(width)) rd_st9_645  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[645]), .rdlo_in(a9_wr[647]),  .coef_in(coef[512]), .rdup_out(a10_wr[645]), .rdlo_out(a10_wr[647]));
			radix2 #(.width(width)) rd_st9_648  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[648]), .rdlo_in(a9_wr[650]),  .coef_in(coef[0]), .rdup_out(a10_wr[648]), .rdlo_out(a10_wr[650]));
			radix2 #(.width(width)) rd_st9_649  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[649]), .rdlo_in(a9_wr[651]),  .coef_in(coef[512]), .rdup_out(a10_wr[649]), .rdlo_out(a10_wr[651]));
			radix2 #(.width(width)) rd_st9_652  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[652]), .rdlo_in(a9_wr[654]),  .coef_in(coef[0]), .rdup_out(a10_wr[652]), .rdlo_out(a10_wr[654]));
			radix2 #(.width(width)) rd_st9_653  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[653]), .rdlo_in(a9_wr[655]),  .coef_in(coef[512]), .rdup_out(a10_wr[653]), .rdlo_out(a10_wr[655]));
			radix2 #(.width(width)) rd_st9_656  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[656]), .rdlo_in(a9_wr[658]),  .coef_in(coef[0]), .rdup_out(a10_wr[656]), .rdlo_out(a10_wr[658]));
			radix2 #(.width(width)) rd_st9_657  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[657]), .rdlo_in(a9_wr[659]),  .coef_in(coef[512]), .rdup_out(a10_wr[657]), .rdlo_out(a10_wr[659]));
			radix2 #(.width(width)) rd_st9_660  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[660]), .rdlo_in(a9_wr[662]),  .coef_in(coef[0]), .rdup_out(a10_wr[660]), .rdlo_out(a10_wr[662]));
			radix2 #(.width(width)) rd_st9_661  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[661]), .rdlo_in(a9_wr[663]),  .coef_in(coef[512]), .rdup_out(a10_wr[661]), .rdlo_out(a10_wr[663]));
			radix2 #(.width(width)) rd_st9_664  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[664]), .rdlo_in(a9_wr[666]),  .coef_in(coef[0]), .rdup_out(a10_wr[664]), .rdlo_out(a10_wr[666]));
			radix2 #(.width(width)) rd_st9_665  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[665]), .rdlo_in(a9_wr[667]),  .coef_in(coef[512]), .rdup_out(a10_wr[665]), .rdlo_out(a10_wr[667]));
			radix2 #(.width(width)) rd_st9_668  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[668]), .rdlo_in(a9_wr[670]),  .coef_in(coef[0]), .rdup_out(a10_wr[668]), .rdlo_out(a10_wr[670]));
			radix2 #(.width(width)) rd_st9_669  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[669]), .rdlo_in(a9_wr[671]),  .coef_in(coef[512]), .rdup_out(a10_wr[669]), .rdlo_out(a10_wr[671]));
			radix2 #(.width(width)) rd_st9_672  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[672]), .rdlo_in(a9_wr[674]),  .coef_in(coef[0]), .rdup_out(a10_wr[672]), .rdlo_out(a10_wr[674]));
			radix2 #(.width(width)) rd_st9_673  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[673]), .rdlo_in(a9_wr[675]),  .coef_in(coef[512]), .rdup_out(a10_wr[673]), .rdlo_out(a10_wr[675]));
			radix2 #(.width(width)) rd_st9_676  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[676]), .rdlo_in(a9_wr[678]),  .coef_in(coef[0]), .rdup_out(a10_wr[676]), .rdlo_out(a10_wr[678]));
			radix2 #(.width(width)) rd_st9_677  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[677]), .rdlo_in(a9_wr[679]),  .coef_in(coef[512]), .rdup_out(a10_wr[677]), .rdlo_out(a10_wr[679]));
			radix2 #(.width(width)) rd_st9_680  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[680]), .rdlo_in(a9_wr[682]),  .coef_in(coef[0]), .rdup_out(a10_wr[680]), .rdlo_out(a10_wr[682]));
			radix2 #(.width(width)) rd_st9_681  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[681]), .rdlo_in(a9_wr[683]),  .coef_in(coef[512]), .rdup_out(a10_wr[681]), .rdlo_out(a10_wr[683]));
			radix2 #(.width(width)) rd_st9_684  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[684]), .rdlo_in(a9_wr[686]),  .coef_in(coef[0]), .rdup_out(a10_wr[684]), .rdlo_out(a10_wr[686]));
			radix2 #(.width(width)) rd_st9_685  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[685]), .rdlo_in(a9_wr[687]),  .coef_in(coef[512]), .rdup_out(a10_wr[685]), .rdlo_out(a10_wr[687]));
			radix2 #(.width(width)) rd_st9_688  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[688]), .rdlo_in(a9_wr[690]),  .coef_in(coef[0]), .rdup_out(a10_wr[688]), .rdlo_out(a10_wr[690]));
			radix2 #(.width(width)) rd_st9_689  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[689]), .rdlo_in(a9_wr[691]),  .coef_in(coef[512]), .rdup_out(a10_wr[689]), .rdlo_out(a10_wr[691]));
			radix2 #(.width(width)) rd_st9_692  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[692]), .rdlo_in(a9_wr[694]),  .coef_in(coef[0]), .rdup_out(a10_wr[692]), .rdlo_out(a10_wr[694]));
			radix2 #(.width(width)) rd_st9_693  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[693]), .rdlo_in(a9_wr[695]),  .coef_in(coef[512]), .rdup_out(a10_wr[693]), .rdlo_out(a10_wr[695]));
			radix2 #(.width(width)) rd_st9_696  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[696]), .rdlo_in(a9_wr[698]),  .coef_in(coef[0]), .rdup_out(a10_wr[696]), .rdlo_out(a10_wr[698]));
			radix2 #(.width(width)) rd_st9_697  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[697]), .rdlo_in(a9_wr[699]),  .coef_in(coef[512]), .rdup_out(a10_wr[697]), .rdlo_out(a10_wr[699]));
			radix2 #(.width(width)) rd_st9_700  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[700]), .rdlo_in(a9_wr[702]),  .coef_in(coef[0]), .rdup_out(a10_wr[700]), .rdlo_out(a10_wr[702]));
			radix2 #(.width(width)) rd_st9_701  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[701]), .rdlo_in(a9_wr[703]),  .coef_in(coef[512]), .rdup_out(a10_wr[701]), .rdlo_out(a10_wr[703]));
			radix2 #(.width(width)) rd_st9_704  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[704]), .rdlo_in(a9_wr[706]),  .coef_in(coef[0]), .rdup_out(a10_wr[704]), .rdlo_out(a10_wr[706]));
			radix2 #(.width(width)) rd_st9_705  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[705]), .rdlo_in(a9_wr[707]),  .coef_in(coef[512]), .rdup_out(a10_wr[705]), .rdlo_out(a10_wr[707]));
			radix2 #(.width(width)) rd_st9_708  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[708]), .rdlo_in(a9_wr[710]),  .coef_in(coef[0]), .rdup_out(a10_wr[708]), .rdlo_out(a10_wr[710]));
			radix2 #(.width(width)) rd_st9_709  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[709]), .rdlo_in(a9_wr[711]),  .coef_in(coef[512]), .rdup_out(a10_wr[709]), .rdlo_out(a10_wr[711]));
			radix2 #(.width(width)) rd_st9_712  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[712]), .rdlo_in(a9_wr[714]),  .coef_in(coef[0]), .rdup_out(a10_wr[712]), .rdlo_out(a10_wr[714]));
			radix2 #(.width(width)) rd_st9_713  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[713]), .rdlo_in(a9_wr[715]),  .coef_in(coef[512]), .rdup_out(a10_wr[713]), .rdlo_out(a10_wr[715]));
			radix2 #(.width(width)) rd_st9_716  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[716]), .rdlo_in(a9_wr[718]),  .coef_in(coef[0]), .rdup_out(a10_wr[716]), .rdlo_out(a10_wr[718]));
			radix2 #(.width(width)) rd_st9_717  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[717]), .rdlo_in(a9_wr[719]),  .coef_in(coef[512]), .rdup_out(a10_wr[717]), .rdlo_out(a10_wr[719]));
			radix2 #(.width(width)) rd_st9_720  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[720]), .rdlo_in(a9_wr[722]),  .coef_in(coef[0]), .rdup_out(a10_wr[720]), .rdlo_out(a10_wr[722]));
			radix2 #(.width(width)) rd_st9_721  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[721]), .rdlo_in(a9_wr[723]),  .coef_in(coef[512]), .rdup_out(a10_wr[721]), .rdlo_out(a10_wr[723]));
			radix2 #(.width(width)) rd_st9_724  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[724]), .rdlo_in(a9_wr[726]),  .coef_in(coef[0]), .rdup_out(a10_wr[724]), .rdlo_out(a10_wr[726]));
			radix2 #(.width(width)) rd_st9_725  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[725]), .rdlo_in(a9_wr[727]),  .coef_in(coef[512]), .rdup_out(a10_wr[725]), .rdlo_out(a10_wr[727]));
			radix2 #(.width(width)) rd_st9_728  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[728]), .rdlo_in(a9_wr[730]),  .coef_in(coef[0]), .rdup_out(a10_wr[728]), .rdlo_out(a10_wr[730]));
			radix2 #(.width(width)) rd_st9_729  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[729]), .rdlo_in(a9_wr[731]),  .coef_in(coef[512]), .rdup_out(a10_wr[729]), .rdlo_out(a10_wr[731]));
			radix2 #(.width(width)) rd_st9_732  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[732]), .rdlo_in(a9_wr[734]),  .coef_in(coef[0]), .rdup_out(a10_wr[732]), .rdlo_out(a10_wr[734]));
			radix2 #(.width(width)) rd_st9_733  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[733]), .rdlo_in(a9_wr[735]),  .coef_in(coef[512]), .rdup_out(a10_wr[733]), .rdlo_out(a10_wr[735]));
			radix2 #(.width(width)) rd_st9_736  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[736]), .rdlo_in(a9_wr[738]),  .coef_in(coef[0]), .rdup_out(a10_wr[736]), .rdlo_out(a10_wr[738]));
			radix2 #(.width(width)) rd_st9_737  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[737]), .rdlo_in(a9_wr[739]),  .coef_in(coef[512]), .rdup_out(a10_wr[737]), .rdlo_out(a10_wr[739]));
			radix2 #(.width(width)) rd_st9_740  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[740]), .rdlo_in(a9_wr[742]),  .coef_in(coef[0]), .rdup_out(a10_wr[740]), .rdlo_out(a10_wr[742]));
			radix2 #(.width(width)) rd_st9_741  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[741]), .rdlo_in(a9_wr[743]),  .coef_in(coef[512]), .rdup_out(a10_wr[741]), .rdlo_out(a10_wr[743]));
			radix2 #(.width(width)) rd_st9_744  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[744]), .rdlo_in(a9_wr[746]),  .coef_in(coef[0]), .rdup_out(a10_wr[744]), .rdlo_out(a10_wr[746]));
			radix2 #(.width(width)) rd_st9_745  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[745]), .rdlo_in(a9_wr[747]),  .coef_in(coef[512]), .rdup_out(a10_wr[745]), .rdlo_out(a10_wr[747]));
			radix2 #(.width(width)) rd_st9_748  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[748]), .rdlo_in(a9_wr[750]),  .coef_in(coef[0]), .rdup_out(a10_wr[748]), .rdlo_out(a10_wr[750]));
			radix2 #(.width(width)) rd_st9_749  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[749]), .rdlo_in(a9_wr[751]),  .coef_in(coef[512]), .rdup_out(a10_wr[749]), .rdlo_out(a10_wr[751]));
			radix2 #(.width(width)) rd_st9_752  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[752]), .rdlo_in(a9_wr[754]),  .coef_in(coef[0]), .rdup_out(a10_wr[752]), .rdlo_out(a10_wr[754]));
			radix2 #(.width(width)) rd_st9_753  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[753]), .rdlo_in(a9_wr[755]),  .coef_in(coef[512]), .rdup_out(a10_wr[753]), .rdlo_out(a10_wr[755]));
			radix2 #(.width(width)) rd_st9_756  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[756]), .rdlo_in(a9_wr[758]),  .coef_in(coef[0]), .rdup_out(a10_wr[756]), .rdlo_out(a10_wr[758]));
			radix2 #(.width(width)) rd_st9_757  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[757]), .rdlo_in(a9_wr[759]),  .coef_in(coef[512]), .rdup_out(a10_wr[757]), .rdlo_out(a10_wr[759]));
			radix2 #(.width(width)) rd_st9_760  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[760]), .rdlo_in(a9_wr[762]),  .coef_in(coef[0]), .rdup_out(a10_wr[760]), .rdlo_out(a10_wr[762]));
			radix2 #(.width(width)) rd_st9_761  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[761]), .rdlo_in(a9_wr[763]),  .coef_in(coef[512]), .rdup_out(a10_wr[761]), .rdlo_out(a10_wr[763]));
			radix2 #(.width(width)) rd_st9_764  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[764]), .rdlo_in(a9_wr[766]),  .coef_in(coef[0]), .rdup_out(a10_wr[764]), .rdlo_out(a10_wr[766]));
			radix2 #(.width(width)) rd_st9_765  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[765]), .rdlo_in(a9_wr[767]),  .coef_in(coef[512]), .rdup_out(a10_wr[765]), .rdlo_out(a10_wr[767]));
			radix2 #(.width(width)) rd_st9_768  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[768]), .rdlo_in(a9_wr[770]),  .coef_in(coef[0]), .rdup_out(a10_wr[768]), .rdlo_out(a10_wr[770]));
			radix2 #(.width(width)) rd_st9_769  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[769]), .rdlo_in(a9_wr[771]),  .coef_in(coef[512]), .rdup_out(a10_wr[769]), .rdlo_out(a10_wr[771]));
			radix2 #(.width(width)) rd_st9_772  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[772]), .rdlo_in(a9_wr[774]),  .coef_in(coef[0]), .rdup_out(a10_wr[772]), .rdlo_out(a10_wr[774]));
			radix2 #(.width(width)) rd_st9_773  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[773]), .rdlo_in(a9_wr[775]),  .coef_in(coef[512]), .rdup_out(a10_wr[773]), .rdlo_out(a10_wr[775]));
			radix2 #(.width(width)) rd_st9_776  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[776]), .rdlo_in(a9_wr[778]),  .coef_in(coef[0]), .rdup_out(a10_wr[776]), .rdlo_out(a10_wr[778]));
			radix2 #(.width(width)) rd_st9_777  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[777]), .rdlo_in(a9_wr[779]),  .coef_in(coef[512]), .rdup_out(a10_wr[777]), .rdlo_out(a10_wr[779]));
			radix2 #(.width(width)) rd_st9_780  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[780]), .rdlo_in(a9_wr[782]),  .coef_in(coef[0]), .rdup_out(a10_wr[780]), .rdlo_out(a10_wr[782]));
			radix2 #(.width(width)) rd_st9_781  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[781]), .rdlo_in(a9_wr[783]),  .coef_in(coef[512]), .rdup_out(a10_wr[781]), .rdlo_out(a10_wr[783]));
			radix2 #(.width(width)) rd_st9_784  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[784]), .rdlo_in(a9_wr[786]),  .coef_in(coef[0]), .rdup_out(a10_wr[784]), .rdlo_out(a10_wr[786]));
			radix2 #(.width(width)) rd_st9_785  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[785]), .rdlo_in(a9_wr[787]),  .coef_in(coef[512]), .rdup_out(a10_wr[785]), .rdlo_out(a10_wr[787]));
			radix2 #(.width(width)) rd_st9_788  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[788]), .rdlo_in(a9_wr[790]),  .coef_in(coef[0]), .rdup_out(a10_wr[788]), .rdlo_out(a10_wr[790]));
			radix2 #(.width(width)) rd_st9_789  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[789]), .rdlo_in(a9_wr[791]),  .coef_in(coef[512]), .rdup_out(a10_wr[789]), .rdlo_out(a10_wr[791]));
			radix2 #(.width(width)) rd_st9_792  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[792]), .rdlo_in(a9_wr[794]),  .coef_in(coef[0]), .rdup_out(a10_wr[792]), .rdlo_out(a10_wr[794]));
			radix2 #(.width(width)) rd_st9_793  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[793]), .rdlo_in(a9_wr[795]),  .coef_in(coef[512]), .rdup_out(a10_wr[793]), .rdlo_out(a10_wr[795]));
			radix2 #(.width(width)) rd_st9_796  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[796]), .rdlo_in(a9_wr[798]),  .coef_in(coef[0]), .rdup_out(a10_wr[796]), .rdlo_out(a10_wr[798]));
			radix2 #(.width(width)) rd_st9_797  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[797]), .rdlo_in(a9_wr[799]),  .coef_in(coef[512]), .rdup_out(a10_wr[797]), .rdlo_out(a10_wr[799]));
			radix2 #(.width(width)) rd_st9_800  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[800]), .rdlo_in(a9_wr[802]),  .coef_in(coef[0]), .rdup_out(a10_wr[800]), .rdlo_out(a10_wr[802]));
			radix2 #(.width(width)) rd_st9_801  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[801]), .rdlo_in(a9_wr[803]),  .coef_in(coef[512]), .rdup_out(a10_wr[801]), .rdlo_out(a10_wr[803]));
			radix2 #(.width(width)) rd_st9_804  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[804]), .rdlo_in(a9_wr[806]),  .coef_in(coef[0]), .rdup_out(a10_wr[804]), .rdlo_out(a10_wr[806]));
			radix2 #(.width(width)) rd_st9_805  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[805]), .rdlo_in(a9_wr[807]),  .coef_in(coef[512]), .rdup_out(a10_wr[805]), .rdlo_out(a10_wr[807]));
			radix2 #(.width(width)) rd_st9_808  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[808]), .rdlo_in(a9_wr[810]),  .coef_in(coef[0]), .rdup_out(a10_wr[808]), .rdlo_out(a10_wr[810]));
			radix2 #(.width(width)) rd_st9_809  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[809]), .rdlo_in(a9_wr[811]),  .coef_in(coef[512]), .rdup_out(a10_wr[809]), .rdlo_out(a10_wr[811]));
			radix2 #(.width(width)) rd_st9_812  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[812]), .rdlo_in(a9_wr[814]),  .coef_in(coef[0]), .rdup_out(a10_wr[812]), .rdlo_out(a10_wr[814]));
			radix2 #(.width(width)) rd_st9_813  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[813]), .rdlo_in(a9_wr[815]),  .coef_in(coef[512]), .rdup_out(a10_wr[813]), .rdlo_out(a10_wr[815]));
			radix2 #(.width(width)) rd_st9_816  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[816]), .rdlo_in(a9_wr[818]),  .coef_in(coef[0]), .rdup_out(a10_wr[816]), .rdlo_out(a10_wr[818]));
			radix2 #(.width(width)) rd_st9_817  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[817]), .rdlo_in(a9_wr[819]),  .coef_in(coef[512]), .rdup_out(a10_wr[817]), .rdlo_out(a10_wr[819]));
			radix2 #(.width(width)) rd_st9_820  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[820]), .rdlo_in(a9_wr[822]),  .coef_in(coef[0]), .rdup_out(a10_wr[820]), .rdlo_out(a10_wr[822]));
			radix2 #(.width(width)) rd_st9_821  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[821]), .rdlo_in(a9_wr[823]),  .coef_in(coef[512]), .rdup_out(a10_wr[821]), .rdlo_out(a10_wr[823]));
			radix2 #(.width(width)) rd_st9_824  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[824]), .rdlo_in(a9_wr[826]),  .coef_in(coef[0]), .rdup_out(a10_wr[824]), .rdlo_out(a10_wr[826]));
			radix2 #(.width(width)) rd_st9_825  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[825]), .rdlo_in(a9_wr[827]),  .coef_in(coef[512]), .rdup_out(a10_wr[825]), .rdlo_out(a10_wr[827]));
			radix2 #(.width(width)) rd_st9_828  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[828]), .rdlo_in(a9_wr[830]),  .coef_in(coef[0]), .rdup_out(a10_wr[828]), .rdlo_out(a10_wr[830]));
			radix2 #(.width(width)) rd_st9_829  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[829]), .rdlo_in(a9_wr[831]),  .coef_in(coef[512]), .rdup_out(a10_wr[829]), .rdlo_out(a10_wr[831]));
			radix2 #(.width(width)) rd_st9_832  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[832]), .rdlo_in(a9_wr[834]),  .coef_in(coef[0]), .rdup_out(a10_wr[832]), .rdlo_out(a10_wr[834]));
			radix2 #(.width(width)) rd_st9_833  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[833]), .rdlo_in(a9_wr[835]),  .coef_in(coef[512]), .rdup_out(a10_wr[833]), .rdlo_out(a10_wr[835]));
			radix2 #(.width(width)) rd_st9_836  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[836]), .rdlo_in(a9_wr[838]),  .coef_in(coef[0]), .rdup_out(a10_wr[836]), .rdlo_out(a10_wr[838]));
			radix2 #(.width(width)) rd_st9_837  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[837]), .rdlo_in(a9_wr[839]),  .coef_in(coef[512]), .rdup_out(a10_wr[837]), .rdlo_out(a10_wr[839]));
			radix2 #(.width(width)) rd_st9_840  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[840]), .rdlo_in(a9_wr[842]),  .coef_in(coef[0]), .rdup_out(a10_wr[840]), .rdlo_out(a10_wr[842]));
			radix2 #(.width(width)) rd_st9_841  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[841]), .rdlo_in(a9_wr[843]),  .coef_in(coef[512]), .rdup_out(a10_wr[841]), .rdlo_out(a10_wr[843]));
			radix2 #(.width(width)) rd_st9_844  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[844]), .rdlo_in(a9_wr[846]),  .coef_in(coef[0]), .rdup_out(a10_wr[844]), .rdlo_out(a10_wr[846]));
			radix2 #(.width(width)) rd_st9_845  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[845]), .rdlo_in(a9_wr[847]),  .coef_in(coef[512]), .rdup_out(a10_wr[845]), .rdlo_out(a10_wr[847]));
			radix2 #(.width(width)) rd_st9_848  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[848]), .rdlo_in(a9_wr[850]),  .coef_in(coef[0]), .rdup_out(a10_wr[848]), .rdlo_out(a10_wr[850]));
			radix2 #(.width(width)) rd_st9_849  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[849]), .rdlo_in(a9_wr[851]),  .coef_in(coef[512]), .rdup_out(a10_wr[849]), .rdlo_out(a10_wr[851]));
			radix2 #(.width(width)) rd_st9_852  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[852]), .rdlo_in(a9_wr[854]),  .coef_in(coef[0]), .rdup_out(a10_wr[852]), .rdlo_out(a10_wr[854]));
			radix2 #(.width(width)) rd_st9_853  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[853]), .rdlo_in(a9_wr[855]),  .coef_in(coef[512]), .rdup_out(a10_wr[853]), .rdlo_out(a10_wr[855]));
			radix2 #(.width(width)) rd_st9_856  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[856]), .rdlo_in(a9_wr[858]),  .coef_in(coef[0]), .rdup_out(a10_wr[856]), .rdlo_out(a10_wr[858]));
			radix2 #(.width(width)) rd_st9_857  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[857]), .rdlo_in(a9_wr[859]),  .coef_in(coef[512]), .rdup_out(a10_wr[857]), .rdlo_out(a10_wr[859]));
			radix2 #(.width(width)) rd_st9_860  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[860]), .rdlo_in(a9_wr[862]),  .coef_in(coef[0]), .rdup_out(a10_wr[860]), .rdlo_out(a10_wr[862]));
			radix2 #(.width(width)) rd_st9_861  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[861]), .rdlo_in(a9_wr[863]),  .coef_in(coef[512]), .rdup_out(a10_wr[861]), .rdlo_out(a10_wr[863]));
			radix2 #(.width(width)) rd_st9_864  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[864]), .rdlo_in(a9_wr[866]),  .coef_in(coef[0]), .rdup_out(a10_wr[864]), .rdlo_out(a10_wr[866]));
			radix2 #(.width(width)) rd_st9_865  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[865]), .rdlo_in(a9_wr[867]),  .coef_in(coef[512]), .rdup_out(a10_wr[865]), .rdlo_out(a10_wr[867]));
			radix2 #(.width(width)) rd_st9_868  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[868]), .rdlo_in(a9_wr[870]),  .coef_in(coef[0]), .rdup_out(a10_wr[868]), .rdlo_out(a10_wr[870]));
			radix2 #(.width(width)) rd_st9_869  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[869]), .rdlo_in(a9_wr[871]),  .coef_in(coef[512]), .rdup_out(a10_wr[869]), .rdlo_out(a10_wr[871]));
			radix2 #(.width(width)) rd_st9_872  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[872]), .rdlo_in(a9_wr[874]),  .coef_in(coef[0]), .rdup_out(a10_wr[872]), .rdlo_out(a10_wr[874]));
			radix2 #(.width(width)) rd_st9_873  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[873]), .rdlo_in(a9_wr[875]),  .coef_in(coef[512]), .rdup_out(a10_wr[873]), .rdlo_out(a10_wr[875]));
			radix2 #(.width(width)) rd_st9_876  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[876]), .rdlo_in(a9_wr[878]),  .coef_in(coef[0]), .rdup_out(a10_wr[876]), .rdlo_out(a10_wr[878]));
			radix2 #(.width(width)) rd_st9_877  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[877]), .rdlo_in(a9_wr[879]),  .coef_in(coef[512]), .rdup_out(a10_wr[877]), .rdlo_out(a10_wr[879]));
			radix2 #(.width(width)) rd_st9_880  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[880]), .rdlo_in(a9_wr[882]),  .coef_in(coef[0]), .rdup_out(a10_wr[880]), .rdlo_out(a10_wr[882]));
			radix2 #(.width(width)) rd_st9_881  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[881]), .rdlo_in(a9_wr[883]),  .coef_in(coef[512]), .rdup_out(a10_wr[881]), .rdlo_out(a10_wr[883]));
			radix2 #(.width(width)) rd_st9_884  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[884]), .rdlo_in(a9_wr[886]),  .coef_in(coef[0]), .rdup_out(a10_wr[884]), .rdlo_out(a10_wr[886]));
			radix2 #(.width(width)) rd_st9_885  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[885]), .rdlo_in(a9_wr[887]),  .coef_in(coef[512]), .rdup_out(a10_wr[885]), .rdlo_out(a10_wr[887]));
			radix2 #(.width(width)) rd_st9_888  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[888]), .rdlo_in(a9_wr[890]),  .coef_in(coef[0]), .rdup_out(a10_wr[888]), .rdlo_out(a10_wr[890]));
			radix2 #(.width(width)) rd_st9_889  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[889]), .rdlo_in(a9_wr[891]),  .coef_in(coef[512]), .rdup_out(a10_wr[889]), .rdlo_out(a10_wr[891]));
			radix2 #(.width(width)) rd_st9_892  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[892]), .rdlo_in(a9_wr[894]),  .coef_in(coef[0]), .rdup_out(a10_wr[892]), .rdlo_out(a10_wr[894]));
			radix2 #(.width(width)) rd_st9_893  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[893]), .rdlo_in(a9_wr[895]),  .coef_in(coef[512]), .rdup_out(a10_wr[893]), .rdlo_out(a10_wr[895]));
			radix2 #(.width(width)) rd_st9_896  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[896]), .rdlo_in(a9_wr[898]),  .coef_in(coef[0]), .rdup_out(a10_wr[896]), .rdlo_out(a10_wr[898]));
			radix2 #(.width(width)) rd_st9_897  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[897]), .rdlo_in(a9_wr[899]),  .coef_in(coef[512]), .rdup_out(a10_wr[897]), .rdlo_out(a10_wr[899]));
			radix2 #(.width(width)) rd_st9_900  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[900]), .rdlo_in(a9_wr[902]),  .coef_in(coef[0]), .rdup_out(a10_wr[900]), .rdlo_out(a10_wr[902]));
			radix2 #(.width(width)) rd_st9_901  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[901]), .rdlo_in(a9_wr[903]),  .coef_in(coef[512]), .rdup_out(a10_wr[901]), .rdlo_out(a10_wr[903]));
			radix2 #(.width(width)) rd_st9_904  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[904]), .rdlo_in(a9_wr[906]),  .coef_in(coef[0]), .rdup_out(a10_wr[904]), .rdlo_out(a10_wr[906]));
			radix2 #(.width(width)) rd_st9_905  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[905]), .rdlo_in(a9_wr[907]),  .coef_in(coef[512]), .rdup_out(a10_wr[905]), .rdlo_out(a10_wr[907]));
			radix2 #(.width(width)) rd_st9_908  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[908]), .rdlo_in(a9_wr[910]),  .coef_in(coef[0]), .rdup_out(a10_wr[908]), .rdlo_out(a10_wr[910]));
			radix2 #(.width(width)) rd_st9_909  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[909]), .rdlo_in(a9_wr[911]),  .coef_in(coef[512]), .rdup_out(a10_wr[909]), .rdlo_out(a10_wr[911]));
			radix2 #(.width(width)) rd_st9_912  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[912]), .rdlo_in(a9_wr[914]),  .coef_in(coef[0]), .rdup_out(a10_wr[912]), .rdlo_out(a10_wr[914]));
			radix2 #(.width(width)) rd_st9_913  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[913]), .rdlo_in(a9_wr[915]),  .coef_in(coef[512]), .rdup_out(a10_wr[913]), .rdlo_out(a10_wr[915]));
			radix2 #(.width(width)) rd_st9_916  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[916]), .rdlo_in(a9_wr[918]),  .coef_in(coef[0]), .rdup_out(a10_wr[916]), .rdlo_out(a10_wr[918]));
			radix2 #(.width(width)) rd_st9_917  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[917]), .rdlo_in(a9_wr[919]),  .coef_in(coef[512]), .rdup_out(a10_wr[917]), .rdlo_out(a10_wr[919]));
			radix2 #(.width(width)) rd_st9_920  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[920]), .rdlo_in(a9_wr[922]),  .coef_in(coef[0]), .rdup_out(a10_wr[920]), .rdlo_out(a10_wr[922]));
			radix2 #(.width(width)) rd_st9_921  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[921]), .rdlo_in(a9_wr[923]),  .coef_in(coef[512]), .rdup_out(a10_wr[921]), .rdlo_out(a10_wr[923]));
			radix2 #(.width(width)) rd_st9_924  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[924]), .rdlo_in(a9_wr[926]),  .coef_in(coef[0]), .rdup_out(a10_wr[924]), .rdlo_out(a10_wr[926]));
			radix2 #(.width(width)) rd_st9_925  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[925]), .rdlo_in(a9_wr[927]),  .coef_in(coef[512]), .rdup_out(a10_wr[925]), .rdlo_out(a10_wr[927]));
			radix2 #(.width(width)) rd_st9_928  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[928]), .rdlo_in(a9_wr[930]),  .coef_in(coef[0]), .rdup_out(a10_wr[928]), .rdlo_out(a10_wr[930]));
			radix2 #(.width(width)) rd_st9_929  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[929]), .rdlo_in(a9_wr[931]),  .coef_in(coef[512]), .rdup_out(a10_wr[929]), .rdlo_out(a10_wr[931]));
			radix2 #(.width(width)) rd_st9_932  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[932]), .rdlo_in(a9_wr[934]),  .coef_in(coef[0]), .rdup_out(a10_wr[932]), .rdlo_out(a10_wr[934]));
			radix2 #(.width(width)) rd_st9_933  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[933]), .rdlo_in(a9_wr[935]),  .coef_in(coef[512]), .rdup_out(a10_wr[933]), .rdlo_out(a10_wr[935]));
			radix2 #(.width(width)) rd_st9_936  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[936]), .rdlo_in(a9_wr[938]),  .coef_in(coef[0]), .rdup_out(a10_wr[936]), .rdlo_out(a10_wr[938]));
			radix2 #(.width(width)) rd_st9_937  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[937]), .rdlo_in(a9_wr[939]),  .coef_in(coef[512]), .rdup_out(a10_wr[937]), .rdlo_out(a10_wr[939]));
			radix2 #(.width(width)) rd_st9_940  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[940]), .rdlo_in(a9_wr[942]),  .coef_in(coef[0]), .rdup_out(a10_wr[940]), .rdlo_out(a10_wr[942]));
			radix2 #(.width(width)) rd_st9_941  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[941]), .rdlo_in(a9_wr[943]),  .coef_in(coef[512]), .rdup_out(a10_wr[941]), .rdlo_out(a10_wr[943]));
			radix2 #(.width(width)) rd_st9_944  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[944]), .rdlo_in(a9_wr[946]),  .coef_in(coef[0]), .rdup_out(a10_wr[944]), .rdlo_out(a10_wr[946]));
			radix2 #(.width(width)) rd_st9_945  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[945]), .rdlo_in(a9_wr[947]),  .coef_in(coef[512]), .rdup_out(a10_wr[945]), .rdlo_out(a10_wr[947]));
			radix2 #(.width(width)) rd_st9_948  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[948]), .rdlo_in(a9_wr[950]),  .coef_in(coef[0]), .rdup_out(a10_wr[948]), .rdlo_out(a10_wr[950]));
			radix2 #(.width(width)) rd_st9_949  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[949]), .rdlo_in(a9_wr[951]),  .coef_in(coef[512]), .rdup_out(a10_wr[949]), .rdlo_out(a10_wr[951]));
			radix2 #(.width(width)) rd_st9_952  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[952]), .rdlo_in(a9_wr[954]),  .coef_in(coef[0]), .rdup_out(a10_wr[952]), .rdlo_out(a10_wr[954]));
			radix2 #(.width(width)) rd_st9_953  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[953]), .rdlo_in(a9_wr[955]),  .coef_in(coef[512]), .rdup_out(a10_wr[953]), .rdlo_out(a10_wr[955]));
			radix2 #(.width(width)) rd_st9_956  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[956]), .rdlo_in(a9_wr[958]),  .coef_in(coef[0]), .rdup_out(a10_wr[956]), .rdlo_out(a10_wr[958]));
			radix2 #(.width(width)) rd_st9_957  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[957]), .rdlo_in(a9_wr[959]),  .coef_in(coef[512]), .rdup_out(a10_wr[957]), .rdlo_out(a10_wr[959]));
			radix2 #(.width(width)) rd_st9_960  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[960]), .rdlo_in(a9_wr[962]),  .coef_in(coef[0]), .rdup_out(a10_wr[960]), .rdlo_out(a10_wr[962]));
			radix2 #(.width(width)) rd_st9_961  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[961]), .rdlo_in(a9_wr[963]),  .coef_in(coef[512]), .rdup_out(a10_wr[961]), .rdlo_out(a10_wr[963]));
			radix2 #(.width(width)) rd_st9_964  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[964]), .rdlo_in(a9_wr[966]),  .coef_in(coef[0]), .rdup_out(a10_wr[964]), .rdlo_out(a10_wr[966]));
			radix2 #(.width(width)) rd_st9_965  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[965]), .rdlo_in(a9_wr[967]),  .coef_in(coef[512]), .rdup_out(a10_wr[965]), .rdlo_out(a10_wr[967]));
			radix2 #(.width(width)) rd_st9_968  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[968]), .rdlo_in(a9_wr[970]),  .coef_in(coef[0]), .rdup_out(a10_wr[968]), .rdlo_out(a10_wr[970]));
			radix2 #(.width(width)) rd_st9_969  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[969]), .rdlo_in(a9_wr[971]),  .coef_in(coef[512]), .rdup_out(a10_wr[969]), .rdlo_out(a10_wr[971]));
			radix2 #(.width(width)) rd_st9_972  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[972]), .rdlo_in(a9_wr[974]),  .coef_in(coef[0]), .rdup_out(a10_wr[972]), .rdlo_out(a10_wr[974]));
			radix2 #(.width(width)) rd_st9_973  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[973]), .rdlo_in(a9_wr[975]),  .coef_in(coef[512]), .rdup_out(a10_wr[973]), .rdlo_out(a10_wr[975]));
			radix2 #(.width(width)) rd_st9_976  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[976]), .rdlo_in(a9_wr[978]),  .coef_in(coef[0]), .rdup_out(a10_wr[976]), .rdlo_out(a10_wr[978]));
			radix2 #(.width(width)) rd_st9_977  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[977]), .rdlo_in(a9_wr[979]),  .coef_in(coef[512]), .rdup_out(a10_wr[977]), .rdlo_out(a10_wr[979]));
			radix2 #(.width(width)) rd_st9_980  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[980]), .rdlo_in(a9_wr[982]),  .coef_in(coef[0]), .rdup_out(a10_wr[980]), .rdlo_out(a10_wr[982]));
			radix2 #(.width(width)) rd_st9_981  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[981]), .rdlo_in(a9_wr[983]),  .coef_in(coef[512]), .rdup_out(a10_wr[981]), .rdlo_out(a10_wr[983]));
			radix2 #(.width(width)) rd_st9_984  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[984]), .rdlo_in(a9_wr[986]),  .coef_in(coef[0]), .rdup_out(a10_wr[984]), .rdlo_out(a10_wr[986]));
			radix2 #(.width(width)) rd_st9_985  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[985]), .rdlo_in(a9_wr[987]),  .coef_in(coef[512]), .rdup_out(a10_wr[985]), .rdlo_out(a10_wr[987]));
			radix2 #(.width(width)) rd_st9_988  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[988]), .rdlo_in(a9_wr[990]),  .coef_in(coef[0]), .rdup_out(a10_wr[988]), .rdlo_out(a10_wr[990]));
			radix2 #(.width(width)) rd_st9_989  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[989]), .rdlo_in(a9_wr[991]),  .coef_in(coef[512]), .rdup_out(a10_wr[989]), .rdlo_out(a10_wr[991]));
			radix2 #(.width(width)) rd_st9_992  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[992]), .rdlo_in(a9_wr[994]),  .coef_in(coef[0]), .rdup_out(a10_wr[992]), .rdlo_out(a10_wr[994]));
			radix2 #(.width(width)) rd_st9_993  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[993]), .rdlo_in(a9_wr[995]),  .coef_in(coef[512]), .rdup_out(a10_wr[993]), .rdlo_out(a10_wr[995]));
			radix2 #(.width(width)) rd_st9_996  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[996]), .rdlo_in(a9_wr[998]),  .coef_in(coef[0]), .rdup_out(a10_wr[996]), .rdlo_out(a10_wr[998]));
			radix2 #(.width(width)) rd_st9_997  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[997]), .rdlo_in(a9_wr[999]),  .coef_in(coef[512]), .rdup_out(a10_wr[997]), .rdlo_out(a10_wr[999]));
			radix2 #(.width(width)) rd_st9_1000  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1000]), .rdlo_in(a9_wr[1002]),  .coef_in(coef[0]), .rdup_out(a10_wr[1000]), .rdlo_out(a10_wr[1002]));
			radix2 #(.width(width)) rd_st9_1001  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1001]), .rdlo_in(a9_wr[1003]),  .coef_in(coef[512]), .rdup_out(a10_wr[1001]), .rdlo_out(a10_wr[1003]));
			radix2 #(.width(width)) rd_st9_1004  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1004]), .rdlo_in(a9_wr[1006]),  .coef_in(coef[0]), .rdup_out(a10_wr[1004]), .rdlo_out(a10_wr[1006]));
			radix2 #(.width(width)) rd_st9_1005  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1005]), .rdlo_in(a9_wr[1007]),  .coef_in(coef[512]), .rdup_out(a10_wr[1005]), .rdlo_out(a10_wr[1007]));
			radix2 #(.width(width)) rd_st9_1008  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1008]), .rdlo_in(a9_wr[1010]),  .coef_in(coef[0]), .rdup_out(a10_wr[1008]), .rdlo_out(a10_wr[1010]));
			radix2 #(.width(width)) rd_st9_1009  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1009]), .rdlo_in(a9_wr[1011]),  .coef_in(coef[512]), .rdup_out(a10_wr[1009]), .rdlo_out(a10_wr[1011]));
			radix2 #(.width(width)) rd_st9_1012  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1012]), .rdlo_in(a9_wr[1014]),  .coef_in(coef[0]), .rdup_out(a10_wr[1012]), .rdlo_out(a10_wr[1014]));
			radix2 #(.width(width)) rd_st9_1013  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1013]), .rdlo_in(a9_wr[1015]),  .coef_in(coef[512]), .rdup_out(a10_wr[1013]), .rdlo_out(a10_wr[1015]));
			radix2 #(.width(width)) rd_st9_1016  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1016]), .rdlo_in(a9_wr[1018]),  .coef_in(coef[0]), .rdup_out(a10_wr[1016]), .rdlo_out(a10_wr[1018]));
			radix2 #(.width(width)) rd_st9_1017  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1017]), .rdlo_in(a9_wr[1019]),  .coef_in(coef[512]), .rdup_out(a10_wr[1017]), .rdlo_out(a10_wr[1019]));
			radix2 #(.width(width)) rd_st9_1020  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1020]), .rdlo_in(a9_wr[1022]),  .coef_in(coef[0]), .rdup_out(a10_wr[1020]), .rdlo_out(a10_wr[1022]));
			radix2 #(.width(width)) rd_st9_1021  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1021]), .rdlo_in(a9_wr[1023]),  .coef_in(coef[512]), .rdup_out(a10_wr[1021]), .rdlo_out(a10_wr[1023]));
			radix2 #(.width(width)) rd_st9_1024  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1024]), .rdlo_in(a9_wr[1026]),  .coef_in(coef[0]), .rdup_out(a10_wr[1024]), .rdlo_out(a10_wr[1026]));
			radix2 #(.width(width)) rd_st9_1025  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1025]), .rdlo_in(a9_wr[1027]),  .coef_in(coef[512]), .rdup_out(a10_wr[1025]), .rdlo_out(a10_wr[1027]));
			radix2 #(.width(width)) rd_st9_1028  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1028]), .rdlo_in(a9_wr[1030]),  .coef_in(coef[0]), .rdup_out(a10_wr[1028]), .rdlo_out(a10_wr[1030]));
			radix2 #(.width(width)) rd_st9_1029  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1029]), .rdlo_in(a9_wr[1031]),  .coef_in(coef[512]), .rdup_out(a10_wr[1029]), .rdlo_out(a10_wr[1031]));
			radix2 #(.width(width)) rd_st9_1032  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1032]), .rdlo_in(a9_wr[1034]),  .coef_in(coef[0]), .rdup_out(a10_wr[1032]), .rdlo_out(a10_wr[1034]));
			radix2 #(.width(width)) rd_st9_1033  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1033]), .rdlo_in(a9_wr[1035]),  .coef_in(coef[512]), .rdup_out(a10_wr[1033]), .rdlo_out(a10_wr[1035]));
			radix2 #(.width(width)) rd_st9_1036  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1036]), .rdlo_in(a9_wr[1038]),  .coef_in(coef[0]), .rdup_out(a10_wr[1036]), .rdlo_out(a10_wr[1038]));
			radix2 #(.width(width)) rd_st9_1037  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1037]), .rdlo_in(a9_wr[1039]),  .coef_in(coef[512]), .rdup_out(a10_wr[1037]), .rdlo_out(a10_wr[1039]));
			radix2 #(.width(width)) rd_st9_1040  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1040]), .rdlo_in(a9_wr[1042]),  .coef_in(coef[0]), .rdup_out(a10_wr[1040]), .rdlo_out(a10_wr[1042]));
			radix2 #(.width(width)) rd_st9_1041  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1041]), .rdlo_in(a9_wr[1043]),  .coef_in(coef[512]), .rdup_out(a10_wr[1041]), .rdlo_out(a10_wr[1043]));
			radix2 #(.width(width)) rd_st9_1044  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1044]), .rdlo_in(a9_wr[1046]),  .coef_in(coef[0]), .rdup_out(a10_wr[1044]), .rdlo_out(a10_wr[1046]));
			radix2 #(.width(width)) rd_st9_1045  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1045]), .rdlo_in(a9_wr[1047]),  .coef_in(coef[512]), .rdup_out(a10_wr[1045]), .rdlo_out(a10_wr[1047]));
			radix2 #(.width(width)) rd_st9_1048  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1048]), .rdlo_in(a9_wr[1050]),  .coef_in(coef[0]), .rdup_out(a10_wr[1048]), .rdlo_out(a10_wr[1050]));
			radix2 #(.width(width)) rd_st9_1049  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1049]), .rdlo_in(a9_wr[1051]),  .coef_in(coef[512]), .rdup_out(a10_wr[1049]), .rdlo_out(a10_wr[1051]));
			radix2 #(.width(width)) rd_st9_1052  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1052]), .rdlo_in(a9_wr[1054]),  .coef_in(coef[0]), .rdup_out(a10_wr[1052]), .rdlo_out(a10_wr[1054]));
			radix2 #(.width(width)) rd_st9_1053  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1053]), .rdlo_in(a9_wr[1055]),  .coef_in(coef[512]), .rdup_out(a10_wr[1053]), .rdlo_out(a10_wr[1055]));
			radix2 #(.width(width)) rd_st9_1056  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1056]), .rdlo_in(a9_wr[1058]),  .coef_in(coef[0]), .rdup_out(a10_wr[1056]), .rdlo_out(a10_wr[1058]));
			radix2 #(.width(width)) rd_st9_1057  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1057]), .rdlo_in(a9_wr[1059]),  .coef_in(coef[512]), .rdup_out(a10_wr[1057]), .rdlo_out(a10_wr[1059]));
			radix2 #(.width(width)) rd_st9_1060  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1060]), .rdlo_in(a9_wr[1062]),  .coef_in(coef[0]), .rdup_out(a10_wr[1060]), .rdlo_out(a10_wr[1062]));
			radix2 #(.width(width)) rd_st9_1061  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1061]), .rdlo_in(a9_wr[1063]),  .coef_in(coef[512]), .rdup_out(a10_wr[1061]), .rdlo_out(a10_wr[1063]));
			radix2 #(.width(width)) rd_st9_1064  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1064]), .rdlo_in(a9_wr[1066]),  .coef_in(coef[0]), .rdup_out(a10_wr[1064]), .rdlo_out(a10_wr[1066]));
			radix2 #(.width(width)) rd_st9_1065  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1065]), .rdlo_in(a9_wr[1067]),  .coef_in(coef[512]), .rdup_out(a10_wr[1065]), .rdlo_out(a10_wr[1067]));
			radix2 #(.width(width)) rd_st9_1068  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1068]), .rdlo_in(a9_wr[1070]),  .coef_in(coef[0]), .rdup_out(a10_wr[1068]), .rdlo_out(a10_wr[1070]));
			radix2 #(.width(width)) rd_st9_1069  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1069]), .rdlo_in(a9_wr[1071]),  .coef_in(coef[512]), .rdup_out(a10_wr[1069]), .rdlo_out(a10_wr[1071]));
			radix2 #(.width(width)) rd_st9_1072  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1072]), .rdlo_in(a9_wr[1074]),  .coef_in(coef[0]), .rdup_out(a10_wr[1072]), .rdlo_out(a10_wr[1074]));
			radix2 #(.width(width)) rd_st9_1073  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1073]), .rdlo_in(a9_wr[1075]),  .coef_in(coef[512]), .rdup_out(a10_wr[1073]), .rdlo_out(a10_wr[1075]));
			radix2 #(.width(width)) rd_st9_1076  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1076]), .rdlo_in(a9_wr[1078]),  .coef_in(coef[0]), .rdup_out(a10_wr[1076]), .rdlo_out(a10_wr[1078]));
			radix2 #(.width(width)) rd_st9_1077  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1077]), .rdlo_in(a9_wr[1079]),  .coef_in(coef[512]), .rdup_out(a10_wr[1077]), .rdlo_out(a10_wr[1079]));
			radix2 #(.width(width)) rd_st9_1080  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1080]), .rdlo_in(a9_wr[1082]),  .coef_in(coef[0]), .rdup_out(a10_wr[1080]), .rdlo_out(a10_wr[1082]));
			radix2 #(.width(width)) rd_st9_1081  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1081]), .rdlo_in(a9_wr[1083]),  .coef_in(coef[512]), .rdup_out(a10_wr[1081]), .rdlo_out(a10_wr[1083]));
			radix2 #(.width(width)) rd_st9_1084  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1084]), .rdlo_in(a9_wr[1086]),  .coef_in(coef[0]), .rdup_out(a10_wr[1084]), .rdlo_out(a10_wr[1086]));
			radix2 #(.width(width)) rd_st9_1085  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1085]), .rdlo_in(a9_wr[1087]),  .coef_in(coef[512]), .rdup_out(a10_wr[1085]), .rdlo_out(a10_wr[1087]));
			radix2 #(.width(width)) rd_st9_1088  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1088]), .rdlo_in(a9_wr[1090]),  .coef_in(coef[0]), .rdup_out(a10_wr[1088]), .rdlo_out(a10_wr[1090]));
			radix2 #(.width(width)) rd_st9_1089  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1089]), .rdlo_in(a9_wr[1091]),  .coef_in(coef[512]), .rdup_out(a10_wr[1089]), .rdlo_out(a10_wr[1091]));
			radix2 #(.width(width)) rd_st9_1092  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1092]), .rdlo_in(a9_wr[1094]),  .coef_in(coef[0]), .rdup_out(a10_wr[1092]), .rdlo_out(a10_wr[1094]));
			radix2 #(.width(width)) rd_st9_1093  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1093]), .rdlo_in(a9_wr[1095]),  .coef_in(coef[512]), .rdup_out(a10_wr[1093]), .rdlo_out(a10_wr[1095]));
			radix2 #(.width(width)) rd_st9_1096  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1096]), .rdlo_in(a9_wr[1098]),  .coef_in(coef[0]), .rdup_out(a10_wr[1096]), .rdlo_out(a10_wr[1098]));
			radix2 #(.width(width)) rd_st9_1097  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1097]), .rdlo_in(a9_wr[1099]),  .coef_in(coef[512]), .rdup_out(a10_wr[1097]), .rdlo_out(a10_wr[1099]));
			radix2 #(.width(width)) rd_st9_1100  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1100]), .rdlo_in(a9_wr[1102]),  .coef_in(coef[0]), .rdup_out(a10_wr[1100]), .rdlo_out(a10_wr[1102]));
			radix2 #(.width(width)) rd_st9_1101  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1101]), .rdlo_in(a9_wr[1103]),  .coef_in(coef[512]), .rdup_out(a10_wr[1101]), .rdlo_out(a10_wr[1103]));
			radix2 #(.width(width)) rd_st9_1104  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1104]), .rdlo_in(a9_wr[1106]),  .coef_in(coef[0]), .rdup_out(a10_wr[1104]), .rdlo_out(a10_wr[1106]));
			radix2 #(.width(width)) rd_st9_1105  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1105]), .rdlo_in(a9_wr[1107]),  .coef_in(coef[512]), .rdup_out(a10_wr[1105]), .rdlo_out(a10_wr[1107]));
			radix2 #(.width(width)) rd_st9_1108  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1108]), .rdlo_in(a9_wr[1110]),  .coef_in(coef[0]), .rdup_out(a10_wr[1108]), .rdlo_out(a10_wr[1110]));
			radix2 #(.width(width)) rd_st9_1109  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1109]), .rdlo_in(a9_wr[1111]),  .coef_in(coef[512]), .rdup_out(a10_wr[1109]), .rdlo_out(a10_wr[1111]));
			radix2 #(.width(width)) rd_st9_1112  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1112]), .rdlo_in(a9_wr[1114]),  .coef_in(coef[0]), .rdup_out(a10_wr[1112]), .rdlo_out(a10_wr[1114]));
			radix2 #(.width(width)) rd_st9_1113  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1113]), .rdlo_in(a9_wr[1115]),  .coef_in(coef[512]), .rdup_out(a10_wr[1113]), .rdlo_out(a10_wr[1115]));
			radix2 #(.width(width)) rd_st9_1116  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1116]), .rdlo_in(a9_wr[1118]),  .coef_in(coef[0]), .rdup_out(a10_wr[1116]), .rdlo_out(a10_wr[1118]));
			radix2 #(.width(width)) rd_st9_1117  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1117]), .rdlo_in(a9_wr[1119]),  .coef_in(coef[512]), .rdup_out(a10_wr[1117]), .rdlo_out(a10_wr[1119]));
			radix2 #(.width(width)) rd_st9_1120  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1120]), .rdlo_in(a9_wr[1122]),  .coef_in(coef[0]), .rdup_out(a10_wr[1120]), .rdlo_out(a10_wr[1122]));
			radix2 #(.width(width)) rd_st9_1121  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1121]), .rdlo_in(a9_wr[1123]),  .coef_in(coef[512]), .rdup_out(a10_wr[1121]), .rdlo_out(a10_wr[1123]));
			radix2 #(.width(width)) rd_st9_1124  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1124]), .rdlo_in(a9_wr[1126]),  .coef_in(coef[0]), .rdup_out(a10_wr[1124]), .rdlo_out(a10_wr[1126]));
			radix2 #(.width(width)) rd_st9_1125  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1125]), .rdlo_in(a9_wr[1127]),  .coef_in(coef[512]), .rdup_out(a10_wr[1125]), .rdlo_out(a10_wr[1127]));
			radix2 #(.width(width)) rd_st9_1128  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1128]), .rdlo_in(a9_wr[1130]),  .coef_in(coef[0]), .rdup_out(a10_wr[1128]), .rdlo_out(a10_wr[1130]));
			radix2 #(.width(width)) rd_st9_1129  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1129]), .rdlo_in(a9_wr[1131]),  .coef_in(coef[512]), .rdup_out(a10_wr[1129]), .rdlo_out(a10_wr[1131]));
			radix2 #(.width(width)) rd_st9_1132  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1132]), .rdlo_in(a9_wr[1134]),  .coef_in(coef[0]), .rdup_out(a10_wr[1132]), .rdlo_out(a10_wr[1134]));
			radix2 #(.width(width)) rd_st9_1133  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1133]), .rdlo_in(a9_wr[1135]),  .coef_in(coef[512]), .rdup_out(a10_wr[1133]), .rdlo_out(a10_wr[1135]));
			radix2 #(.width(width)) rd_st9_1136  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1136]), .rdlo_in(a9_wr[1138]),  .coef_in(coef[0]), .rdup_out(a10_wr[1136]), .rdlo_out(a10_wr[1138]));
			radix2 #(.width(width)) rd_st9_1137  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1137]), .rdlo_in(a9_wr[1139]),  .coef_in(coef[512]), .rdup_out(a10_wr[1137]), .rdlo_out(a10_wr[1139]));
			radix2 #(.width(width)) rd_st9_1140  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1140]), .rdlo_in(a9_wr[1142]),  .coef_in(coef[0]), .rdup_out(a10_wr[1140]), .rdlo_out(a10_wr[1142]));
			radix2 #(.width(width)) rd_st9_1141  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1141]), .rdlo_in(a9_wr[1143]),  .coef_in(coef[512]), .rdup_out(a10_wr[1141]), .rdlo_out(a10_wr[1143]));
			radix2 #(.width(width)) rd_st9_1144  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1144]), .rdlo_in(a9_wr[1146]),  .coef_in(coef[0]), .rdup_out(a10_wr[1144]), .rdlo_out(a10_wr[1146]));
			radix2 #(.width(width)) rd_st9_1145  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1145]), .rdlo_in(a9_wr[1147]),  .coef_in(coef[512]), .rdup_out(a10_wr[1145]), .rdlo_out(a10_wr[1147]));
			radix2 #(.width(width)) rd_st9_1148  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1148]), .rdlo_in(a9_wr[1150]),  .coef_in(coef[0]), .rdup_out(a10_wr[1148]), .rdlo_out(a10_wr[1150]));
			radix2 #(.width(width)) rd_st9_1149  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1149]), .rdlo_in(a9_wr[1151]),  .coef_in(coef[512]), .rdup_out(a10_wr[1149]), .rdlo_out(a10_wr[1151]));
			radix2 #(.width(width)) rd_st9_1152  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1152]), .rdlo_in(a9_wr[1154]),  .coef_in(coef[0]), .rdup_out(a10_wr[1152]), .rdlo_out(a10_wr[1154]));
			radix2 #(.width(width)) rd_st9_1153  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1153]), .rdlo_in(a9_wr[1155]),  .coef_in(coef[512]), .rdup_out(a10_wr[1153]), .rdlo_out(a10_wr[1155]));
			radix2 #(.width(width)) rd_st9_1156  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1156]), .rdlo_in(a9_wr[1158]),  .coef_in(coef[0]), .rdup_out(a10_wr[1156]), .rdlo_out(a10_wr[1158]));
			radix2 #(.width(width)) rd_st9_1157  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1157]), .rdlo_in(a9_wr[1159]),  .coef_in(coef[512]), .rdup_out(a10_wr[1157]), .rdlo_out(a10_wr[1159]));
			radix2 #(.width(width)) rd_st9_1160  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1160]), .rdlo_in(a9_wr[1162]),  .coef_in(coef[0]), .rdup_out(a10_wr[1160]), .rdlo_out(a10_wr[1162]));
			radix2 #(.width(width)) rd_st9_1161  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1161]), .rdlo_in(a9_wr[1163]),  .coef_in(coef[512]), .rdup_out(a10_wr[1161]), .rdlo_out(a10_wr[1163]));
			radix2 #(.width(width)) rd_st9_1164  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1164]), .rdlo_in(a9_wr[1166]),  .coef_in(coef[0]), .rdup_out(a10_wr[1164]), .rdlo_out(a10_wr[1166]));
			radix2 #(.width(width)) rd_st9_1165  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1165]), .rdlo_in(a9_wr[1167]),  .coef_in(coef[512]), .rdup_out(a10_wr[1165]), .rdlo_out(a10_wr[1167]));
			radix2 #(.width(width)) rd_st9_1168  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1168]), .rdlo_in(a9_wr[1170]),  .coef_in(coef[0]), .rdup_out(a10_wr[1168]), .rdlo_out(a10_wr[1170]));
			radix2 #(.width(width)) rd_st9_1169  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1169]), .rdlo_in(a9_wr[1171]),  .coef_in(coef[512]), .rdup_out(a10_wr[1169]), .rdlo_out(a10_wr[1171]));
			radix2 #(.width(width)) rd_st9_1172  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1172]), .rdlo_in(a9_wr[1174]),  .coef_in(coef[0]), .rdup_out(a10_wr[1172]), .rdlo_out(a10_wr[1174]));
			radix2 #(.width(width)) rd_st9_1173  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1173]), .rdlo_in(a9_wr[1175]),  .coef_in(coef[512]), .rdup_out(a10_wr[1173]), .rdlo_out(a10_wr[1175]));
			radix2 #(.width(width)) rd_st9_1176  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1176]), .rdlo_in(a9_wr[1178]),  .coef_in(coef[0]), .rdup_out(a10_wr[1176]), .rdlo_out(a10_wr[1178]));
			radix2 #(.width(width)) rd_st9_1177  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1177]), .rdlo_in(a9_wr[1179]),  .coef_in(coef[512]), .rdup_out(a10_wr[1177]), .rdlo_out(a10_wr[1179]));
			radix2 #(.width(width)) rd_st9_1180  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1180]), .rdlo_in(a9_wr[1182]),  .coef_in(coef[0]), .rdup_out(a10_wr[1180]), .rdlo_out(a10_wr[1182]));
			radix2 #(.width(width)) rd_st9_1181  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1181]), .rdlo_in(a9_wr[1183]),  .coef_in(coef[512]), .rdup_out(a10_wr[1181]), .rdlo_out(a10_wr[1183]));
			radix2 #(.width(width)) rd_st9_1184  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1184]), .rdlo_in(a9_wr[1186]),  .coef_in(coef[0]), .rdup_out(a10_wr[1184]), .rdlo_out(a10_wr[1186]));
			radix2 #(.width(width)) rd_st9_1185  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1185]), .rdlo_in(a9_wr[1187]),  .coef_in(coef[512]), .rdup_out(a10_wr[1185]), .rdlo_out(a10_wr[1187]));
			radix2 #(.width(width)) rd_st9_1188  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1188]), .rdlo_in(a9_wr[1190]),  .coef_in(coef[0]), .rdup_out(a10_wr[1188]), .rdlo_out(a10_wr[1190]));
			radix2 #(.width(width)) rd_st9_1189  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1189]), .rdlo_in(a9_wr[1191]),  .coef_in(coef[512]), .rdup_out(a10_wr[1189]), .rdlo_out(a10_wr[1191]));
			radix2 #(.width(width)) rd_st9_1192  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1192]), .rdlo_in(a9_wr[1194]),  .coef_in(coef[0]), .rdup_out(a10_wr[1192]), .rdlo_out(a10_wr[1194]));
			radix2 #(.width(width)) rd_st9_1193  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1193]), .rdlo_in(a9_wr[1195]),  .coef_in(coef[512]), .rdup_out(a10_wr[1193]), .rdlo_out(a10_wr[1195]));
			radix2 #(.width(width)) rd_st9_1196  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1196]), .rdlo_in(a9_wr[1198]),  .coef_in(coef[0]), .rdup_out(a10_wr[1196]), .rdlo_out(a10_wr[1198]));
			radix2 #(.width(width)) rd_st9_1197  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1197]), .rdlo_in(a9_wr[1199]),  .coef_in(coef[512]), .rdup_out(a10_wr[1197]), .rdlo_out(a10_wr[1199]));
			radix2 #(.width(width)) rd_st9_1200  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1200]), .rdlo_in(a9_wr[1202]),  .coef_in(coef[0]), .rdup_out(a10_wr[1200]), .rdlo_out(a10_wr[1202]));
			radix2 #(.width(width)) rd_st9_1201  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1201]), .rdlo_in(a9_wr[1203]),  .coef_in(coef[512]), .rdup_out(a10_wr[1201]), .rdlo_out(a10_wr[1203]));
			radix2 #(.width(width)) rd_st9_1204  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1204]), .rdlo_in(a9_wr[1206]),  .coef_in(coef[0]), .rdup_out(a10_wr[1204]), .rdlo_out(a10_wr[1206]));
			radix2 #(.width(width)) rd_st9_1205  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1205]), .rdlo_in(a9_wr[1207]),  .coef_in(coef[512]), .rdup_out(a10_wr[1205]), .rdlo_out(a10_wr[1207]));
			radix2 #(.width(width)) rd_st9_1208  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1208]), .rdlo_in(a9_wr[1210]),  .coef_in(coef[0]), .rdup_out(a10_wr[1208]), .rdlo_out(a10_wr[1210]));
			radix2 #(.width(width)) rd_st9_1209  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1209]), .rdlo_in(a9_wr[1211]),  .coef_in(coef[512]), .rdup_out(a10_wr[1209]), .rdlo_out(a10_wr[1211]));
			radix2 #(.width(width)) rd_st9_1212  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1212]), .rdlo_in(a9_wr[1214]),  .coef_in(coef[0]), .rdup_out(a10_wr[1212]), .rdlo_out(a10_wr[1214]));
			radix2 #(.width(width)) rd_st9_1213  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1213]), .rdlo_in(a9_wr[1215]),  .coef_in(coef[512]), .rdup_out(a10_wr[1213]), .rdlo_out(a10_wr[1215]));
			radix2 #(.width(width)) rd_st9_1216  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1216]), .rdlo_in(a9_wr[1218]),  .coef_in(coef[0]), .rdup_out(a10_wr[1216]), .rdlo_out(a10_wr[1218]));
			radix2 #(.width(width)) rd_st9_1217  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1217]), .rdlo_in(a9_wr[1219]),  .coef_in(coef[512]), .rdup_out(a10_wr[1217]), .rdlo_out(a10_wr[1219]));
			radix2 #(.width(width)) rd_st9_1220  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1220]), .rdlo_in(a9_wr[1222]),  .coef_in(coef[0]), .rdup_out(a10_wr[1220]), .rdlo_out(a10_wr[1222]));
			radix2 #(.width(width)) rd_st9_1221  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1221]), .rdlo_in(a9_wr[1223]),  .coef_in(coef[512]), .rdup_out(a10_wr[1221]), .rdlo_out(a10_wr[1223]));
			radix2 #(.width(width)) rd_st9_1224  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1224]), .rdlo_in(a9_wr[1226]),  .coef_in(coef[0]), .rdup_out(a10_wr[1224]), .rdlo_out(a10_wr[1226]));
			radix2 #(.width(width)) rd_st9_1225  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1225]), .rdlo_in(a9_wr[1227]),  .coef_in(coef[512]), .rdup_out(a10_wr[1225]), .rdlo_out(a10_wr[1227]));
			radix2 #(.width(width)) rd_st9_1228  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1228]), .rdlo_in(a9_wr[1230]),  .coef_in(coef[0]), .rdup_out(a10_wr[1228]), .rdlo_out(a10_wr[1230]));
			radix2 #(.width(width)) rd_st9_1229  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1229]), .rdlo_in(a9_wr[1231]),  .coef_in(coef[512]), .rdup_out(a10_wr[1229]), .rdlo_out(a10_wr[1231]));
			radix2 #(.width(width)) rd_st9_1232  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1232]), .rdlo_in(a9_wr[1234]),  .coef_in(coef[0]), .rdup_out(a10_wr[1232]), .rdlo_out(a10_wr[1234]));
			radix2 #(.width(width)) rd_st9_1233  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1233]), .rdlo_in(a9_wr[1235]),  .coef_in(coef[512]), .rdup_out(a10_wr[1233]), .rdlo_out(a10_wr[1235]));
			radix2 #(.width(width)) rd_st9_1236  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1236]), .rdlo_in(a9_wr[1238]),  .coef_in(coef[0]), .rdup_out(a10_wr[1236]), .rdlo_out(a10_wr[1238]));
			radix2 #(.width(width)) rd_st9_1237  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1237]), .rdlo_in(a9_wr[1239]),  .coef_in(coef[512]), .rdup_out(a10_wr[1237]), .rdlo_out(a10_wr[1239]));
			radix2 #(.width(width)) rd_st9_1240  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1240]), .rdlo_in(a9_wr[1242]),  .coef_in(coef[0]), .rdup_out(a10_wr[1240]), .rdlo_out(a10_wr[1242]));
			radix2 #(.width(width)) rd_st9_1241  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1241]), .rdlo_in(a9_wr[1243]),  .coef_in(coef[512]), .rdup_out(a10_wr[1241]), .rdlo_out(a10_wr[1243]));
			radix2 #(.width(width)) rd_st9_1244  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1244]), .rdlo_in(a9_wr[1246]),  .coef_in(coef[0]), .rdup_out(a10_wr[1244]), .rdlo_out(a10_wr[1246]));
			radix2 #(.width(width)) rd_st9_1245  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1245]), .rdlo_in(a9_wr[1247]),  .coef_in(coef[512]), .rdup_out(a10_wr[1245]), .rdlo_out(a10_wr[1247]));
			radix2 #(.width(width)) rd_st9_1248  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1248]), .rdlo_in(a9_wr[1250]),  .coef_in(coef[0]), .rdup_out(a10_wr[1248]), .rdlo_out(a10_wr[1250]));
			radix2 #(.width(width)) rd_st9_1249  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1249]), .rdlo_in(a9_wr[1251]),  .coef_in(coef[512]), .rdup_out(a10_wr[1249]), .rdlo_out(a10_wr[1251]));
			radix2 #(.width(width)) rd_st9_1252  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1252]), .rdlo_in(a9_wr[1254]),  .coef_in(coef[0]), .rdup_out(a10_wr[1252]), .rdlo_out(a10_wr[1254]));
			radix2 #(.width(width)) rd_st9_1253  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1253]), .rdlo_in(a9_wr[1255]),  .coef_in(coef[512]), .rdup_out(a10_wr[1253]), .rdlo_out(a10_wr[1255]));
			radix2 #(.width(width)) rd_st9_1256  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1256]), .rdlo_in(a9_wr[1258]),  .coef_in(coef[0]), .rdup_out(a10_wr[1256]), .rdlo_out(a10_wr[1258]));
			radix2 #(.width(width)) rd_st9_1257  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1257]), .rdlo_in(a9_wr[1259]),  .coef_in(coef[512]), .rdup_out(a10_wr[1257]), .rdlo_out(a10_wr[1259]));
			radix2 #(.width(width)) rd_st9_1260  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1260]), .rdlo_in(a9_wr[1262]),  .coef_in(coef[0]), .rdup_out(a10_wr[1260]), .rdlo_out(a10_wr[1262]));
			radix2 #(.width(width)) rd_st9_1261  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1261]), .rdlo_in(a9_wr[1263]),  .coef_in(coef[512]), .rdup_out(a10_wr[1261]), .rdlo_out(a10_wr[1263]));
			radix2 #(.width(width)) rd_st9_1264  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1264]), .rdlo_in(a9_wr[1266]),  .coef_in(coef[0]), .rdup_out(a10_wr[1264]), .rdlo_out(a10_wr[1266]));
			radix2 #(.width(width)) rd_st9_1265  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1265]), .rdlo_in(a9_wr[1267]),  .coef_in(coef[512]), .rdup_out(a10_wr[1265]), .rdlo_out(a10_wr[1267]));
			radix2 #(.width(width)) rd_st9_1268  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1268]), .rdlo_in(a9_wr[1270]),  .coef_in(coef[0]), .rdup_out(a10_wr[1268]), .rdlo_out(a10_wr[1270]));
			radix2 #(.width(width)) rd_st9_1269  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1269]), .rdlo_in(a9_wr[1271]),  .coef_in(coef[512]), .rdup_out(a10_wr[1269]), .rdlo_out(a10_wr[1271]));
			radix2 #(.width(width)) rd_st9_1272  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1272]), .rdlo_in(a9_wr[1274]),  .coef_in(coef[0]), .rdup_out(a10_wr[1272]), .rdlo_out(a10_wr[1274]));
			radix2 #(.width(width)) rd_st9_1273  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1273]), .rdlo_in(a9_wr[1275]),  .coef_in(coef[512]), .rdup_out(a10_wr[1273]), .rdlo_out(a10_wr[1275]));
			radix2 #(.width(width)) rd_st9_1276  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1276]), .rdlo_in(a9_wr[1278]),  .coef_in(coef[0]), .rdup_out(a10_wr[1276]), .rdlo_out(a10_wr[1278]));
			radix2 #(.width(width)) rd_st9_1277  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1277]), .rdlo_in(a9_wr[1279]),  .coef_in(coef[512]), .rdup_out(a10_wr[1277]), .rdlo_out(a10_wr[1279]));
			radix2 #(.width(width)) rd_st9_1280  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1280]), .rdlo_in(a9_wr[1282]),  .coef_in(coef[0]), .rdup_out(a10_wr[1280]), .rdlo_out(a10_wr[1282]));
			radix2 #(.width(width)) rd_st9_1281  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1281]), .rdlo_in(a9_wr[1283]),  .coef_in(coef[512]), .rdup_out(a10_wr[1281]), .rdlo_out(a10_wr[1283]));
			radix2 #(.width(width)) rd_st9_1284  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1284]), .rdlo_in(a9_wr[1286]),  .coef_in(coef[0]), .rdup_out(a10_wr[1284]), .rdlo_out(a10_wr[1286]));
			radix2 #(.width(width)) rd_st9_1285  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1285]), .rdlo_in(a9_wr[1287]),  .coef_in(coef[512]), .rdup_out(a10_wr[1285]), .rdlo_out(a10_wr[1287]));
			radix2 #(.width(width)) rd_st9_1288  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1288]), .rdlo_in(a9_wr[1290]),  .coef_in(coef[0]), .rdup_out(a10_wr[1288]), .rdlo_out(a10_wr[1290]));
			radix2 #(.width(width)) rd_st9_1289  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1289]), .rdlo_in(a9_wr[1291]),  .coef_in(coef[512]), .rdup_out(a10_wr[1289]), .rdlo_out(a10_wr[1291]));
			radix2 #(.width(width)) rd_st9_1292  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1292]), .rdlo_in(a9_wr[1294]),  .coef_in(coef[0]), .rdup_out(a10_wr[1292]), .rdlo_out(a10_wr[1294]));
			radix2 #(.width(width)) rd_st9_1293  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1293]), .rdlo_in(a9_wr[1295]),  .coef_in(coef[512]), .rdup_out(a10_wr[1293]), .rdlo_out(a10_wr[1295]));
			radix2 #(.width(width)) rd_st9_1296  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1296]), .rdlo_in(a9_wr[1298]),  .coef_in(coef[0]), .rdup_out(a10_wr[1296]), .rdlo_out(a10_wr[1298]));
			radix2 #(.width(width)) rd_st9_1297  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1297]), .rdlo_in(a9_wr[1299]),  .coef_in(coef[512]), .rdup_out(a10_wr[1297]), .rdlo_out(a10_wr[1299]));
			radix2 #(.width(width)) rd_st9_1300  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1300]), .rdlo_in(a9_wr[1302]),  .coef_in(coef[0]), .rdup_out(a10_wr[1300]), .rdlo_out(a10_wr[1302]));
			radix2 #(.width(width)) rd_st9_1301  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1301]), .rdlo_in(a9_wr[1303]),  .coef_in(coef[512]), .rdup_out(a10_wr[1301]), .rdlo_out(a10_wr[1303]));
			radix2 #(.width(width)) rd_st9_1304  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1304]), .rdlo_in(a9_wr[1306]),  .coef_in(coef[0]), .rdup_out(a10_wr[1304]), .rdlo_out(a10_wr[1306]));
			radix2 #(.width(width)) rd_st9_1305  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1305]), .rdlo_in(a9_wr[1307]),  .coef_in(coef[512]), .rdup_out(a10_wr[1305]), .rdlo_out(a10_wr[1307]));
			radix2 #(.width(width)) rd_st9_1308  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1308]), .rdlo_in(a9_wr[1310]),  .coef_in(coef[0]), .rdup_out(a10_wr[1308]), .rdlo_out(a10_wr[1310]));
			radix2 #(.width(width)) rd_st9_1309  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1309]), .rdlo_in(a9_wr[1311]),  .coef_in(coef[512]), .rdup_out(a10_wr[1309]), .rdlo_out(a10_wr[1311]));
			radix2 #(.width(width)) rd_st9_1312  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1312]), .rdlo_in(a9_wr[1314]),  .coef_in(coef[0]), .rdup_out(a10_wr[1312]), .rdlo_out(a10_wr[1314]));
			radix2 #(.width(width)) rd_st9_1313  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1313]), .rdlo_in(a9_wr[1315]),  .coef_in(coef[512]), .rdup_out(a10_wr[1313]), .rdlo_out(a10_wr[1315]));
			radix2 #(.width(width)) rd_st9_1316  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1316]), .rdlo_in(a9_wr[1318]),  .coef_in(coef[0]), .rdup_out(a10_wr[1316]), .rdlo_out(a10_wr[1318]));
			radix2 #(.width(width)) rd_st9_1317  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1317]), .rdlo_in(a9_wr[1319]),  .coef_in(coef[512]), .rdup_out(a10_wr[1317]), .rdlo_out(a10_wr[1319]));
			radix2 #(.width(width)) rd_st9_1320  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1320]), .rdlo_in(a9_wr[1322]),  .coef_in(coef[0]), .rdup_out(a10_wr[1320]), .rdlo_out(a10_wr[1322]));
			radix2 #(.width(width)) rd_st9_1321  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1321]), .rdlo_in(a9_wr[1323]),  .coef_in(coef[512]), .rdup_out(a10_wr[1321]), .rdlo_out(a10_wr[1323]));
			radix2 #(.width(width)) rd_st9_1324  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1324]), .rdlo_in(a9_wr[1326]),  .coef_in(coef[0]), .rdup_out(a10_wr[1324]), .rdlo_out(a10_wr[1326]));
			radix2 #(.width(width)) rd_st9_1325  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1325]), .rdlo_in(a9_wr[1327]),  .coef_in(coef[512]), .rdup_out(a10_wr[1325]), .rdlo_out(a10_wr[1327]));
			radix2 #(.width(width)) rd_st9_1328  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1328]), .rdlo_in(a9_wr[1330]),  .coef_in(coef[0]), .rdup_out(a10_wr[1328]), .rdlo_out(a10_wr[1330]));
			radix2 #(.width(width)) rd_st9_1329  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1329]), .rdlo_in(a9_wr[1331]),  .coef_in(coef[512]), .rdup_out(a10_wr[1329]), .rdlo_out(a10_wr[1331]));
			radix2 #(.width(width)) rd_st9_1332  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1332]), .rdlo_in(a9_wr[1334]),  .coef_in(coef[0]), .rdup_out(a10_wr[1332]), .rdlo_out(a10_wr[1334]));
			radix2 #(.width(width)) rd_st9_1333  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1333]), .rdlo_in(a9_wr[1335]),  .coef_in(coef[512]), .rdup_out(a10_wr[1333]), .rdlo_out(a10_wr[1335]));
			radix2 #(.width(width)) rd_st9_1336  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1336]), .rdlo_in(a9_wr[1338]),  .coef_in(coef[0]), .rdup_out(a10_wr[1336]), .rdlo_out(a10_wr[1338]));
			radix2 #(.width(width)) rd_st9_1337  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1337]), .rdlo_in(a9_wr[1339]),  .coef_in(coef[512]), .rdup_out(a10_wr[1337]), .rdlo_out(a10_wr[1339]));
			radix2 #(.width(width)) rd_st9_1340  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1340]), .rdlo_in(a9_wr[1342]),  .coef_in(coef[0]), .rdup_out(a10_wr[1340]), .rdlo_out(a10_wr[1342]));
			radix2 #(.width(width)) rd_st9_1341  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1341]), .rdlo_in(a9_wr[1343]),  .coef_in(coef[512]), .rdup_out(a10_wr[1341]), .rdlo_out(a10_wr[1343]));
			radix2 #(.width(width)) rd_st9_1344  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1344]), .rdlo_in(a9_wr[1346]),  .coef_in(coef[0]), .rdup_out(a10_wr[1344]), .rdlo_out(a10_wr[1346]));
			radix2 #(.width(width)) rd_st9_1345  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1345]), .rdlo_in(a9_wr[1347]),  .coef_in(coef[512]), .rdup_out(a10_wr[1345]), .rdlo_out(a10_wr[1347]));
			radix2 #(.width(width)) rd_st9_1348  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1348]), .rdlo_in(a9_wr[1350]),  .coef_in(coef[0]), .rdup_out(a10_wr[1348]), .rdlo_out(a10_wr[1350]));
			radix2 #(.width(width)) rd_st9_1349  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1349]), .rdlo_in(a9_wr[1351]),  .coef_in(coef[512]), .rdup_out(a10_wr[1349]), .rdlo_out(a10_wr[1351]));
			radix2 #(.width(width)) rd_st9_1352  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1352]), .rdlo_in(a9_wr[1354]),  .coef_in(coef[0]), .rdup_out(a10_wr[1352]), .rdlo_out(a10_wr[1354]));
			radix2 #(.width(width)) rd_st9_1353  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1353]), .rdlo_in(a9_wr[1355]),  .coef_in(coef[512]), .rdup_out(a10_wr[1353]), .rdlo_out(a10_wr[1355]));
			radix2 #(.width(width)) rd_st9_1356  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1356]), .rdlo_in(a9_wr[1358]),  .coef_in(coef[0]), .rdup_out(a10_wr[1356]), .rdlo_out(a10_wr[1358]));
			radix2 #(.width(width)) rd_st9_1357  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1357]), .rdlo_in(a9_wr[1359]),  .coef_in(coef[512]), .rdup_out(a10_wr[1357]), .rdlo_out(a10_wr[1359]));
			radix2 #(.width(width)) rd_st9_1360  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1360]), .rdlo_in(a9_wr[1362]),  .coef_in(coef[0]), .rdup_out(a10_wr[1360]), .rdlo_out(a10_wr[1362]));
			radix2 #(.width(width)) rd_st9_1361  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1361]), .rdlo_in(a9_wr[1363]),  .coef_in(coef[512]), .rdup_out(a10_wr[1361]), .rdlo_out(a10_wr[1363]));
			radix2 #(.width(width)) rd_st9_1364  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1364]), .rdlo_in(a9_wr[1366]),  .coef_in(coef[0]), .rdup_out(a10_wr[1364]), .rdlo_out(a10_wr[1366]));
			radix2 #(.width(width)) rd_st9_1365  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1365]), .rdlo_in(a9_wr[1367]),  .coef_in(coef[512]), .rdup_out(a10_wr[1365]), .rdlo_out(a10_wr[1367]));
			radix2 #(.width(width)) rd_st9_1368  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1368]), .rdlo_in(a9_wr[1370]),  .coef_in(coef[0]), .rdup_out(a10_wr[1368]), .rdlo_out(a10_wr[1370]));
			radix2 #(.width(width)) rd_st9_1369  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1369]), .rdlo_in(a9_wr[1371]),  .coef_in(coef[512]), .rdup_out(a10_wr[1369]), .rdlo_out(a10_wr[1371]));
			radix2 #(.width(width)) rd_st9_1372  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1372]), .rdlo_in(a9_wr[1374]),  .coef_in(coef[0]), .rdup_out(a10_wr[1372]), .rdlo_out(a10_wr[1374]));
			radix2 #(.width(width)) rd_st9_1373  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1373]), .rdlo_in(a9_wr[1375]),  .coef_in(coef[512]), .rdup_out(a10_wr[1373]), .rdlo_out(a10_wr[1375]));
			radix2 #(.width(width)) rd_st9_1376  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1376]), .rdlo_in(a9_wr[1378]),  .coef_in(coef[0]), .rdup_out(a10_wr[1376]), .rdlo_out(a10_wr[1378]));
			radix2 #(.width(width)) rd_st9_1377  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1377]), .rdlo_in(a9_wr[1379]),  .coef_in(coef[512]), .rdup_out(a10_wr[1377]), .rdlo_out(a10_wr[1379]));
			radix2 #(.width(width)) rd_st9_1380  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1380]), .rdlo_in(a9_wr[1382]),  .coef_in(coef[0]), .rdup_out(a10_wr[1380]), .rdlo_out(a10_wr[1382]));
			radix2 #(.width(width)) rd_st9_1381  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1381]), .rdlo_in(a9_wr[1383]),  .coef_in(coef[512]), .rdup_out(a10_wr[1381]), .rdlo_out(a10_wr[1383]));
			radix2 #(.width(width)) rd_st9_1384  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1384]), .rdlo_in(a9_wr[1386]),  .coef_in(coef[0]), .rdup_out(a10_wr[1384]), .rdlo_out(a10_wr[1386]));
			radix2 #(.width(width)) rd_st9_1385  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1385]), .rdlo_in(a9_wr[1387]),  .coef_in(coef[512]), .rdup_out(a10_wr[1385]), .rdlo_out(a10_wr[1387]));
			radix2 #(.width(width)) rd_st9_1388  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1388]), .rdlo_in(a9_wr[1390]),  .coef_in(coef[0]), .rdup_out(a10_wr[1388]), .rdlo_out(a10_wr[1390]));
			radix2 #(.width(width)) rd_st9_1389  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1389]), .rdlo_in(a9_wr[1391]),  .coef_in(coef[512]), .rdup_out(a10_wr[1389]), .rdlo_out(a10_wr[1391]));
			radix2 #(.width(width)) rd_st9_1392  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1392]), .rdlo_in(a9_wr[1394]),  .coef_in(coef[0]), .rdup_out(a10_wr[1392]), .rdlo_out(a10_wr[1394]));
			radix2 #(.width(width)) rd_st9_1393  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1393]), .rdlo_in(a9_wr[1395]),  .coef_in(coef[512]), .rdup_out(a10_wr[1393]), .rdlo_out(a10_wr[1395]));
			radix2 #(.width(width)) rd_st9_1396  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1396]), .rdlo_in(a9_wr[1398]),  .coef_in(coef[0]), .rdup_out(a10_wr[1396]), .rdlo_out(a10_wr[1398]));
			radix2 #(.width(width)) rd_st9_1397  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1397]), .rdlo_in(a9_wr[1399]),  .coef_in(coef[512]), .rdup_out(a10_wr[1397]), .rdlo_out(a10_wr[1399]));
			radix2 #(.width(width)) rd_st9_1400  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1400]), .rdlo_in(a9_wr[1402]),  .coef_in(coef[0]), .rdup_out(a10_wr[1400]), .rdlo_out(a10_wr[1402]));
			radix2 #(.width(width)) rd_st9_1401  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1401]), .rdlo_in(a9_wr[1403]),  .coef_in(coef[512]), .rdup_out(a10_wr[1401]), .rdlo_out(a10_wr[1403]));
			radix2 #(.width(width)) rd_st9_1404  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1404]), .rdlo_in(a9_wr[1406]),  .coef_in(coef[0]), .rdup_out(a10_wr[1404]), .rdlo_out(a10_wr[1406]));
			radix2 #(.width(width)) rd_st9_1405  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1405]), .rdlo_in(a9_wr[1407]),  .coef_in(coef[512]), .rdup_out(a10_wr[1405]), .rdlo_out(a10_wr[1407]));
			radix2 #(.width(width)) rd_st9_1408  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1408]), .rdlo_in(a9_wr[1410]),  .coef_in(coef[0]), .rdup_out(a10_wr[1408]), .rdlo_out(a10_wr[1410]));
			radix2 #(.width(width)) rd_st9_1409  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1409]), .rdlo_in(a9_wr[1411]),  .coef_in(coef[512]), .rdup_out(a10_wr[1409]), .rdlo_out(a10_wr[1411]));
			radix2 #(.width(width)) rd_st9_1412  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1412]), .rdlo_in(a9_wr[1414]),  .coef_in(coef[0]), .rdup_out(a10_wr[1412]), .rdlo_out(a10_wr[1414]));
			radix2 #(.width(width)) rd_st9_1413  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1413]), .rdlo_in(a9_wr[1415]),  .coef_in(coef[512]), .rdup_out(a10_wr[1413]), .rdlo_out(a10_wr[1415]));
			radix2 #(.width(width)) rd_st9_1416  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1416]), .rdlo_in(a9_wr[1418]),  .coef_in(coef[0]), .rdup_out(a10_wr[1416]), .rdlo_out(a10_wr[1418]));
			radix2 #(.width(width)) rd_st9_1417  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1417]), .rdlo_in(a9_wr[1419]),  .coef_in(coef[512]), .rdup_out(a10_wr[1417]), .rdlo_out(a10_wr[1419]));
			radix2 #(.width(width)) rd_st9_1420  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1420]), .rdlo_in(a9_wr[1422]),  .coef_in(coef[0]), .rdup_out(a10_wr[1420]), .rdlo_out(a10_wr[1422]));
			radix2 #(.width(width)) rd_st9_1421  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1421]), .rdlo_in(a9_wr[1423]),  .coef_in(coef[512]), .rdup_out(a10_wr[1421]), .rdlo_out(a10_wr[1423]));
			radix2 #(.width(width)) rd_st9_1424  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1424]), .rdlo_in(a9_wr[1426]),  .coef_in(coef[0]), .rdup_out(a10_wr[1424]), .rdlo_out(a10_wr[1426]));
			radix2 #(.width(width)) rd_st9_1425  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1425]), .rdlo_in(a9_wr[1427]),  .coef_in(coef[512]), .rdup_out(a10_wr[1425]), .rdlo_out(a10_wr[1427]));
			radix2 #(.width(width)) rd_st9_1428  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1428]), .rdlo_in(a9_wr[1430]),  .coef_in(coef[0]), .rdup_out(a10_wr[1428]), .rdlo_out(a10_wr[1430]));
			radix2 #(.width(width)) rd_st9_1429  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1429]), .rdlo_in(a9_wr[1431]),  .coef_in(coef[512]), .rdup_out(a10_wr[1429]), .rdlo_out(a10_wr[1431]));
			radix2 #(.width(width)) rd_st9_1432  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1432]), .rdlo_in(a9_wr[1434]),  .coef_in(coef[0]), .rdup_out(a10_wr[1432]), .rdlo_out(a10_wr[1434]));
			radix2 #(.width(width)) rd_st9_1433  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1433]), .rdlo_in(a9_wr[1435]),  .coef_in(coef[512]), .rdup_out(a10_wr[1433]), .rdlo_out(a10_wr[1435]));
			radix2 #(.width(width)) rd_st9_1436  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1436]), .rdlo_in(a9_wr[1438]),  .coef_in(coef[0]), .rdup_out(a10_wr[1436]), .rdlo_out(a10_wr[1438]));
			radix2 #(.width(width)) rd_st9_1437  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1437]), .rdlo_in(a9_wr[1439]),  .coef_in(coef[512]), .rdup_out(a10_wr[1437]), .rdlo_out(a10_wr[1439]));
			radix2 #(.width(width)) rd_st9_1440  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1440]), .rdlo_in(a9_wr[1442]),  .coef_in(coef[0]), .rdup_out(a10_wr[1440]), .rdlo_out(a10_wr[1442]));
			radix2 #(.width(width)) rd_st9_1441  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1441]), .rdlo_in(a9_wr[1443]),  .coef_in(coef[512]), .rdup_out(a10_wr[1441]), .rdlo_out(a10_wr[1443]));
			radix2 #(.width(width)) rd_st9_1444  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1444]), .rdlo_in(a9_wr[1446]),  .coef_in(coef[0]), .rdup_out(a10_wr[1444]), .rdlo_out(a10_wr[1446]));
			radix2 #(.width(width)) rd_st9_1445  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1445]), .rdlo_in(a9_wr[1447]),  .coef_in(coef[512]), .rdup_out(a10_wr[1445]), .rdlo_out(a10_wr[1447]));
			radix2 #(.width(width)) rd_st9_1448  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1448]), .rdlo_in(a9_wr[1450]),  .coef_in(coef[0]), .rdup_out(a10_wr[1448]), .rdlo_out(a10_wr[1450]));
			radix2 #(.width(width)) rd_st9_1449  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1449]), .rdlo_in(a9_wr[1451]),  .coef_in(coef[512]), .rdup_out(a10_wr[1449]), .rdlo_out(a10_wr[1451]));
			radix2 #(.width(width)) rd_st9_1452  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1452]), .rdlo_in(a9_wr[1454]),  .coef_in(coef[0]), .rdup_out(a10_wr[1452]), .rdlo_out(a10_wr[1454]));
			radix2 #(.width(width)) rd_st9_1453  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1453]), .rdlo_in(a9_wr[1455]),  .coef_in(coef[512]), .rdup_out(a10_wr[1453]), .rdlo_out(a10_wr[1455]));
			radix2 #(.width(width)) rd_st9_1456  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1456]), .rdlo_in(a9_wr[1458]),  .coef_in(coef[0]), .rdup_out(a10_wr[1456]), .rdlo_out(a10_wr[1458]));
			radix2 #(.width(width)) rd_st9_1457  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1457]), .rdlo_in(a9_wr[1459]),  .coef_in(coef[512]), .rdup_out(a10_wr[1457]), .rdlo_out(a10_wr[1459]));
			radix2 #(.width(width)) rd_st9_1460  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1460]), .rdlo_in(a9_wr[1462]),  .coef_in(coef[0]), .rdup_out(a10_wr[1460]), .rdlo_out(a10_wr[1462]));
			radix2 #(.width(width)) rd_st9_1461  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1461]), .rdlo_in(a9_wr[1463]),  .coef_in(coef[512]), .rdup_out(a10_wr[1461]), .rdlo_out(a10_wr[1463]));
			radix2 #(.width(width)) rd_st9_1464  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1464]), .rdlo_in(a9_wr[1466]),  .coef_in(coef[0]), .rdup_out(a10_wr[1464]), .rdlo_out(a10_wr[1466]));
			radix2 #(.width(width)) rd_st9_1465  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1465]), .rdlo_in(a9_wr[1467]),  .coef_in(coef[512]), .rdup_out(a10_wr[1465]), .rdlo_out(a10_wr[1467]));
			radix2 #(.width(width)) rd_st9_1468  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1468]), .rdlo_in(a9_wr[1470]),  .coef_in(coef[0]), .rdup_out(a10_wr[1468]), .rdlo_out(a10_wr[1470]));
			radix2 #(.width(width)) rd_st9_1469  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1469]), .rdlo_in(a9_wr[1471]),  .coef_in(coef[512]), .rdup_out(a10_wr[1469]), .rdlo_out(a10_wr[1471]));
			radix2 #(.width(width)) rd_st9_1472  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1472]), .rdlo_in(a9_wr[1474]),  .coef_in(coef[0]), .rdup_out(a10_wr[1472]), .rdlo_out(a10_wr[1474]));
			radix2 #(.width(width)) rd_st9_1473  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1473]), .rdlo_in(a9_wr[1475]),  .coef_in(coef[512]), .rdup_out(a10_wr[1473]), .rdlo_out(a10_wr[1475]));
			radix2 #(.width(width)) rd_st9_1476  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1476]), .rdlo_in(a9_wr[1478]),  .coef_in(coef[0]), .rdup_out(a10_wr[1476]), .rdlo_out(a10_wr[1478]));
			radix2 #(.width(width)) rd_st9_1477  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1477]), .rdlo_in(a9_wr[1479]),  .coef_in(coef[512]), .rdup_out(a10_wr[1477]), .rdlo_out(a10_wr[1479]));
			radix2 #(.width(width)) rd_st9_1480  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1480]), .rdlo_in(a9_wr[1482]),  .coef_in(coef[0]), .rdup_out(a10_wr[1480]), .rdlo_out(a10_wr[1482]));
			radix2 #(.width(width)) rd_st9_1481  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1481]), .rdlo_in(a9_wr[1483]),  .coef_in(coef[512]), .rdup_out(a10_wr[1481]), .rdlo_out(a10_wr[1483]));
			radix2 #(.width(width)) rd_st9_1484  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1484]), .rdlo_in(a9_wr[1486]),  .coef_in(coef[0]), .rdup_out(a10_wr[1484]), .rdlo_out(a10_wr[1486]));
			radix2 #(.width(width)) rd_st9_1485  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1485]), .rdlo_in(a9_wr[1487]),  .coef_in(coef[512]), .rdup_out(a10_wr[1485]), .rdlo_out(a10_wr[1487]));
			radix2 #(.width(width)) rd_st9_1488  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1488]), .rdlo_in(a9_wr[1490]),  .coef_in(coef[0]), .rdup_out(a10_wr[1488]), .rdlo_out(a10_wr[1490]));
			radix2 #(.width(width)) rd_st9_1489  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1489]), .rdlo_in(a9_wr[1491]),  .coef_in(coef[512]), .rdup_out(a10_wr[1489]), .rdlo_out(a10_wr[1491]));
			radix2 #(.width(width)) rd_st9_1492  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1492]), .rdlo_in(a9_wr[1494]),  .coef_in(coef[0]), .rdup_out(a10_wr[1492]), .rdlo_out(a10_wr[1494]));
			radix2 #(.width(width)) rd_st9_1493  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1493]), .rdlo_in(a9_wr[1495]),  .coef_in(coef[512]), .rdup_out(a10_wr[1493]), .rdlo_out(a10_wr[1495]));
			radix2 #(.width(width)) rd_st9_1496  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1496]), .rdlo_in(a9_wr[1498]),  .coef_in(coef[0]), .rdup_out(a10_wr[1496]), .rdlo_out(a10_wr[1498]));
			radix2 #(.width(width)) rd_st9_1497  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1497]), .rdlo_in(a9_wr[1499]),  .coef_in(coef[512]), .rdup_out(a10_wr[1497]), .rdlo_out(a10_wr[1499]));
			radix2 #(.width(width)) rd_st9_1500  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1500]), .rdlo_in(a9_wr[1502]),  .coef_in(coef[0]), .rdup_out(a10_wr[1500]), .rdlo_out(a10_wr[1502]));
			radix2 #(.width(width)) rd_st9_1501  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1501]), .rdlo_in(a9_wr[1503]),  .coef_in(coef[512]), .rdup_out(a10_wr[1501]), .rdlo_out(a10_wr[1503]));
			radix2 #(.width(width)) rd_st9_1504  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1504]), .rdlo_in(a9_wr[1506]),  .coef_in(coef[0]), .rdup_out(a10_wr[1504]), .rdlo_out(a10_wr[1506]));
			radix2 #(.width(width)) rd_st9_1505  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1505]), .rdlo_in(a9_wr[1507]),  .coef_in(coef[512]), .rdup_out(a10_wr[1505]), .rdlo_out(a10_wr[1507]));
			radix2 #(.width(width)) rd_st9_1508  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1508]), .rdlo_in(a9_wr[1510]),  .coef_in(coef[0]), .rdup_out(a10_wr[1508]), .rdlo_out(a10_wr[1510]));
			radix2 #(.width(width)) rd_st9_1509  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1509]), .rdlo_in(a9_wr[1511]),  .coef_in(coef[512]), .rdup_out(a10_wr[1509]), .rdlo_out(a10_wr[1511]));
			radix2 #(.width(width)) rd_st9_1512  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1512]), .rdlo_in(a9_wr[1514]),  .coef_in(coef[0]), .rdup_out(a10_wr[1512]), .rdlo_out(a10_wr[1514]));
			radix2 #(.width(width)) rd_st9_1513  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1513]), .rdlo_in(a9_wr[1515]),  .coef_in(coef[512]), .rdup_out(a10_wr[1513]), .rdlo_out(a10_wr[1515]));
			radix2 #(.width(width)) rd_st9_1516  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1516]), .rdlo_in(a9_wr[1518]),  .coef_in(coef[0]), .rdup_out(a10_wr[1516]), .rdlo_out(a10_wr[1518]));
			radix2 #(.width(width)) rd_st9_1517  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1517]), .rdlo_in(a9_wr[1519]),  .coef_in(coef[512]), .rdup_out(a10_wr[1517]), .rdlo_out(a10_wr[1519]));
			radix2 #(.width(width)) rd_st9_1520  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1520]), .rdlo_in(a9_wr[1522]),  .coef_in(coef[0]), .rdup_out(a10_wr[1520]), .rdlo_out(a10_wr[1522]));
			radix2 #(.width(width)) rd_st9_1521  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1521]), .rdlo_in(a9_wr[1523]),  .coef_in(coef[512]), .rdup_out(a10_wr[1521]), .rdlo_out(a10_wr[1523]));
			radix2 #(.width(width)) rd_st9_1524  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1524]), .rdlo_in(a9_wr[1526]),  .coef_in(coef[0]), .rdup_out(a10_wr[1524]), .rdlo_out(a10_wr[1526]));
			radix2 #(.width(width)) rd_st9_1525  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1525]), .rdlo_in(a9_wr[1527]),  .coef_in(coef[512]), .rdup_out(a10_wr[1525]), .rdlo_out(a10_wr[1527]));
			radix2 #(.width(width)) rd_st9_1528  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1528]), .rdlo_in(a9_wr[1530]),  .coef_in(coef[0]), .rdup_out(a10_wr[1528]), .rdlo_out(a10_wr[1530]));
			radix2 #(.width(width)) rd_st9_1529  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1529]), .rdlo_in(a9_wr[1531]),  .coef_in(coef[512]), .rdup_out(a10_wr[1529]), .rdlo_out(a10_wr[1531]));
			radix2 #(.width(width)) rd_st9_1532  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1532]), .rdlo_in(a9_wr[1534]),  .coef_in(coef[0]), .rdup_out(a10_wr[1532]), .rdlo_out(a10_wr[1534]));
			radix2 #(.width(width)) rd_st9_1533  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1533]), .rdlo_in(a9_wr[1535]),  .coef_in(coef[512]), .rdup_out(a10_wr[1533]), .rdlo_out(a10_wr[1535]));
			radix2 #(.width(width)) rd_st9_1536  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1536]), .rdlo_in(a9_wr[1538]),  .coef_in(coef[0]), .rdup_out(a10_wr[1536]), .rdlo_out(a10_wr[1538]));
			radix2 #(.width(width)) rd_st9_1537  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1537]), .rdlo_in(a9_wr[1539]),  .coef_in(coef[512]), .rdup_out(a10_wr[1537]), .rdlo_out(a10_wr[1539]));
			radix2 #(.width(width)) rd_st9_1540  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1540]), .rdlo_in(a9_wr[1542]),  .coef_in(coef[0]), .rdup_out(a10_wr[1540]), .rdlo_out(a10_wr[1542]));
			radix2 #(.width(width)) rd_st9_1541  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1541]), .rdlo_in(a9_wr[1543]),  .coef_in(coef[512]), .rdup_out(a10_wr[1541]), .rdlo_out(a10_wr[1543]));
			radix2 #(.width(width)) rd_st9_1544  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1544]), .rdlo_in(a9_wr[1546]),  .coef_in(coef[0]), .rdup_out(a10_wr[1544]), .rdlo_out(a10_wr[1546]));
			radix2 #(.width(width)) rd_st9_1545  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1545]), .rdlo_in(a9_wr[1547]),  .coef_in(coef[512]), .rdup_out(a10_wr[1545]), .rdlo_out(a10_wr[1547]));
			radix2 #(.width(width)) rd_st9_1548  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1548]), .rdlo_in(a9_wr[1550]),  .coef_in(coef[0]), .rdup_out(a10_wr[1548]), .rdlo_out(a10_wr[1550]));
			radix2 #(.width(width)) rd_st9_1549  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1549]), .rdlo_in(a9_wr[1551]),  .coef_in(coef[512]), .rdup_out(a10_wr[1549]), .rdlo_out(a10_wr[1551]));
			radix2 #(.width(width)) rd_st9_1552  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1552]), .rdlo_in(a9_wr[1554]),  .coef_in(coef[0]), .rdup_out(a10_wr[1552]), .rdlo_out(a10_wr[1554]));
			radix2 #(.width(width)) rd_st9_1553  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1553]), .rdlo_in(a9_wr[1555]),  .coef_in(coef[512]), .rdup_out(a10_wr[1553]), .rdlo_out(a10_wr[1555]));
			radix2 #(.width(width)) rd_st9_1556  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1556]), .rdlo_in(a9_wr[1558]),  .coef_in(coef[0]), .rdup_out(a10_wr[1556]), .rdlo_out(a10_wr[1558]));
			radix2 #(.width(width)) rd_st9_1557  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1557]), .rdlo_in(a9_wr[1559]),  .coef_in(coef[512]), .rdup_out(a10_wr[1557]), .rdlo_out(a10_wr[1559]));
			radix2 #(.width(width)) rd_st9_1560  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1560]), .rdlo_in(a9_wr[1562]),  .coef_in(coef[0]), .rdup_out(a10_wr[1560]), .rdlo_out(a10_wr[1562]));
			radix2 #(.width(width)) rd_st9_1561  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1561]), .rdlo_in(a9_wr[1563]),  .coef_in(coef[512]), .rdup_out(a10_wr[1561]), .rdlo_out(a10_wr[1563]));
			radix2 #(.width(width)) rd_st9_1564  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1564]), .rdlo_in(a9_wr[1566]),  .coef_in(coef[0]), .rdup_out(a10_wr[1564]), .rdlo_out(a10_wr[1566]));
			radix2 #(.width(width)) rd_st9_1565  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1565]), .rdlo_in(a9_wr[1567]),  .coef_in(coef[512]), .rdup_out(a10_wr[1565]), .rdlo_out(a10_wr[1567]));
			radix2 #(.width(width)) rd_st9_1568  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1568]), .rdlo_in(a9_wr[1570]),  .coef_in(coef[0]), .rdup_out(a10_wr[1568]), .rdlo_out(a10_wr[1570]));
			radix2 #(.width(width)) rd_st9_1569  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1569]), .rdlo_in(a9_wr[1571]),  .coef_in(coef[512]), .rdup_out(a10_wr[1569]), .rdlo_out(a10_wr[1571]));
			radix2 #(.width(width)) rd_st9_1572  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1572]), .rdlo_in(a9_wr[1574]),  .coef_in(coef[0]), .rdup_out(a10_wr[1572]), .rdlo_out(a10_wr[1574]));
			radix2 #(.width(width)) rd_st9_1573  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1573]), .rdlo_in(a9_wr[1575]),  .coef_in(coef[512]), .rdup_out(a10_wr[1573]), .rdlo_out(a10_wr[1575]));
			radix2 #(.width(width)) rd_st9_1576  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1576]), .rdlo_in(a9_wr[1578]),  .coef_in(coef[0]), .rdup_out(a10_wr[1576]), .rdlo_out(a10_wr[1578]));
			radix2 #(.width(width)) rd_st9_1577  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1577]), .rdlo_in(a9_wr[1579]),  .coef_in(coef[512]), .rdup_out(a10_wr[1577]), .rdlo_out(a10_wr[1579]));
			radix2 #(.width(width)) rd_st9_1580  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1580]), .rdlo_in(a9_wr[1582]),  .coef_in(coef[0]), .rdup_out(a10_wr[1580]), .rdlo_out(a10_wr[1582]));
			radix2 #(.width(width)) rd_st9_1581  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1581]), .rdlo_in(a9_wr[1583]),  .coef_in(coef[512]), .rdup_out(a10_wr[1581]), .rdlo_out(a10_wr[1583]));
			radix2 #(.width(width)) rd_st9_1584  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1584]), .rdlo_in(a9_wr[1586]),  .coef_in(coef[0]), .rdup_out(a10_wr[1584]), .rdlo_out(a10_wr[1586]));
			radix2 #(.width(width)) rd_st9_1585  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1585]), .rdlo_in(a9_wr[1587]),  .coef_in(coef[512]), .rdup_out(a10_wr[1585]), .rdlo_out(a10_wr[1587]));
			radix2 #(.width(width)) rd_st9_1588  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1588]), .rdlo_in(a9_wr[1590]),  .coef_in(coef[0]), .rdup_out(a10_wr[1588]), .rdlo_out(a10_wr[1590]));
			radix2 #(.width(width)) rd_st9_1589  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1589]), .rdlo_in(a9_wr[1591]),  .coef_in(coef[512]), .rdup_out(a10_wr[1589]), .rdlo_out(a10_wr[1591]));
			radix2 #(.width(width)) rd_st9_1592  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1592]), .rdlo_in(a9_wr[1594]),  .coef_in(coef[0]), .rdup_out(a10_wr[1592]), .rdlo_out(a10_wr[1594]));
			radix2 #(.width(width)) rd_st9_1593  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1593]), .rdlo_in(a9_wr[1595]),  .coef_in(coef[512]), .rdup_out(a10_wr[1593]), .rdlo_out(a10_wr[1595]));
			radix2 #(.width(width)) rd_st9_1596  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1596]), .rdlo_in(a9_wr[1598]),  .coef_in(coef[0]), .rdup_out(a10_wr[1596]), .rdlo_out(a10_wr[1598]));
			radix2 #(.width(width)) rd_st9_1597  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1597]), .rdlo_in(a9_wr[1599]),  .coef_in(coef[512]), .rdup_out(a10_wr[1597]), .rdlo_out(a10_wr[1599]));
			radix2 #(.width(width)) rd_st9_1600  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1600]), .rdlo_in(a9_wr[1602]),  .coef_in(coef[0]), .rdup_out(a10_wr[1600]), .rdlo_out(a10_wr[1602]));
			radix2 #(.width(width)) rd_st9_1601  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1601]), .rdlo_in(a9_wr[1603]),  .coef_in(coef[512]), .rdup_out(a10_wr[1601]), .rdlo_out(a10_wr[1603]));
			radix2 #(.width(width)) rd_st9_1604  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1604]), .rdlo_in(a9_wr[1606]),  .coef_in(coef[0]), .rdup_out(a10_wr[1604]), .rdlo_out(a10_wr[1606]));
			radix2 #(.width(width)) rd_st9_1605  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1605]), .rdlo_in(a9_wr[1607]),  .coef_in(coef[512]), .rdup_out(a10_wr[1605]), .rdlo_out(a10_wr[1607]));
			radix2 #(.width(width)) rd_st9_1608  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1608]), .rdlo_in(a9_wr[1610]),  .coef_in(coef[0]), .rdup_out(a10_wr[1608]), .rdlo_out(a10_wr[1610]));
			radix2 #(.width(width)) rd_st9_1609  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1609]), .rdlo_in(a9_wr[1611]),  .coef_in(coef[512]), .rdup_out(a10_wr[1609]), .rdlo_out(a10_wr[1611]));
			radix2 #(.width(width)) rd_st9_1612  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1612]), .rdlo_in(a9_wr[1614]),  .coef_in(coef[0]), .rdup_out(a10_wr[1612]), .rdlo_out(a10_wr[1614]));
			radix2 #(.width(width)) rd_st9_1613  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1613]), .rdlo_in(a9_wr[1615]),  .coef_in(coef[512]), .rdup_out(a10_wr[1613]), .rdlo_out(a10_wr[1615]));
			radix2 #(.width(width)) rd_st9_1616  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1616]), .rdlo_in(a9_wr[1618]),  .coef_in(coef[0]), .rdup_out(a10_wr[1616]), .rdlo_out(a10_wr[1618]));
			radix2 #(.width(width)) rd_st9_1617  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1617]), .rdlo_in(a9_wr[1619]),  .coef_in(coef[512]), .rdup_out(a10_wr[1617]), .rdlo_out(a10_wr[1619]));
			radix2 #(.width(width)) rd_st9_1620  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1620]), .rdlo_in(a9_wr[1622]),  .coef_in(coef[0]), .rdup_out(a10_wr[1620]), .rdlo_out(a10_wr[1622]));
			radix2 #(.width(width)) rd_st9_1621  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1621]), .rdlo_in(a9_wr[1623]),  .coef_in(coef[512]), .rdup_out(a10_wr[1621]), .rdlo_out(a10_wr[1623]));
			radix2 #(.width(width)) rd_st9_1624  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1624]), .rdlo_in(a9_wr[1626]),  .coef_in(coef[0]), .rdup_out(a10_wr[1624]), .rdlo_out(a10_wr[1626]));
			radix2 #(.width(width)) rd_st9_1625  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1625]), .rdlo_in(a9_wr[1627]),  .coef_in(coef[512]), .rdup_out(a10_wr[1625]), .rdlo_out(a10_wr[1627]));
			radix2 #(.width(width)) rd_st9_1628  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1628]), .rdlo_in(a9_wr[1630]),  .coef_in(coef[0]), .rdup_out(a10_wr[1628]), .rdlo_out(a10_wr[1630]));
			radix2 #(.width(width)) rd_st9_1629  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1629]), .rdlo_in(a9_wr[1631]),  .coef_in(coef[512]), .rdup_out(a10_wr[1629]), .rdlo_out(a10_wr[1631]));
			radix2 #(.width(width)) rd_st9_1632  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1632]), .rdlo_in(a9_wr[1634]),  .coef_in(coef[0]), .rdup_out(a10_wr[1632]), .rdlo_out(a10_wr[1634]));
			radix2 #(.width(width)) rd_st9_1633  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1633]), .rdlo_in(a9_wr[1635]),  .coef_in(coef[512]), .rdup_out(a10_wr[1633]), .rdlo_out(a10_wr[1635]));
			radix2 #(.width(width)) rd_st9_1636  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1636]), .rdlo_in(a9_wr[1638]),  .coef_in(coef[0]), .rdup_out(a10_wr[1636]), .rdlo_out(a10_wr[1638]));
			radix2 #(.width(width)) rd_st9_1637  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1637]), .rdlo_in(a9_wr[1639]),  .coef_in(coef[512]), .rdup_out(a10_wr[1637]), .rdlo_out(a10_wr[1639]));
			radix2 #(.width(width)) rd_st9_1640  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1640]), .rdlo_in(a9_wr[1642]),  .coef_in(coef[0]), .rdup_out(a10_wr[1640]), .rdlo_out(a10_wr[1642]));
			radix2 #(.width(width)) rd_st9_1641  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1641]), .rdlo_in(a9_wr[1643]),  .coef_in(coef[512]), .rdup_out(a10_wr[1641]), .rdlo_out(a10_wr[1643]));
			radix2 #(.width(width)) rd_st9_1644  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1644]), .rdlo_in(a9_wr[1646]),  .coef_in(coef[0]), .rdup_out(a10_wr[1644]), .rdlo_out(a10_wr[1646]));
			radix2 #(.width(width)) rd_st9_1645  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1645]), .rdlo_in(a9_wr[1647]),  .coef_in(coef[512]), .rdup_out(a10_wr[1645]), .rdlo_out(a10_wr[1647]));
			radix2 #(.width(width)) rd_st9_1648  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1648]), .rdlo_in(a9_wr[1650]),  .coef_in(coef[0]), .rdup_out(a10_wr[1648]), .rdlo_out(a10_wr[1650]));
			radix2 #(.width(width)) rd_st9_1649  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1649]), .rdlo_in(a9_wr[1651]),  .coef_in(coef[512]), .rdup_out(a10_wr[1649]), .rdlo_out(a10_wr[1651]));
			radix2 #(.width(width)) rd_st9_1652  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1652]), .rdlo_in(a9_wr[1654]),  .coef_in(coef[0]), .rdup_out(a10_wr[1652]), .rdlo_out(a10_wr[1654]));
			radix2 #(.width(width)) rd_st9_1653  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1653]), .rdlo_in(a9_wr[1655]),  .coef_in(coef[512]), .rdup_out(a10_wr[1653]), .rdlo_out(a10_wr[1655]));
			radix2 #(.width(width)) rd_st9_1656  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1656]), .rdlo_in(a9_wr[1658]),  .coef_in(coef[0]), .rdup_out(a10_wr[1656]), .rdlo_out(a10_wr[1658]));
			radix2 #(.width(width)) rd_st9_1657  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1657]), .rdlo_in(a9_wr[1659]),  .coef_in(coef[512]), .rdup_out(a10_wr[1657]), .rdlo_out(a10_wr[1659]));
			radix2 #(.width(width)) rd_st9_1660  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1660]), .rdlo_in(a9_wr[1662]),  .coef_in(coef[0]), .rdup_out(a10_wr[1660]), .rdlo_out(a10_wr[1662]));
			radix2 #(.width(width)) rd_st9_1661  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1661]), .rdlo_in(a9_wr[1663]),  .coef_in(coef[512]), .rdup_out(a10_wr[1661]), .rdlo_out(a10_wr[1663]));
			radix2 #(.width(width)) rd_st9_1664  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1664]), .rdlo_in(a9_wr[1666]),  .coef_in(coef[0]), .rdup_out(a10_wr[1664]), .rdlo_out(a10_wr[1666]));
			radix2 #(.width(width)) rd_st9_1665  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1665]), .rdlo_in(a9_wr[1667]),  .coef_in(coef[512]), .rdup_out(a10_wr[1665]), .rdlo_out(a10_wr[1667]));
			radix2 #(.width(width)) rd_st9_1668  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1668]), .rdlo_in(a9_wr[1670]),  .coef_in(coef[0]), .rdup_out(a10_wr[1668]), .rdlo_out(a10_wr[1670]));
			radix2 #(.width(width)) rd_st9_1669  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1669]), .rdlo_in(a9_wr[1671]),  .coef_in(coef[512]), .rdup_out(a10_wr[1669]), .rdlo_out(a10_wr[1671]));
			radix2 #(.width(width)) rd_st9_1672  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1672]), .rdlo_in(a9_wr[1674]),  .coef_in(coef[0]), .rdup_out(a10_wr[1672]), .rdlo_out(a10_wr[1674]));
			radix2 #(.width(width)) rd_st9_1673  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1673]), .rdlo_in(a9_wr[1675]),  .coef_in(coef[512]), .rdup_out(a10_wr[1673]), .rdlo_out(a10_wr[1675]));
			radix2 #(.width(width)) rd_st9_1676  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1676]), .rdlo_in(a9_wr[1678]),  .coef_in(coef[0]), .rdup_out(a10_wr[1676]), .rdlo_out(a10_wr[1678]));
			radix2 #(.width(width)) rd_st9_1677  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1677]), .rdlo_in(a9_wr[1679]),  .coef_in(coef[512]), .rdup_out(a10_wr[1677]), .rdlo_out(a10_wr[1679]));
			radix2 #(.width(width)) rd_st9_1680  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1680]), .rdlo_in(a9_wr[1682]),  .coef_in(coef[0]), .rdup_out(a10_wr[1680]), .rdlo_out(a10_wr[1682]));
			radix2 #(.width(width)) rd_st9_1681  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1681]), .rdlo_in(a9_wr[1683]),  .coef_in(coef[512]), .rdup_out(a10_wr[1681]), .rdlo_out(a10_wr[1683]));
			radix2 #(.width(width)) rd_st9_1684  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1684]), .rdlo_in(a9_wr[1686]),  .coef_in(coef[0]), .rdup_out(a10_wr[1684]), .rdlo_out(a10_wr[1686]));
			radix2 #(.width(width)) rd_st9_1685  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1685]), .rdlo_in(a9_wr[1687]),  .coef_in(coef[512]), .rdup_out(a10_wr[1685]), .rdlo_out(a10_wr[1687]));
			radix2 #(.width(width)) rd_st9_1688  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1688]), .rdlo_in(a9_wr[1690]),  .coef_in(coef[0]), .rdup_out(a10_wr[1688]), .rdlo_out(a10_wr[1690]));
			radix2 #(.width(width)) rd_st9_1689  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1689]), .rdlo_in(a9_wr[1691]),  .coef_in(coef[512]), .rdup_out(a10_wr[1689]), .rdlo_out(a10_wr[1691]));
			radix2 #(.width(width)) rd_st9_1692  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1692]), .rdlo_in(a9_wr[1694]),  .coef_in(coef[0]), .rdup_out(a10_wr[1692]), .rdlo_out(a10_wr[1694]));
			radix2 #(.width(width)) rd_st9_1693  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1693]), .rdlo_in(a9_wr[1695]),  .coef_in(coef[512]), .rdup_out(a10_wr[1693]), .rdlo_out(a10_wr[1695]));
			radix2 #(.width(width)) rd_st9_1696  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1696]), .rdlo_in(a9_wr[1698]),  .coef_in(coef[0]), .rdup_out(a10_wr[1696]), .rdlo_out(a10_wr[1698]));
			radix2 #(.width(width)) rd_st9_1697  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1697]), .rdlo_in(a9_wr[1699]),  .coef_in(coef[512]), .rdup_out(a10_wr[1697]), .rdlo_out(a10_wr[1699]));
			radix2 #(.width(width)) rd_st9_1700  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1700]), .rdlo_in(a9_wr[1702]),  .coef_in(coef[0]), .rdup_out(a10_wr[1700]), .rdlo_out(a10_wr[1702]));
			radix2 #(.width(width)) rd_st9_1701  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1701]), .rdlo_in(a9_wr[1703]),  .coef_in(coef[512]), .rdup_out(a10_wr[1701]), .rdlo_out(a10_wr[1703]));
			radix2 #(.width(width)) rd_st9_1704  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1704]), .rdlo_in(a9_wr[1706]),  .coef_in(coef[0]), .rdup_out(a10_wr[1704]), .rdlo_out(a10_wr[1706]));
			radix2 #(.width(width)) rd_st9_1705  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1705]), .rdlo_in(a9_wr[1707]),  .coef_in(coef[512]), .rdup_out(a10_wr[1705]), .rdlo_out(a10_wr[1707]));
			radix2 #(.width(width)) rd_st9_1708  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1708]), .rdlo_in(a9_wr[1710]),  .coef_in(coef[0]), .rdup_out(a10_wr[1708]), .rdlo_out(a10_wr[1710]));
			radix2 #(.width(width)) rd_st9_1709  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1709]), .rdlo_in(a9_wr[1711]),  .coef_in(coef[512]), .rdup_out(a10_wr[1709]), .rdlo_out(a10_wr[1711]));
			radix2 #(.width(width)) rd_st9_1712  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1712]), .rdlo_in(a9_wr[1714]),  .coef_in(coef[0]), .rdup_out(a10_wr[1712]), .rdlo_out(a10_wr[1714]));
			radix2 #(.width(width)) rd_st9_1713  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1713]), .rdlo_in(a9_wr[1715]),  .coef_in(coef[512]), .rdup_out(a10_wr[1713]), .rdlo_out(a10_wr[1715]));
			radix2 #(.width(width)) rd_st9_1716  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1716]), .rdlo_in(a9_wr[1718]),  .coef_in(coef[0]), .rdup_out(a10_wr[1716]), .rdlo_out(a10_wr[1718]));
			radix2 #(.width(width)) rd_st9_1717  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1717]), .rdlo_in(a9_wr[1719]),  .coef_in(coef[512]), .rdup_out(a10_wr[1717]), .rdlo_out(a10_wr[1719]));
			radix2 #(.width(width)) rd_st9_1720  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1720]), .rdlo_in(a9_wr[1722]),  .coef_in(coef[0]), .rdup_out(a10_wr[1720]), .rdlo_out(a10_wr[1722]));
			radix2 #(.width(width)) rd_st9_1721  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1721]), .rdlo_in(a9_wr[1723]),  .coef_in(coef[512]), .rdup_out(a10_wr[1721]), .rdlo_out(a10_wr[1723]));
			radix2 #(.width(width)) rd_st9_1724  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1724]), .rdlo_in(a9_wr[1726]),  .coef_in(coef[0]), .rdup_out(a10_wr[1724]), .rdlo_out(a10_wr[1726]));
			radix2 #(.width(width)) rd_st9_1725  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1725]), .rdlo_in(a9_wr[1727]),  .coef_in(coef[512]), .rdup_out(a10_wr[1725]), .rdlo_out(a10_wr[1727]));
			radix2 #(.width(width)) rd_st9_1728  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1728]), .rdlo_in(a9_wr[1730]),  .coef_in(coef[0]), .rdup_out(a10_wr[1728]), .rdlo_out(a10_wr[1730]));
			radix2 #(.width(width)) rd_st9_1729  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1729]), .rdlo_in(a9_wr[1731]),  .coef_in(coef[512]), .rdup_out(a10_wr[1729]), .rdlo_out(a10_wr[1731]));
			radix2 #(.width(width)) rd_st9_1732  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1732]), .rdlo_in(a9_wr[1734]),  .coef_in(coef[0]), .rdup_out(a10_wr[1732]), .rdlo_out(a10_wr[1734]));
			radix2 #(.width(width)) rd_st9_1733  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1733]), .rdlo_in(a9_wr[1735]),  .coef_in(coef[512]), .rdup_out(a10_wr[1733]), .rdlo_out(a10_wr[1735]));
			radix2 #(.width(width)) rd_st9_1736  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1736]), .rdlo_in(a9_wr[1738]),  .coef_in(coef[0]), .rdup_out(a10_wr[1736]), .rdlo_out(a10_wr[1738]));
			radix2 #(.width(width)) rd_st9_1737  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1737]), .rdlo_in(a9_wr[1739]),  .coef_in(coef[512]), .rdup_out(a10_wr[1737]), .rdlo_out(a10_wr[1739]));
			radix2 #(.width(width)) rd_st9_1740  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1740]), .rdlo_in(a9_wr[1742]),  .coef_in(coef[0]), .rdup_out(a10_wr[1740]), .rdlo_out(a10_wr[1742]));
			radix2 #(.width(width)) rd_st9_1741  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1741]), .rdlo_in(a9_wr[1743]),  .coef_in(coef[512]), .rdup_out(a10_wr[1741]), .rdlo_out(a10_wr[1743]));
			radix2 #(.width(width)) rd_st9_1744  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1744]), .rdlo_in(a9_wr[1746]),  .coef_in(coef[0]), .rdup_out(a10_wr[1744]), .rdlo_out(a10_wr[1746]));
			radix2 #(.width(width)) rd_st9_1745  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1745]), .rdlo_in(a9_wr[1747]),  .coef_in(coef[512]), .rdup_out(a10_wr[1745]), .rdlo_out(a10_wr[1747]));
			radix2 #(.width(width)) rd_st9_1748  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1748]), .rdlo_in(a9_wr[1750]),  .coef_in(coef[0]), .rdup_out(a10_wr[1748]), .rdlo_out(a10_wr[1750]));
			radix2 #(.width(width)) rd_st9_1749  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1749]), .rdlo_in(a9_wr[1751]),  .coef_in(coef[512]), .rdup_out(a10_wr[1749]), .rdlo_out(a10_wr[1751]));
			radix2 #(.width(width)) rd_st9_1752  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1752]), .rdlo_in(a9_wr[1754]),  .coef_in(coef[0]), .rdup_out(a10_wr[1752]), .rdlo_out(a10_wr[1754]));
			radix2 #(.width(width)) rd_st9_1753  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1753]), .rdlo_in(a9_wr[1755]),  .coef_in(coef[512]), .rdup_out(a10_wr[1753]), .rdlo_out(a10_wr[1755]));
			radix2 #(.width(width)) rd_st9_1756  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1756]), .rdlo_in(a9_wr[1758]),  .coef_in(coef[0]), .rdup_out(a10_wr[1756]), .rdlo_out(a10_wr[1758]));
			radix2 #(.width(width)) rd_st9_1757  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1757]), .rdlo_in(a9_wr[1759]),  .coef_in(coef[512]), .rdup_out(a10_wr[1757]), .rdlo_out(a10_wr[1759]));
			radix2 #(.width(width)) rd_st9_1760  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1760]), .rdlo_in(a9_wr[1762]),  .coef_in(coef[0]), .rdup_out(a10_wr[1760]), .rdlo_out(a10_wr[1762]));
			radix2 #(.width(width)) rd_st9_1761  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1761]), .rdlo_in(a9_wr[1763]),  .coef_in(coef[512]), .rdup_out(a10_wr[1761]), .rdlo_out(a10_wr[1763]));
			radix2 #(.width(width)) rd_st9_1764  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1764]), .rdlo_in(a9_wr[1766]),  .coef_in(coef[0]), .rdup_out(a10_wr[1764]), .rdlo_out(a10_wr[1766]));
			radix2 #(.width(width)) rd_st9_1765  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1765]), .rdlo_in(a9_wr[1767]),  .coef_in(coef[512]), .rdup_out(a10_wr[1765]), .rdlo_out(a10_wr[1767]));
			radix2 #(.width(width)) rd_st9_1768  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1768]), .rdlo_in(a9_wr[1770]),  .coef_in(coef[0]), .rdup_out(a10_wr[1768]), .rdlo_out(a10_wr[1770]));
			radix2 #(.width(width)) rd_st9_1769  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1769]), .rdlo_in(a9_wr[1771]),  .coef_in(coef[512]), .rdup_out(a10_wr[1769]), .rdlo_out(a10_wr[1771]));
			radix2 #(.width(width)) rd_st9_1772  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1772]), .rdlo_in(a9_wr[1774]),  .coef_in(coef[0]), .rdup_out(a10_wr[1772]), .rdlo_out(a10_wr[1774]));
			radix2 #(.width(width)) rd_st9_1773  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1773]), .rdlo_in(a9_wr[1775]),  .coef_in(coef[512]), .rdup_out(a10_wr[1773]), .rdlo_out(a10_wr[1775]));
			radix2 #(.width(width)) rd_st9_1776  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1776]), .rdlo_in(a9_wr[1778]),  .coef_in(coef[0]), .rdup_out(a10_wr[1776]), .rdlo_out(a10_wr[1778]));
			radix2 #(.width(width)) rd_st9_1777  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1777]), .rdlo_in(a9_wr[1779]),  .coef_in(coef[512]), .rdup_out(a10_wr[1777]), .rdlo_out(a10_wr[1779]));
			radix2 #(.width(width)) rd_st9_1780  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1780]), .rdlo_in(a9_wr[1782]),  .coef_in(coef[0]), .rdup_out(a10_wr[1780]), .rdlo_out(a10_wr[1782]));
			radix2 #(.width(width)) rd_st9_1781  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1781]), .rdlo_in(a9_wr[1783]),  .coef_in(coef[512]), .rdup_out(a10_wr[1781]), .rdlo_out(a10_wr[1783]));
			radix2 #(.width(width)) rd_st9_1784  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1784]), .rdlo_in(a9_wr[1786]),  .coef_in(coef[0]), .rdup_out(a10_wr[1784]), .rdlo_out(a10_wr[1786]));
			radix2 #(.width(width)) rd_st9_1785  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1785]), .rdlo_in(a9_wr[1787]),  .coef_in(coef[512]), .rdup_out(a10_wr[1785]), .rdlo_out(a10_wr[1787]));
			radix2 #(.width(width)) rd_st9_1788  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1788]), .rdlo_in(a9_wr[1790]),  .coef_in(coef[0]), .rdup_out(a10_wr[1788]), .rdlo_out(a10_wr[1790]));
			radix2 #(.width(width)) rd_st9_1789  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1789]), .rdlo_in(a9_wr[1791]),  .coef_in(coef[512]), .rdup_out(a10_wr[1789]), .rdlo_out(a10_wr[1791]));
			radix2 #(.width(width)) rd_st9_1792  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1792]), .rdlo_in(a9_wr[1794]),  .coef_in(coef[0]), .rdup_out(a10_wr[1792]), .rdlo_out(a10_wr[1794]));
			radix2 #(.width(width)) rd_st9_1793  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1793]), .rdlo_in(a9_wr[1795]),  .coef_in(coef[512]), .rdup_out(a10_wr[1793]), .rdlo_out(a10_wr[1795]));
			radix2 #(.width(width)) rd_st9_1796  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1796]), .rdlo_in(a9_wr[1798]),  .coef_in(coef[0]), .rdup_out(a10_wr[1796]), .rdlo_out(a10_wr[1798]));
			radix2 #(.width(width)) rd_st9_1797  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1797]), .rdlo_in(a9_wr[1799]),  .coef_in(coef[512]), .rdup_out(a10_wr[1797]), .rdlo_out(a10_wr[1799]));
			radix2 #(.width(width)) rd_st9_1800  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1800]), .rdlo_in(a9_wr[1802]),  .coef_in(coef[0]), .rdup_out(a10_wr[1800]), .rdlo_out(a10_wr[1802]));
			radix2 #(.width(width)) rd_st9_1801  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1801]), .rdlo_in(a9_wr[1803]),  .coef_in(coef[512]), .rdup_out(a10_wr[1801]), .rdlo_out(a10_wr[1803]));
			radix2 #(.width(width)) rd_st9_1804  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1804]), .rdlo_in(a9_wr[1806]),  .coef_in(coef[0]), .rdup_out(a10_wr[1804]), .rdlo_out(a10_wr[1806]));
			radix2 #(.width(width)) rd_st9_1805  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1805]), .rdlo_in(a9_wr[1807]),  .coef_in(coef[512]), .rdup_out(a10_wr[1805]), .rdlo_out(a10_wr[1807]));
			radix2 #(.width(width)) rd_st9_1808  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1808]), .rdlo_in(a9_wr[1810]),  .coef_in(coef[0]), .rdup_out(a10_wr[1808]), .rdlo_out(a10_wr[1810]));
			radix2 #(.width(width)) rd_st9_1809  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1809]), .rdlo_in(a9_wr[1811]),  .coef_in(coef[512]), .rdup_out(a10_wr[1809]), .rdlo_out(a10_wr[1811]));
			radix2 #(.width(width)) rd_st9_1812  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1812]), .rdlo_in(a9_wr[1814]),  .coef_in(coef[0]), .rdup_out(a10_wr[1812]), .rdlo_out(a10_wr[1814]));
			radix2 #(.width(width)) rd_st9_1813  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1813]), .rdlo_in(a9_wr[1815]),  .coef_in(coef[512]), .rdup_out(a10_wr[1813]), .rdlo_out(a10_wr[1815]));
			radix2 #(.width(width)) rd_st9_1816  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1816]), .rdlo_in(a9_wr[1818]),  .coef_in(coef[0]), .rdup_out(a10_wr[1816]), .rdlo_out(a10_wr[1818]));
			radix2 #(.width(width)) rd_st9_1817  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1817]), .rdlo_in(a9_wr[1819]),  .coef_in(coef[512]), .rdup_out(a10_wr[1817]), .rdlo_out(a10_wr[1819]));
			radix2 #(.width(width)) rd_st9_1820  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1820]), .rdlo_in(a9_wr[1822]),  .coef_in(coef[0]), .rdup_out(a10_wr[1820]), .rdlo_out(a10_wr[1822]));
			radix2 #(.width(width)) rd_st9_1821  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1821]), .rdlo_in(a9_wr[1823]),  .coef_in(coef[512]), .rdup_out(a10_wr[1821]), .rdlo_out(a10_wr[1823]));
			radix2 #(.width(width)) rd_st9_1824  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1824]), .rdlo_in(a9_wr[1826]),  .coef_in(coef[0]), .rdup_out(a10_wr[1824]), .rdlo_out(a10_wr[1826]));
			radix2 #(.width(width)) rd_st9_1825  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1825]), .rdlo_in(a9_wr[1827]),  .coef_in(coef[512]), .rdup_out(a10_wr[1825]), .rdlo_out(a10_wr[1827]));
			radix2 #(.width(width)) rd_st9_1828  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1828]), .rdlo_in(a9_wr[1830]),  .coef_in(coef[0]), .rdup_out(a10_wr[1828]), .rdlo_out(a10_wr[1830]));
			radix2 #(.width(width)) rd_st9_1829  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1829]), .rdlo_in(a9_wr[1831]),  .coef_in(coef[512]), .rdup_out(a10_wr[1829]), .rdlo_out(a10_wr[1831]));
			radix2 #(.width(width)) rd_st9_1832  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1832]), .rdlo_in(a9_wr[1834]),  .coef_in(coef[0]), .rdup_out(a10_wr[1832]), .rdlo_out(a10_wr[1834]));
			radix2 #(.width(width)) rd_st9_1833  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1833]), .rdlo_in(a9_wr[1835]),  .coef_in(coef[512]), .rdup_out(a10_wr[1833]), .rdlo_out(a10_wr[1835]));
			radix2 #(.width(width)) rd_st9_1836  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1836]), .rdlo_in(a9_wr[1838]),  .coef_in(coef[0]), .rdup_out(a10_wr[1836]), .rdlo_out(a10_wr[1838]));
			radix2 #(.width(width)) rd_st9_1837  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1837]), .rdlo_in(a9_wr[1839]),  .coef_in(coef[512]), .rdup_out(a10_wr[1837]), .rdlo_out(a10_wr[1839]));
			radix2 #(.width(width)) rd_st9_1840  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1840]), .rdlo_in(a9_wr[1842]),  .coef_in(coef[0]), .rdup_out(a10_wr[1840]), .rdlo_out(a10_wr[1842]));
			radix2 #(.width(width)) rd_st9_1841  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1841]), .rdlo_in(a9_wr[1843]),  .coef_in(coef[512]), .rdup_out(a10_wr[1841]), .rdlo_out(a10_wr[1843]));
			radix2 #(.width(width)) rd_st9_1844  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1844]), .rdlo_in(a9_wr[1846]),  .coef_in(coef[0]), .rdup_out(a10_wr[1844]), .rdlo_out(a10_wr[1846]));
			radix2 #(.width(width)) rd_st9_1845  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1845]), .rdlo_in(a9_wr[1847]),  .coef_in(coef[512]), .rdup_out(a10_wr[1845]), .rdlo_out(a10_wr[1847]));
			radix2 #(.width(width)) rd_st9_1848  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1848]), .rdlo_in(a9_wr[1850]),  .coef_in(coef[0]), .rdup_out(a10_wr[1848]), .rdlo_out(a10_wr[1850]));
			radix2 #(.width(width)) rd_st9_1849  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1849]), .rdlo_in(a9_wr[1851]),  .coef_in(coef[512]), .rdup_out(a10_wr[1849]), .rdlo_out(a10_wr[1851]));
			radix2 #(.width(width)) rd_st9_1852  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1852]), .rdlo_in(a9_wr[1854]),  .coef_in(coef[0]), .rdup_out(a10_wr[1852]), .rdlo_out(a10_wr[1854]));
			radix2 #(.width(width)) rd_st9_1853  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1853]), .rdlo_in(a9_wr[1855]),  .coef_in(coef[512]), .rdup_out(a10_wr[1853]), .rdlo_out(a10_wr[1855]));
			radix2 #(.width(width)) rd_st9_1856  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1856]), .rdlo_in(a9_wr[1858]),  .coef_in(coef[0]), .rdup_out(a10_wr[1856]), .rdlo_out(a10_wr[1858]));
			radix2 #(.width(width)) rd_st9_1857  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1857]), .rdlo_in(a9_wr[1859]),  .coef_in(coef[512]), .rdup_out(a10_wr[1857]), .rdlo_out(a10_wr[1859]));
			radix2 #(.width(width)) rd_st9_1860  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1860]), .rdlo_in(a9_wr[1862]),  .coef_in(coef[0]), .rdup_out(a10_wr[1860]), .rdlo_out(a10_wr[1862]));
			radix2 #(.width(width)) rd_st9_1861  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1861]), .rdlo_in(a9_wr[1863]),  .coef_in(coef[512]), .rdup_out(a10_wr[1861]), .rdlo_out(a10_wr[1863]));
			radix2 #(.width(width)) rd_st9_1864  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1864]), .rdlo_in(a9_wr[1866]),  .coef_in(coef[0]), .rdup_out(a10_wr[1864]), .rdlo_out(a10_wr[1866]));
			radix2 #(.width(width)) rd_st9_1865  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1865]), .rdlo_in(a9_wr[1867]),  .coef_in(coef[512]), .rdup_out(a10_wr[1865]), .rdlo_out(a10_wr[1867]));
			radix2 #(.width(width)) rd_st9_1868  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1868]), .rdlo_in(a9_wr[1870]),  .coef_in(coef[0]), .rdup_out(a10_wr[1868]), .rdlo_out(a10_wr[1870]));
			radix2 #(.width(width)) rd_st9_1869  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1869]), .rdlo_in(a9_wr[1871]),  .coef_in(coef[512]), .rdup_out(a10_wr[1869]), .rdlo_out(a10_wr[1871]));
			radix2 #(.width(width)) rd_st9_1872  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1872]), .rdlo_in(a9_wr[1874]),  .coef_in(coef[0]), .rdup_out(a10_wr[1872]), .rdlo_out(a10_wr[1874]));
			radix2 #(.width(width)) rd_st9_1873  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1873]), .rdlo_in(a9_wr[1875]),  .coef_in(coef[512]), .rdup_out(a10_wr[1873]), .rdlo_out(a10_wr[1875]));
			radix2 #(.width(width)) rd_st9_1876  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1876]), .rdlo_in(a9_wr[1878]),  .coef_in(coef[0]), .rdup_out(a10_wr[1876]), .rdlo_out(a10_wr[1878]));
			radix2 #(.width(width)) rd_st9_1877  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1877]), .rdlo_in(a9_wr[1879]),  .coef_in(coef[512]), .rdup_out(a10_wr[1877]), .rdlo_out(a10_wr[1879]));
			radix2 #(.width(width)) rd_st9_1880  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1880]), .rdlo_in(a9_wr[1882]),  .coef_in(coef[0]), .rdup_out(a10_wr[1880]), .rdlo_out(a10_wr[1882]));
			radix2 #(.width(width)) rd_st9_1881  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1881]), .rdlo_in(a9_wr[1883]),  .coef_in(coef[512]), .rdup_out(a10_wr[1881]), .rdlo_out(a10_wr[1883]));
			radix2 #(.width(width)) rd_st9_1884  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1884]), .rdlo_in(a9_wr[1886]),  .coef_in(coef[0]), .rdup_out(a10_wr[1884]), .rdlo_out(a10_wr[1886]));
			radix2 #(.width(width)) rd_st9_1885  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1885]), .rdlo_in(a9_wr[1887]),  .coef_in(coef[512]), .rdup_out(a10_wr[1885]), .rdlo_out(a10_wr[1887]));
			radix2 #(.width(width)) rd_st9_1888  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1888]), .rdlo_in(a9_wr[1890]),  .coef_in(coef[0]), .rdup_out(a10_wr[1888]), .rdlo_out(a10_wr[1890]));
			radix2 #(.width(width)) rd_st9_1889  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1889]), .rdlo_in(a9_wr[1891]),  .coef_in(coef[512]), .rdup_out(a10_wr[1889]), .rdlo_out(a10_wr[1891]));
			radix2 #(.width(width)) rd_st9_1892  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1892]), .rdlo_in(a9_wr[1894]),  .coef_in(coef[0]), .rdup_out(a10_wr[1892]), .rdlo_out(a10_wr[1894]));
			radix2 #(.width(width)) rd_st9_1893  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1893]), .rdlo_in(a9_wr[1895]),  .coef_in(coef[512]), .rdup_out(a10_wr[1893]), .rdlo_out(a10_wr[1895]));
			radix2 #(.width(width)) rd_st9_1896  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1896]), .rdlo_in(a9_wr[1898]),  .coef_in(coef[0]), .rdup_out(a10_wr[1896]), .rdlo_out(a10_wr[1898]));
			radix2 #(.width(width)) rd_st9_1897  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1897]), .rdlo_in(a9_wr[1899]),  .coef_in(coef[512]), .rdup_out(a10_wr[1897]), .rdlo_out(a10_wr[1899]));
			radix2 #(.width(width)) rd_st9_1900  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1900]), .rdlo_in(a9_wr[1902]),  .coef_in(coef[0]), .rdup_out(a10_wr[1900]), .rdlo_out(a10_wr[1902]));
			radix2 #(.width(width)) rd_st9_1901  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1901]), .rdlo_in(a9_wr[1903]),  .coef_in(coef[512]), .rdup_out(a10_wr[1901]), .rdlo_out(a10_wr[1903]));
			radix2 #(.width(width)) rd_st9_1904  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1904]), .rdlo_in(a9_wr[1906]),  .coef_in(coef[0]), .rdup_out(a10_wr[1904]), .rdlo_out(a10_wr[1906]));
			radix2 #(.width(width)) rd_st9_1905  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1905]), .rdlo_in(a9_wr[1907]),  .coef_in(coef[512]), .rdup_out(a10_wr[1905]), .rdlo_out(a10_wr[1907]));
			radix2 #(.width(width)) rd_st9_1908  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1908]), .rdlo_in(a9_wr[1910]),  .coef_in(coef[0]), .rdup_out(a10_wr[1908]), .rdlo_out(a10_wr[1910]));
			radix2 #(.width(width)) rd_st9_1909  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1909]), .rdlo_in(a9_wr[1911]),  .coef_in(coef[512]), .rdup_out(a10_wr[1909]), .rdlo_out(a10_wr[1911]));
			radix2 #(.width(width)) rd_st9_1912  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1912]), .rdlo_in(a9_wr[1914]),  .coef_in(coef[0]), .rdup_out(a10_wr[1912]), .rdlo_out(a10_wr[1914]));
			radix2 #(.width(width)) rd_st9_1913  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1913]), .rdlo_in(a9_wr[1915]),  .coef_in(coef[512]), .rdup_out(a10_wr[1913]), .rdlo_out(a10_wr[1915]));
			radix2 #(.width(width)) rd_st9_1916  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1916]), .rdlo_in(a9_wr[1918]),  .coef_in(coef[0]), .rdup_out(a10_wr[1916]), .rdlo_out(a10_wr[1918]));
			radix2 #(.width(width)) rd_st9_1917  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1917]), .rdlo_in(a9_wr[1919]),  .coef_in(coef[512]), .rdup_out(a10_wr[1917]), .rdlo_out(a10_wr[1919]));
			radix2 #(.width(width)) rd_st9_1920  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1920]), .rdlo_in(a9_wr[1922]),  .coef_in(coef[0]), .rdup_out(a10_wr[1920]), .rdlo_out(a10_wr[1922]));
			radix2 #(.width(width)) rd_st9_1921  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1921]), .rdlo_in(a9_wr[1923]),  .coef_in(coef[512]), .rdup_out(a10_wr[1921]), .rdlo_out(a10_wr[1923]));
			radix2 #(.width(width)) rd_st9_1924  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1924]), .rdlo_in(a9_wr[1926]),  .coef_in(coef[0]), .rdup_out(a10_wr[1924]), .rdlo_out(a10_wr[1926]));
			radix2 #(.width(width)) rd_st9_1925  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1925]), .rdlo_in(a9_wr[1927]),  .coef_in(coef[512]), .rdup_out(a10_wr[1925]), .rdlo_out(a10_wr[1927]));
			radix2 #(.width(width)) rd_st9_1928  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1928]), .rdlo_in(a9_wr[1930]),  .coef_in(coef[0]), .rdup_out(a10_wr[1928]), .rdlo_out(a10_wr[1930]));
			radix2 #(.width(width)) rd_st9_1929  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1929]), .rdlo_in(a9_wr[1931]),  .coef_in(coef[512]), .rdup_out(a10_wr[1929]), .rdlo_out(a10_wr[1931]));
			radix2 #(.width(width)) rd_st9_1932  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1932]), .rdlo_in(a9_wr[1934]),  .coef_in(coef[0]), .rdup_out(a10_wr[1932]), .rdlo_out(a10_wr[1934]));
			radix2 #(.width(width)) rd_st9_1933  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1933]), .rdlo_in(a9_wr[1935]),  .coef_in(coef[512]), .rdup_out(a10_wr[1933]), .rdlo_out(a10_wr[1935]));
			radix2 #(.width(width)) rd_st9_1936  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1936]), .rdlo_in(a9_wr[1938]),  .coef_in(coef[0]), .rdup_out(a10_wr[1936]), .rdlo_out(a10_wr[1938]));
			radix2 #(.width(width)) rd_st9_1937  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1937]), .rdlo_in(a9_wr[1939]),  .coef_in(coef[512]), .rdup_out(a10_wr[1937]), .rdlo_out(a10_wr[1939]));
			radix2 #(.width(width)) rd_st9_1940  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1940]), .rdlo_in(a9_wr[1942]),  .coef_in(coef[0]), .rdup_out(a10_wr[1940]), .rdlo_out(a10_wr[1942]));
			radix2 #(.width(width)) rd_st9_1941  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1941]), .rdlo_in(a9_wr[1943]),  .coef_in(coef[512]), .rdup_out(a10_wr[1941]), .rdlo_out(a10_wr[1943]));
			radix2 #(.width(width)) rd_st9_1944  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1944]), .rdlo_in(a9_wr[1946]),  .coef_in(coef[0]), .rdup_out(a10_wr[1944]), .rdlo_out(a10_wr[1946]));
			radix2 #(.width(width)) rd_st9_1945  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1945]), .rdlo_in(a9_wr[1947]),  .coef_in(coef[512]), .rdup_out(a10_wr[1945]), .rdlo_out(a10_wr[1947]));
			radix2 #(.width(width)) rd_st9_1948  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1948]), .rdlo_in(a9_wr[1950]),  .coef_in(coef[0]), .rdup_out(a10_wr[1948]), .rdlo_out(a10_wr[1950]));
			radix2 #(.width(width)) rd_st9_1949  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1949]), .rdlo_in(a9_wr[1951]),  .coef_in(coef[512]), .rdup_out(a10_wr[1949]), .rdlo_out(a10_wr[1951]));
			radix2 #(.width(width)) rd_st9_1952  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1952]), .rdlo_in(a9_wr[1954]),  .coef_in(coef[0]), .rdup_out(a10_wr[1952]), .rdlo_out(a10_wr[1954]));
			radix2 #(.width(width)) rd_st9_1953  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1953]), .rdlo_in(a9_wr[1955]),  .coef_in(coef[512]), .rdup_out(a10_wr[1953]), .rdlo_out(a10_wr[1955]));
			radix2 #(.width(width)) rd_st9_1956  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1956]), .rdlo_in(a9_wr[1958]),  .coef_in(coef[0]), .rdup_out(a10_wr[1956]), .rdlo_out(a10_wr[1958]));
			radix2 #(.width(width)) rd_st9_1957  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1957]), .rdlo_in(a9_wr[1959]),  .coef_in(coef[512]), .rdup_out(a10_wr[1957]), .rdlo_out(a10_wr[1959]));
			radix2 #(.width(width)) rd_st9_1960  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1960]), .rdlo_in(a9_wr[1962]),  .coef_in(coef[0]), .rdup_out(a10_wr[1960]), .rdlo_out(a10_wr[1962]));
			radix2 #(.width(width)) rd_st9_1961  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1961]), .rdlo_in(a9_wr[1963]),  .coef_in(coef[512]), .rdup_out(a10_wr[1961]), .rdlo_out(a10_wr[1963]));
			radix2 #(.width(width)) rd_st9_1964  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1964]), .rdlo_in(a9_wr[1966]),  .coef_in(coef[0]), .rdup_out(a10_wr[1964]), .rdlo_out(a10_wr[1966]));
			radix2 #(.width(width)) rd_st9_1965  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1965]), .rdlo_in(a9_wr[1967]),  .coef_in(coef[512]), .rdup_out(a10_wr[1965]), .rdlo_out(a10_wr[1967]));
			radix2 #(.width(width)) rd_st9_1968  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1968]), .rdlo_in(a9_wr[1970]),  .coef_in(coef[0]), .rdup_out(a10_wr[1968]), .rdlo_out(a10_wr[1970]));
			radix2 #(.width(width)) rd_st9_1969  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1969]), .rdlo_in(a9_wr[1971]),  .coef_in(coef[512]), .rdup_out(a10_wr[1969]), .rdlo_out(a10_wr[1971]));
			radix2 #(.width(width)) rd_st9_1972  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1972]), .rdlo_in(a9_wr[1974]),  .coef_in(coef[0]), .rdup_out(a10_wr[1972]), .rdlo_out(a10_wr[1974]));
			radix2 #(.width(width)) rd_st9_1973  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1973]), .rdlo_in(a9_wr[1975]),  .coef_in(coef[512]), .rdup_out(a10_wr[1973]), .rdlo_out(a10_wr[1975]));
			radix2 #(.width(width)) rd_st9_1976  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1976]), .rdlo_in(a9_wr[1978]),  .coef_in(coef[0]), .rdup_out(a10_wr[1976]), .rdlo_out(a10_wr[1978]));
			radix2 #(.width(width)) rd_st9_1977  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1977]), .rdlo_in(a9_wr[1979]),  .coef_in(coef[512]), .rdup_out(a10_wr[1977]), .rdlo_out(a10_wr[1979]));
			radix2 #(.width(width)) rd_st9_1980  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1980]), .rdlo_in(a9_wr[1982]),  .coef_in(coef[0]), .rdup_out(a10_wr[1980]), .rdlo_out(a10_wr[1982]));
			radix2 #(.width(width)) rd_st9_1981  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1981]), .rdlo_in(a9_wr[1983]),  .coef_in(coef[512]), .rdup_out(a10_wr[1981]), .rdlo_out(a10_wr[1983]));
			radix2 #(.width(width)) rd_st9_1984  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1984]), .rdlo_in(a9_wr[1986]),  .coef_in(coef[0]), .rdup_out(a10_wr[1984]), .rdlo_out(a10_wr[1986]));
			radix2 #(.width(width)) rd_st9_1985  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1985]), .rdlo_in(a9_wr[1987]),  .coef_in(coef[512]), .rdup_out(a10_wr[1985]), .rdlo_out(a10_wr[1987]));
			radix2 #(.width(width)) rd_st9_1988  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1988]), .rdlo_in(a9_wr[1990]),  .coef_in(coef[0]), .rdup_out(a10_wr[1988]), .rdlo_out(a10_wr[1990]));
			radix2 #(.width(width)) rd_st9_1989  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1989]), .rdlo_in(a9_wr[1991]),  .coef_in(coef[512]), .rdup_out(a10_wr[1989]), .rdlo_out(a10_wr[1991]));
			radix2 #(.width(width)) rd_st9_1992  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1992]), .rdlo_in(a9_wr[1994]),  .coef_in(coef[0]), .rdup_out(a10_wr[1992]), .rdlo_out(a10_wr[1994]));
			radix2 #(.width(width)) rd_st9_1993  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1993]), .rdlo_in(a9_wr[1995]),  .coef_in(coef[512]), .rdup_out(a10_wr[1993]), .rdlo_out(a10_wr[1995]));
			radix2 #(.width(width)) rd_st9_1996  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1996]), .rdlo_in(a9_wr[1998]),  .coef_in(coef[0]), .rdup_out(a10_wr[1996]), .rdlo_out(a10_wr[1998]));
			radix2 #(.width(width)) rd_st9_1997  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[1997]), .rdlo_in(a9_wr[1999]),  .coef_in(coef[512]), .rdup_out(a10_wr[1997]), .rdlo_out(a10_wr[1999]));
			radix2 #(.width(width)) rd_st9_2000  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[2000]), .rdlo_in(a9_wr[2002]),  .coef_in(coef[0]), .rdup_out(a10_wr[2000]), .rdlo_out(a10_wr[2002]));
			radix2 #(.width(width)) rd_st9_2001  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[2001]), .rdlo_in(a9_wr[2003]),  .coef_in(coef[512]), .rdup_out(a10_wr[2001]), .rdlo_out(a10_wr[2003]));
			radix2 #(.width(width)) rd_st9_2004  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[2004]), .rdlo_in(a9_wr[2006]),  .coef_in(coef[0]), .rdup_out(a10_wr[2004]), .rdlo_out(a10_wr[2006]));
			radix2 #(.width(width)) rd_st9_2005  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[2005]), .rdlo_in(a9_wr[2007]),  .coef_in(coef[512]), .rdup_out(a10_wr[2005]), .rdlo_out(a10_wr[2007]));
			radix2 #(.width(width)) rd_st9_2008  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[2008]), .rdlo_in(a9_wr[2010]),  .coef_in(coef[0]), .rdup_out(a10_wr[2008]), .rdlo_out(a10_wr[2010]));
			radix2 #(.width(width)) rd_st9_2009  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[2009]), .rdlo_in(a9_wr[2011]),  .coef_in(coef[512]), .rdup_out(a10_wr[2009]), .rdlo_out(a10_wr[2011]));
			radix2 #(.width(width)) rd_st9_2012  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[2012]), .rdlo_in(a9_wr[2014]),  .coef_in(coef[0]), .rdup_out(a10_wr[2012]), .rdlo_out(a10_wr[2014]));
			radix2 #(.width(width)) rd_st9_2013  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[2013]), .rdlo_in(a9_wr[2015]),  .coef_in(coef[512]), .rdup_out(a10_wr[2013]), .rdlo_out(a10_wr[2015]));
			radix2 #(.width(width)) rd_st9_2016  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[2016]), .rdlo_in(a9_wr[2018]),  .coef_in(coef[0]), .rdup_out(a10_wr[2016]), .rdlo_out(a10_wr[2018]));
			radix2 #(.width(width)) rd_st9_2017  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[2017]), .rdlo_in(a9_wr[2019]),  .coef_in(coef[512]), .rdup_out(a10_wr[2017]), .rdlo_out(a10_wr[2019]));
			radix2 #(.width(width)) rd_st9_2020  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[2020]), .rdlo_in(a9_wr[2022]),  .coef_in(coef[0]), .rdup_out(a10_wr[2020]), .rdlo_out(a10_wr[2022]));
			radix2 #(.width(width)) rd_st9_2021  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[2021]), .rdlo_in(a9_wr[2023]),  .coef_in(coef[512]), .rdup_out(a10_wr[2021]), .rdlo_out(a10_wr[2023]));
			radix2 #(.width(width)) rd_st9_2024  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[2024]), .rdlo_in(a9_wr[2026]),  .coef_in(coef[0]), .rdup_out(a10_wr[2024]), .rdlo_out(a10_wr[2026]));
			radix2 #(.width(width)) rd_st9_2025  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[2025]), .rdlo_in(a9_wr[2027]),  .coef_in(coef[512]), .rdup_out(a10_wr[2025]), .rdlo_out(a10_wr[2027]));
			radix2 #(.width(width)) rd_st9_2028  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[2028]), .rdlo_in(a9_wr[2030]),  .coef_in(coef[0]), .rdup_out(a10_wr[2028]), .rdlo_out(a10_wr[2030]));
			radix2 #(.width(width)) rd_st9_2029  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[2029]), .rdlo_in(a9_wr[2031]),  .coef_in(coef[512]), .rdup_out(a10_wr[2029]), .rdlo_out(a10_wr[2031]));
			radix2 #(.width(width)) rd_st9_2032  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[2032]), .rdlo_in(a9_wr[2034]),  .coef_in(coef[0]), .rdup_out(a10_wr[2032]), .rdlo_out(a10_wr[2034]));
			radix2 #(.width(width)) rd_st9_2033  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[2033]), .rdlo_in(a9_wr[2035]),  .coef_in(coef[512]), .rdup_out(a10_wr[2033]), .rdlo_out(a10_wr[2035]));
			radix2 #(.width(width)) rd_st9_2036  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[2036]), .rdlo_in(a9_wr[2038]),  .coef_in(coef[0]), .rdup_out(a10_wr[2036]), .rdlo_out(a10_wr[2038]));
			radix2 #(.width(width)) rd_st9_2037  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[2037]), .rdlo_in(a9_wr[2039]),  .coef_in(coef[512]), .rdup_out(a10_wr[2037]), .rdlo_out(a10_wr[2039]));
			radix2 #(.width(width)) rd_st9_2040  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[2040]), .rdlo_in(a9_wr[2042]),  .coef_in(coef[0]), .rdup_out(a10_wr[2040]), .rdlo_out(a10_wr[2042]));
			radix2 #(.width(width)) rd_st9_2041  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[2041]), .rdlo_in(a9_wr[2043]),  .coef_in(coef[512]), .rdup_out(a10_wr[2041]), .rdlo_out(a10_wr[2043]));
			radix2 #(.width(width)) rd_st9_2044  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[2044]), .rdlo_in(a9_wr[2046]),  .coef_in(coef[0]), .rdup_out(a10_wr[2044]), .rdlo_out(a10_wr[2046]));
			radix2 #(.width(width)) rd_st9_2045  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a9_wr[2045]), .rdlo_in(a9_wr[2047]),  .coef_in(coef[512]), .rdup_out(a10_wr[2045]), .rdlo_out(a10_wr[2047]));

		//--- radix stage 10
			radix2 #(.width(width)) rd_st10_0  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[0]), .rdlo_in(a10_wr[1]),  .coef_in(coef[0]), .rdup_out(a11_wr[0]), .rdlo_out(a11_wr[1]));
			radix2 #(.width(width)) rd_st10_2  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[2]), .rdlo_in(a10_wr[3]),  .coef_in(coef[0]), .rdup_out(a11_wr[2]), .rdlo_out(a11_wr[3]));
			radix2 #(.width(width)) rd_st10_4  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[4]), .rdlo_in(a10_wr[5]),  .coef_in(coef[0]), .rdup_out(a11_wr[4]), .rdlo_out(a11_wr[5]));
			radix2 #(.width(width)) rd_st10_6  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[6]), .rdlo_in(a10_wr[7]),  .coef_in(coef[0]), .rdup_out(a11_wr[6]), .rdlo_out(a11_wr[7]));
			radix2 #(.width(width)) rd_st10_8  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[8]), .rdlo_in(a10_wr[9]),  .coef_in(coef[0]), .rdup_out(a11_wr[8]), .rdlo_out(a11_wr[9]));
			radix2 #(.width(width)) rd_st10_10  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[10]), .rdlo_in(a10_wr[11]),  .coef_in(coef[0]), .rdup_out(a11_wr[10]), .rdlo_out(a11_wr[11]));
			radix2 #(.width(width)) rd_st10_12  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[12]), .rdlo_in(a10_wr[13]),  .coef_in(coef[0]), .rdup_out(a11_wr[12]), .rdlo_out(a11_wr[13]));
			radix2 #(.width(width)) rd_st10_14  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[14]), .rdlo_in(a10_wr[15]),  .coef_in(coef[0]), .rdup_out(a11_wr[14]), .rdlo_out(a11_wr[15]));
			radix2 #(.width(width)) rd_st10_16  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[16]), .rdlo_in(a10_wr[17]),  .coef_in(coef[0]), .rdup_out(a11_wr[16]), .rdlo_out(a11_wr[17]));
			radix2 #(.width(width)) rd_st10_18  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[18]), .rdlo_in(a10_wr[19]),  .coef_in(coef[0]), .rdup_out(a11_wr[18]), .rdlo_out(a11_wr[19]));
			radix2 #(.width(width)) rd_st10_20  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[20]), .rdlo_in(a10_wr[21]),  .coef_in(coef[0]), .rdup_out(a11_wr[20]), .rdlo_out(a11_wr[21]));
			radix2 #(.width(width)) rd_st10_22  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[22]), .rdlo_in(a10_wr[23]),  .coef_in(coef[0]), .rdup_out(a11_wr[22]), .rdlo_out(a11_wr[23]));
			radix2 #(.width(width)) rd_st10_24  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[24]), .rdlo_in(a10_wr[25]),  .coef_in(coef[0]), .rdup_out(a11_wr[24]), .rdlo_out(a11_wr[25]));
			radix2 #(.width(width)) rd_st10_26  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[26]), .rdlo_in(a10_wr[27]),  .coef_in(coef[0]), .rdup_out(a11_wr[26]), .rdlo_out(a11_wr[27]));
			radix2 #(.width(width)) rd_st10_28  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[28]), .rdlo_in(a10_wr[29]),  .coef_in(coef[0]), .rdup_out(a11_wr[28]), .rdlo_out(a11_wr[29]));
			radix2 #(.width(width)) rd_st10_30  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[30]), .rdlo_in(a10_wr[31]),  .coef_in(coef[0]), .rdup_out(a11_wr[30]), .rdlo_out(a11_wr[31]));
			radix2 #(.width(width)) rd_st10_32  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[32]), .rdlo_in(a10_wr[33]),  .coef_in(coef[0]), .rdup_out(a11_wr[32]), .rdlo_out(a11_wr[33]));
			radix2 #(.width(width)) rd_st10_34  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[34]), .rdlo_in(a10_wr[35]),  .coef_in(coef[0]), .rdup_out(a11_wr[34]), .rdlo_out(a11_wr[35]));
			radix2 #(.width(width)) rd_st10_36  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[36]), .rdlo_in(a10_wr[37]),  .coef_in(coef[0]), .rdup_out(a11_wr[36]), .rdlo_out(a11_wr[37]));
			radix2 #(.width(width)) rd_st10_38  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[38]), .rdlo_in(a10_wr[39]),  .coef_in(coef[0]), .rdup_out(a11_wr[38]), .rdlo_out(a11_wr[39]));
			radix2 #(.width(width)) rd_st10_40  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[40]), .rdlo_in(a10_wr[41]),  .coef_in(coef[0]), .rdup_out(a11_wr[40]), .rdlo_out(a11_wr[41]));
			radix2 #(.width(width)) rd_st10_42  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[42]), .rdlo_in(a10_wr[43]),  .coef_in(coef[0]), .rdup_out(a11_wr[42]), .rdlo_out(a11_wr[43]));
			radix2 #(.width(width)) rd_st10_44  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[44]), .rdlo_in(a10_wr[45]),  .coef_in(coef[0]), .rdup_out(a11_wr[44]), .rdlo_out(a11_wr[45]));
			radix2 #(.width(width)) rd_st10_46  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[46]), .rdlo_in(a10_wr[47]),  .coef_in(coef[0]), .rdup_out(a11_wr[46]), .rdlo_out(a11_wr[47]));
			radix2 #(.width(width)) rd_st10_48  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[48]), .rdlo_in(a10_wr[49]),  .coef_in(coef[0]), .rdup_out(a11_wr[48]), .rdlo_out(a11_wr[49]));
			radix2 #(.width(width)) rd_st10_50  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[50]), .rdlo_in(a10_wr[51]),  .coef_in(coef[0]), .rdup_out(a11_wr[50]), .rdlo_out(a11_wr[51]));
			radix2 #(.width(width)) rd_st10_52  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[52]), .rdlo_in(a10_wr[53]),  .coef_in(coef[0]), .rdup_out(a11_wr[52]), .rdlo_out(a11_wr[53]));
			radix2 #(.width(width)) rd_st10_54  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[54]), .rdlo_in(a10_wr[55]),  .coef_in(coef[0]), .rdup_out(a11_wr[54]), .rdlo_out(a11_wr[55]));
			radix2 #(.width(width)) rd_st10_56  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[56]), .rdlo_in(a10_wr[57]),  .coef_in(coef[0]), .rdup_out(a11_wr[56]), .rdlo_out(a11_wr[57]));
			radix2 #(.width(width)) rd_st10_58  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[58]), .rdlo_in(a10_wr[59]),  .coef_in(coef[0]), .rdup_out(a11_wr[58]), .rdlo_out(a11_wr[59]));
			radix2 #(.width(width)) rd_st10_60  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[60]), .rdlo_in(a10_wr[61]),  .coef_in(coef[0]), .rdup_out(a11_wr[60]), .rdlo_out(a11_wr[61]));
			radix2 #(.width(width)) rd_st10_62  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[62]), .rdlo_in(a10_wr[63]),  .coef_in(coef[0]), .rdup_out(a11_wr[62]), .rdlo_out(a11_wr[63]));
			radix2 #(.width(width)) rd_st10_64  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[64]), .rdlo_in(a10_wr[65]),  .coef_in(coef[0]), .rdup_out(a11_wr[64]), .rdlo_out(a11_wr[65]));
			radix2 #(.width(width)) rd_st10_66  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[66]), .rdlo_in(a10_wr[67]),  .coef_in(coef[0]), .rdup_out(a11_wr[66]), .rdlo_out(a11_wr[67]));
			radix2 #(.width(width)) rd_st10_68  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[68]), .rdlo_in(a10_wr[69]),  .coef_in(coef[0]), .rdup_out(a11_wr[68]), .rdlo_out(a11_wr[69]));
			radix2 #(.width(width)) rd_st10_70  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[70]), .rdlo_in(a10_wr[71]),  .coef_in(coef[0]), .rdup_out(a11_wr[70]), .rdlo_out(a11_wr[71]));
			radix2 #(.width(width)) rd_st10_72  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[72]), .rdlo_in(a10_wr[73]),  .coef_in(coef[0]), .rdup_out(a11_wr[72]), .rdlo_out(a11_wr[73]));
			radix2 #(.width(width)) rd_st10_74  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[74]), .rdlo_in(a10_wr[75]),  .coef_in(coef[0]), .rdup_out(a11_wr[74]), .rdlo_out(a11_wr[75]));
			radix2 #(.width(width)) rd_st10_76  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[76]), .rdlo_in(a10_wr[77]),  .coef_in(coef[0]), .rdup_out(a11_wr[76]), .rdlo_out(a11_wr[77]));
			radix2 #(.width(width)) rd_st10_78  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[78]), .rdlo_in(a10_wr[79]),  .coef_in(coef[0]), .rdup_out(a11_wr[78]), .rdlo_out(a11_wr[79]));
			radix2 #(.width(width)) rd_st10_80  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[80]), .rdlo_in(a10_wr[81]),  .coef_in(coef[0]), .rdup_out(a11_wr[80]), .rdlo_out(a11_wr[81]));
			radix2 #(.width(width)) rd_st10_82  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[82]), .rdlo_in(a10_wr[83]),  .coef_in(coef[0]), .rdup_out(a11_wr[82]), .rdlo_out(a11_wr[83]));
			radix2 #(.width(width)) rd_st10_84  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[84]), .rdlo_in(a10_wr[85]),  .coef_in(coef[0]), .rdup_out(a11_wr[84]), .rdlo_out(a11_wr[85]));
			radix2 #(.width(width)) rd_st10_86  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[86]), .rdlo_in(a10_wr[87]),  .coef_in(coef[0]), .rdup_out(a11_wr[86]), .rdlo_out(a11_wr[87]));
			radix2 #(.width(width)) rd_st10_88  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[88]), .rdlo_in(a10_wr[89]),  .coef_in(coef[0]), .rdup_out(a11_wr[88]), .rdlo_out(a11_wr[89]));
			radix2 #(.width(width)) rd_st10_90  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[90]), .rdlo_in(a10_wr[91]),  .coef_in(coef[0]), .rdup_out(a11_wr[90]), .rdlo_out(a11_wr[91]));
			radix2 #(.width(width)) rd_st10_92  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[92]), .rdlo_in(a10_wr[93]),  .coef_in(coef[0]), .rdup_out(a11_wr[92]), .rdlo_out(a11_wr[93]));
			radix2 #(.width(width)) rd_st10_94  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[94]), .rdlo_in(a10_wr[95]),  .coef_in(coef[0]), .rdup_out(a11_wr[94]), .rdlo_out(a11_wr[95]));
			radix2 #(.width(width)) rd_st10_96  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[96]), .rdlo_in(a10_wr[97]),  .coef_in(coef[0]), .rdup_out(a11_wr[96]), .rdlo_out(a11_wr[97]));
			radix2 #(.width(width)) rd_st10_98  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[98]), .rdlo_in(a10_wr[99]),  .coef_in(coef[0]), .rdup_out(a11_wr[98]), .rdlo_out(a11_wr[99]));
			radix2 #(.width(width)) rd_st10_100  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[100]), .rdlo_in(a10_wr[101]),  .coef_in(coef[0]), .rdup_out(a11_wr[100]), .rdlo_out(a11_wr[101]));
			radix2 #(.width(width)) rd_st10_102  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[102]), .rdlo_in(a10_wr[103]),  .coef_in(coef[0]), .rdup_out(a11_wr[102]), .rdlo_out(a11_wr[103]));
			radix2 #(.width(width)) rd_st10_104  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[104]), .rdlo_in(a10_wr[105]),  .coef_in(coef[0]), .rdup_out(a11_wr[104]), .rdlo_out(a11_wr[105]));
			radix2 #(.width(width)) rd_st10_106  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[106]), .rdlo_in(a10_wr[107]),  .coef_in(coef[0]), .rdup_out(a11_wr[106]), .rdlo_out(a11_wr[107]));
			radix2 #(.width(width)) rd_st10_108  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[108]), .rdlo_in(a10_wr[109]),  .coef_in(coef[0]), .rdup_out(a11_wr[108]), .rdlo_out(a11_wr[109]));
			radix2 #(.width(width)) rd_st10_110  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[110]), .rdlo_in(a10_wr[111]),  .coef_in(coef[0]), .rdup_out(a11_wr[110]), .rdlo_out(a11_wr[111]));
			radix2 #(.width(width)) rd_st10_112  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[112]), .rdlo_in(a10_wr[113]),  .coef_in(coef[0]), .rdup_out(a11_wr[112]), .rdlo_out(a11_wr[113]));
			radix2 #(.width(width)) rd_st10_114  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[114]), .rdlo_in(a10_wr[115]),  .coef_in(coef[0]), .rdup_out(a11_wr[114]), .rdlo_out(a11_wr[115]));
			radix2 #(.width(width)) rd_st10_116  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[116]), .rdlo_in(a10_wr[117]),  .coef_in(coef[0]), .rdup_out(a11_wr[116]), .rdlo_out(a11_wr[117]));
			radix2 #(.width(width)) rd_st10_118  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[118]), .rdlo_in(a10_wr[119]),  .coef_in(coef[0]), .rdup_out(a11_wr[118]), .rdlo_out(a11_wr[119]));
			radix2 #(.width(width)) rd_st10_120  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[120]), .rdlo_in(a10_wr[121]),  .coef_in(coef[0]), .rdup_out(a11_wr[120]), .rdlo_out(a11_wr[121]));
			radix2 #(.width(width)) rd_st10_122  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[122]), .rdlo_in(a10_wr[123]),  .coef_in(coef[0]), .rdup_out(a11_wr[122]), .rdlo_out(a11_wr[123]));
			radix2 #(.width(width)) rd_st10_124  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[124]), .rdlo_in(a10_wr[125]),  .coef_in(coef[0]), .rdup_out(a11_wr[124]), .rdlo_out(a11_wr[125]));
			radix2 #(.width(width)) rd_st10_126  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[126]), .rdlo_in(a10_wr[127]),  .coef_in(coef[0]), .rdup_out(a11_wr[126]), .rdlo_out(a11_wr[127]));
			radix2 #(.width(width)) rd_st10_128  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[128]), .rdlo_in(a10_wr[129]),  .coef_in(coef[0]), .rdup_out(a11_wr[128]), .rdlo_out(a11_wr[129]));
			radix2 #(.width(width)) rd_st10_130  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[130]), .rdlo_in(a10_wr[131]),  .coef_in(coef[0]), .rdup_out(a11_wr[130]), .rdlo_out(a11_wr[131]));
			radix2 #(.width(width)) rd_st10_132  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[132]), .rdlo_in(a10_wr[133]),  .coef_in(coef[0]), .rdup_out(a11_wr[132]), .rdlo_out(a11_wr[133]));
			radix2 #(.width(width)) rd_st10_134  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[134]), .rdlo_in(a10_wr[135]),  .coef_in(coef[0]), .rdup_out(a11_wr[134]), .rdlo_out(a11_wr[135]));
			radix2 #(.width(width)) rd_st10_136  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[136]), .rdlo_in(a10_wr[137]),  .coef_in(coef[0]), .rdup_out(a11_wr[136]), .rdlo_out(a11_wr[137]));
			radix2 #(.width(width)) rd_st10_138  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[138]), .rdlo_in(a10_wr[139]),  .coef_in(coef[0]), .rdup_out(a11_wr[138]), .rdlo_out(a11_wr[139]));
			radix2 #(.width(width)) rd_st10_140  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[140]), .rdlo_in(a10_wr[141]),  .coef_in(coef[0]), .rdup_out(a11_wr[140]), .rdlo_out(a11_wr[141]));
			radix2 #(.width(width)) rd_st10_142  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[142]), .rdlo_in(a10_wr[143]),  .coef_in(coef[0]), .rdup_out(a11_wr[142]), .rdlo_out(a11_wr[143]));
			radix2 #(.width(width)) rd_st10_144  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[144]), .rdlo_in(a10_wr[145]),  .coef_in(coef[0]), .rdup_out(a11_wr[144]), .rdlo_out(a11_wr[145]));
			radix2 #(.width(width)) rd_st10_146  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[146]), .rdlo_in(a10_wr[147]),  .coef_in(coef[0]), .rdup_out(a11_wr[146]), .rdlo_out(a11_wr[147]));
			radix2 #(.width(width)) rd_st10_148  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[148]), .rdlo_in(a10_wr[149]),  .coef_in(coef[0]), .rdup_out(a11_wr[148]), .rdlo_out(a11_wr[149]));
			radix2 #(.width(width)) rd_st10_150  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[150]), .rdlo_in(a10_wr[151]),  .coef_in(coef[0]), .rdup_out(a11_wr[150]), .rdlo_out(a11_wr[151]));
			radix2 #(.width(width)) rd_st10_152  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[152]), .rdlo_in(a10_wr[153]),  .coef_in(coef[0]), .rdup_out(a11_wr[152]), .rdlo_out(a11_wr[153]));
			radix2 #(.width(width)) rd_st10_154  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[154]), .rdlo_in(a10_wr[155]),  .coef_in(coef[0]), .rdup_out(a11_wr[154]), .rdlo_out(a11_wr[155]));
			radix2 #(.width(width)) rd_st10_156  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[156]), .rdlo_in(a10_wr[157]),  .coef_in(coef[0]), .rdup_out(a11_wr[156]), .rdlo_out(a11_wr[157]));
			radix2 #(.width(width)) rd_st10_158  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[158]), .rdlo_in(a10_wr[159]),  .coef_in(coef[0]), .rdup_out(a11_wr[158]), .rdlo_out(a11_wr[159]));
			radix2 #(.width(width)) rd_st10_160  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[160]), .rdlo_in(a10_wr[161]),  .coef_in(coef[0]), .rdup_out(a11_wr[160]), .rdlo_out(a11_wr[161]));
			radix2 #(.width(width)) rd_st10_162  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[162]), .rdlo_in(a10_wr[163]),  .coef_in(coef[0]), .rdup_out(a11_wr[162]), .rdlo_out(a11_wr[163]));
			radix2 #(.width(width)) rd_st10_164  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[164]), .rdlo_in(a10_wr[165]),  .coef_in(coef[0]), .rdup_out(a11_wr[164]), .rdlo_out(a11_wr[165]));
			radix2 #(.width(width)) rd_st10_166  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[166]), .rdlo_in(a10_wr[167]),  .coef_in(coef[0]), .rdup_out(a11_wr[166]), .rdlo_out(a11_wr[167]));
			radix2 #(.width(width)) rd_st10_168  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[168]), .rdlo_in(a10_wr[169]),  .coef_in(coef[0]), .rdup_out(a11_wr[168]), .rdlo_out(a11_wr[169]));
			radix2 #(.width(width)) rd_st10_170  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[170]), .rdlo_in(a10_wr[171]),  .coef_in(coef[0]), .rdup_out(a11_wr[170]), .rdlo_out(a11_wr[171]));
			radix2 #(.width(width)) rd_st10_172  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[172]), .rdlo_in(a10_wr[173]),  .coef_in(coef[0]), .rdup_out(a11_wr[172]), .rdlo_out(a11_wr[173]));
			radix2 #(.width(width)) rd_st10_174  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[174]), .rdlo_in(a10_wr[175]),  .coef_in(coef[0]), .rdup_out(a11_wr[174]), .rdlo_out(a11_wr[175]));
			radix2 #(.width(width)) rd_st10_176  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[176]), .rdlo_in(a10_wr[177]),  .coef_in(coef[0]), .rdup_out(a11_wr[176]), .rdlo_out(a11_wr[177]));
			radix2 #(.width(width)) rd_st10_178  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[178]), .rdlo_in(a10_wr[179]),  .coef_in(coef[0]), .rdup_out(a11_wr[178]), .rdlo_out(a11_wr[179]));
			radix2 #(.width(width)) rd_st10_180  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[180]), .rdlo_in(a10_wr[181]),  .coef_in(coef[0]), .rdup_out(a11_wr[180]), .rdlo_out(a11_wr[181]));
			radix2 #(.width(width)) rd_st10_182  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[182]), .rdlo_in(a10_wr[183]),  .coef_in(coef[0]), .rdup_out(a11_wr[182]), .rdlo_out(a11_wr[183]));
			radix2 #(.width(width)) rd_st10_184  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[184]), .rdlo_in(a10_wr[185]),  .coef_in(coef[0]), .rdup_out(a11_wr[184]), .rdlo_out(a11_wr[185]));
			radix2 #(.width(width)) rd_st10_186  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[186]), .rdlo_in(a10_wr[187]),  .coef_in(coef[0]), .rdup_out(a11_wr[186]), .rdlo_out(a11_wr[187]));
			radix2 #(.width(width)) rd_st10_188  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[188]), .rdlo_in(a10_wr[189]),  .coef_in(coef[0]), .rdup_out(a11_wr[188]), .rdlo_out(a11_wr[189]));
			radix2 #(.width(width)) rd_st10_190  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[190]), .rdlo_in(a10_wr[191]),  .coef_in(coef[0]), .rdup_out(a11_wr[190]), .rdlo_out(a11_wr[191]));
			radix2 #(.width(width)) rd_st10_192  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[192]), .rdlo_in(a10_wr[193]),  .coef_in(coef[0]), .rdup_out(a11_wr[192]), .rdlo_out(a11_wr[193]));
			radix2 #(.width(width)) rd_st10_194  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[194]), .rdlo_in(a10_wr[195]),  .coef_in(coef[0]), .rdup_out(a11_wr[194]), .rdlo_out(a11_wr[195]));
			radix2 #(.width(width)) rd_st10_196  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[196]), .rdlo_in(a10_wr[197]),  .coef_in(coef[0]), .rdup_out(a11_wr[196]), .rdlo_out(a11_wr[197]));
			radix2 #(.width(width)) rd_st10_198  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[198]), .rdlo_in(a10_wr[199]),  .coef_in(coef[0]), .rdup_out(a11_wr[198]), .rdlo_out(a11_wr[199]));
			radix2 #(.width(width)) rd_st10_200  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[200]), .rdlo_in(a10_wr[201]),  .coef_in(coef[0]), .rdup_out(a11_wr[200]), .rdlo_out(a11_wr[201]));
			radix2 #(.width(width)) rd_st10_202  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[202]), .rdlo_in(a10_wr[203]),  .coef_in(coef[0]), .rdup_out(a11_wr[202]), .rdlo_out(a11_wr[203]));
			radix2 #(.width(width)) rd_st10_204  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[204]), .rdlo_in(a10_wr[205]),  .coef_in(coef[0]), .rdup_out(a11_wr[204]), .rdlo_out(a11_wr[205]));
			radix2 #(.width(width)) rd_st10_206  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[206]), .rdlo_in(a10_wr[207]),  .coef_in(coef[0]), .rdup_out(a11_wr[206]), .rdlo_out(a11_wr[207]));
			radix2 #(.width(width)) rd_st10_208  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[208]), .rdlo_in(a10_wr[209]),  .coef_in(coef[0]), .rdup_out(a11_wr[208]), .rdlo_out(a11_wr[209]));
			radix2 #(.width(width)) rd_st10_210  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[210]), .rdlo_in(a10_wr[211]),  .coef_in(coef[0]), .rdup_out(a11_wr[210]), .rdlo_out(a11_wr[211]));
			radix2 #(.width(width)) rd_st10_212  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[212]), .rdlo_in(a10_wr[213]),  .coef_in(coef[0]), .rdup_out(a11_wr[212]), .rdlo_out(a11_wr[213]));
			radix2 #(.width(width)) rd_st10_214  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[214]), .rdlo_in(a10_wr[215]),  .coef_in(coef[0]), .rdup_out(a11_wr[214]), .rdlo_out(a11_wr[215]));
			radix2 #(.width(width)) rd_st10_216  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[216]), .rdlo_in(a10_wr[217]),  .coef_in(coef[0]), .rdup_out(a11_wr[216]), .rdlo_out(a11_wr[217]));
			radix2 #(.width(width)) rd_st10_218  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[218]), .rdlo_in(a10_wr[219]),  .coef_in(coef[0]), .rdup_out(a11_wr[218]), .rdlo_out(a11_wr[219]));
			radix2 #(.width(width)) rd_st10_220  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[220]), .rdlo_in(a10_wr[221]),  .coef_in(coef[0]), .rdup_out(a11_wr[220]), .rdlo_out(a11_wr[221]));
			radix2 #(.width(width)) rd_st10_222  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[222]), .rdlo_in(a10_wr[223]),  .coef_in(coef[0]), .rdup_out(a11_wr[222]), .rdlo_out(a11_wr[223]));
			radix2 #(.width(width)) rd_st10_224  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[224]), .rdlo_in(a10_wr[225]),  .coef_in(coef[0]), .rdup_out(a11_wr[224]), .rdlo_out(a11_wr[225]));
			radix2 #(.width(width)) rd_st10_226  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[226]), .rdlo_in(a10_wr[227]),  .coef_in(coef[0]), .rdup_out(a11_wr[226]), .rdlo_out(a11_wr[227]));
			radix2 #(.width(width)) rd_st10_228  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[228]), .rdlo_in(a10_wr[229]),  .coef_in(coef[0]), .rdup_out(a11_wr[228]), .rdlo_out(a11_wr[229]));
			radix2 #(.width(width)) rd_st10_230  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[230]), .rdlo_in(a10_wr[231]),  .coef_in(coef[0]), .rdup_out(a11_wr[230]), .rdlo_out(a11_wr[231]));
			radix2 #(.width(width)) rd_st10_232  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[232]), .rdlo_in(a10_wr[233]),  .coef_in(coef[0]), .rdup_out(a11_wr[232]), .rdlo_out(a11_wr[233]));
			radix2 #(.width(width)) rd_st10_234  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[234]), .rdlo_in(a10_wr[235]),  .coef_in(coef[0]), .rdup_out(a11_wr[234]), .rdlo_out(a11_wr[235]));
			radix2 #(.width(width)) rd_st10_236  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[236]), .rdlo_in(a10_wr[237]),  .coef_in(coef[0]), .rdup_out(a11_wr[236]), .rdlo_out(a11_wr[237]));
			radix2 #(.width(width)) rd_st10_238  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[238]), .rdlo_in(a10_wr[239]),  .coef_in(coef[0]), .rdup_out(a11_wr[238]), .rdlo_out(a11_wr[239]));
			radix2 #(.width(width)) rd_st10_240  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[240]), .rdlo_in(a10_wr[241]),  .coef_in(coef[0]), .rdup_out(a11_wr[240]), .rdlo_out(a11_wr[241]));
			radix2 #(.width(width)) rd_st10_242  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[242]), .rdlo_in(a10_wr[243]),  .coef_in(coef[0]), .rdup_out(a11_wr[242]), .rdlo_out(a11_wr[243]));
			radix2 #(.width(width)) rd_st10_244  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[244]), .rdlo_in(a10_wr[245]),  .coef_in(coef[0]), .rdup_out(a11_wr[244]), .rdlo_out(a11_wr[245]));
			radix2 #(.width(width)) rd_st10_246  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[246]), .rdlo_in(a10_wr[247]),  .coef_in(coef[0]), .rdup_out(a11_wr[246]), .rdlo_out(a11_wr[247]));
			radix2 #(.width(width)) rd_st10_248  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[248]), .rdlo_in(a10_wr[249]),  .coef_in(coef[0]), .rdup_out(a11_wr[248]), .rdlo_out(a11_wr[249]));
			radix2 #(.width(width)) rd_st10_250  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[250]), .rdlo_in(a10_wr[251]),  .coef_in(coef[0]), .rdup_out(a11_wr[250]), .rdlo_out(a11_wr[251]));
			radix2 #(.width(width)) rd_st10_252  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[252]), .rdlo_in(a10_wr[253]),  .coef_in(coef[0]), .rdup_out(a11_wr[252]), .rdlo_out(a11_wr[253]));
			radix2 #(.width(width)) rd_st10_254  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[254]), .rdlo_in(a10_wr[255]),  .coef_in(coef[0]), .rdup_out(a11_wr[254]), .rdlo_out(a11_wr[255]));
			radix2 #(.width(width)) rd_st10_256  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[256]), .rdlo_in(a10_wr[257]),  .coef_in(coef[0]), .rdup_out(a11_wr[256]), .rdlo_out(a11_wr[257]));
			radix2 #(.width(width)) rd_st10_258  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[258]), .rdlo_in(a10_wr[259]),  .coef_in(coef[0]), .rdup_out(a11_wr[258]), .rdlo_out(a11_wr[259]));
			radix2 #(.width(width)) rd_st10_260  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[260]), .rdlo_in(a10_wr[261]),  .coef_in(coef[0]), .rdup_out(a11_wr[260]), .rdlo_out(a11_wr[261]));
			radix2 #(.width(width)) rd_st10_262  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[262]), .rdlo_in(a10_wr[263]),  .coef_in(coef[0]), .rdup_out(a11_wr[262]), .rdlo_out(a11_wr[263]));
			radix2 #(.width(width)) rd_st10_264  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[264]), .rdlo_in(a10_wr[265]),  .coef_in(coef[0]), .rdup_out(a11_wr[264]), .rdlo_out(a11_wr[265]));
			radix2 #(.width(width)) rd_st10_266  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[266]), .rdlo_in(a10_wr[267]),  .coef_in(coef[0]), .rdup_out(a11_wr[266]), .rdlo_out(a11_wr[267]));
			radix2 #(.width(width)) rd_st10_268  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[268]), .rdlo_in(a10_wr[269]),  .coef_in(coef[0]), .rdup_out(a11_wr[268]), .rdlo_out(a11_wr[269]));
			radix2 #(.width(width)) rd_st10_270  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[270]), .rdlo_in(a10_wr[271]),  .coef_in(coef[0]), .rdup_out(a11_wr[270]), .rdlo_out(a11_wr[271]));
			radix2 #(.width(width)) rd_st10_272  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[272]), .rdlo_in(a10_wr[273]),  .coef_in(coef[0]), .rdup_out(a11_wr[272]), .rdlo_out(a11_wr[273]));
			radix2 #(.width(width)) rd_st10_274  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[274]), .rdlo_in(a10_wr[275]),  .coef_in(coef[0]), .rdup_out(a11_wr[274]), .rdlo_out(a11_wr[275]));
			radix2 #(.width(width)) rd_st10_276  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[276]), .rdlo_in(a10_wr[277]),  .coef_in(coef[0]), .rdup_out(a11_wr[276]), .rdlo_out(a11_wr[277]));
			radix2 #(.width(width)) rd_st10_278  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[278]), .rdlo_in(a10_wr[279]),  .coef_in(coef[0]), .rdup_out(a11_wr[278]), .rdlo_out(a11_wr[279]));
			radix2 #(.width(width)) rd_st10_280  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[280]), .rdlo_in(a10_wr[281]),  .coef_in(coef[0]), .rdup_out(a11_wr[280]), .rdlo_out(a11_wr[281]));
			radix2 #(.width(width)) rd_st10_282  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[282]), .rdlo_in(a10_wr[283]),  .coef_in(coef[0]), .rdup_out(a11_wr[282]), .rdlo_out(a11_wr[283]));
			radix2 #(.width(width)) rd_st10_284  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[284]), .rdlo_in(a10_wr[285]),  .coef_in(coef[0]), .rdup_out(a11_wr[284]), .rdlo_out(a11_wr[285]));
			radix2 #(.width(width)) rd_st10_286  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[286]), .rdlo_in(a10_wr[287]),  .coef_in(coef[0]), .rdup_out(a11_wr[286]), .rdlo_out(a11_wr[287]));
			radix2 #(.width(width)) rd_st10_288  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[288]), .rdlo_in(a10_wr[289]),  .coef_in(coef[0]), .rdup_out(a11_wr[288]), .rdlo_out(a11_wr[289]));
			radix2 #(.width(width)) rd_st10_290  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[290]), .rdlo_in(a10_wr[291]),  .coef_in(coef[0]), .rdup_out(a11_wr[290]), .rdlo_out(a11_wr[291]));
			radix2 #(.width(width)) rd_st10_292  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[292]), .rdlo_in(a10_wr[293]),  .coef_in(coef[0]), .rdup_out(a11_wr[292]), .rdlo_out(a11_wr[293]));
			radix2 #(.width(width)) rd_st10_294  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[294]), .rdlo_in(a10_wr[295]),  .coef_in(coef[0]), .rdup_out(a11_wr[294]), .rdlo_out(a11_wr[295]));
			radix2 #(.width(width)) rd_st10_296  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[296]), .rdlo_in(a10_wr[297]),  .coef_in(coef[0]), .rdup_out(a11_wr[296]), .rdlo_out(a11_wr[297]));
			radix2 #(.width(width)) rd_st10_298  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[298]), .rdlo_in(a10_wr[299]),  .coef_in(coef[0]), .rdup_out(a11_wr[298]), .rdlo_out(a11_wr[299]));
			radix2 #(.width(width)) rd_st10_300  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[300]), .rdlo_in(a10_wr[301]),  .coef_in(coef[0]), .rdup_out(a11_wr[300]), .rdlo_out(a11_wr[301]));
			radix2 #(.width(width)) rd_st10_302  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[302]), .rdlo_in(a10_wr[303]),  .coef_in(coef[0]), .rdup_out(a11_wr[302]), .rdlo_out(a11_wr[303]));
			radix2 #(.width(width)) rd_st10_304  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[304]), .rdlo_in(a10_wr[305]),  .coef_in(coef[0]), .rdup_out(a11_wr[304]), .rdlo_out(a11_wr[305]));
			radix2 #(.width(width)) rd_st10_306  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[306]), .rdlo_in(a10_wr[307]),  .coef_in(coef[0]), .rdup_out(a11_wr[306]), .rdlo_out(a11_wr[307]));
			radix2 #(.width(width)) rd_st10_308  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[308]), .rdlo_in(a10_wr[309]),  .coef_in(coef[0]), .rdup_out(a11_wr[308]), .rdlo_out(a11_wr[309]));
			radix2 #(.width(width)) rd_st10_310  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[310]), .rdlo_in(a10_wr[311]),  .coef_in(coef[0]), .rdup_out(a11_wr[310]), .rdlo_out(a11_wr[311]));
			radix2 #(.width(width)) rd_st10_312  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[312]), .rdlo_in(a10_wr[313]),  .coef_in(coef[0]), .rdup_out(a11_wr[312]), .rdlo_out(a11_wr[313]));
			radix2 #(.width(width)) rd_st10_314  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[314]), .rdlo_in(a10_wr[315]),  .coef_in(coef[0]), .rdup_out(a11_wr[314]), .rdlo_out(a11_wr[315]));
			radix2 #(.width(width)) rd_st10_316  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[316]), .rdlo_in(a10_wr[317]),  .coef_in(coef[0]), .rdup_out(a11_wr[316]), .rdlo_out(a11_wr[317]));
			radix2 #(.width(width)) rd_st10_318  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[318]), .rdlo_in(a10_wr[319]),  .coef_in(coef[0]), .rdup_out(a11_wr[318]), .rdlo_out(a11_wr[319]));
			radix2 #(.width(width)) rd_st10_320  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[320]), .rdlo_in(a10_wr[321]),  .coef_in(coef[0]), .rdup_out(a11_wr[320]), .rdlo_out(a11_wr[321]));
			radix2 #(.width(width)) rd_st10_322  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[322]), .rdlo_in(a10_wr[323]),  .coef_in(coef[0]), .rdup_out(a11_wr[322]), .rdlo_out(a11_wr[323]));
			radix2 #(.width(width)) rd_st10_324  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[324]), .rdlo_in(a10_wr[325]),  .coef_in(coef[0]), .rdup_out(a11_wr[324]), .rdlo_out(a11_wr[325]));
			radix2 #(.width(width)) rd_st10_326  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[326]), .rdlo_in(a10_wr[327]),  .coef_in(coef[0]), .rdup_out(a11_wr[326]), .rdlo_out(a11_wr[327]));
			radix2 #(.width(width)) rd_st10_328  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[328]), .rdlo_in(a10_wr[329]),  .coef_in(coef[0]), .rdup_out(a11_wr[328]), .rdlo_out(a11_wr[329]));
			radix2 #(.width(width)) rd_st10_330  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[330]), .rdlo_in(a10_wr[331]),  .coef_in(coef[0]), .rdup_out(a11_wr[330]), .rdlo_out(a11_wr[331]));
			radix2 #(.width(width)) rd_st10_332  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[332]), .rdlo_in(a10_wr[333]),  .coef_in(coef[0]), .rdup_out(a11_wr[332]), .rdlo_out(a11_wr[333]));
			radix2 #(.width(width)) rd_st10_334  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[334]), .rdlo_in(a10_wr[335]),  .coef_in(coef[0]), .rdup_out(a11_wr[334]), .rdlo_out(a11_wr[335]));
			radix2 #(.width(width)) rd_st10_336  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[336]), .rdlo_in(a10_wr[337]),  .coef_in(coef[0]), .rdup_out(a11_wr[336]), .rdlo_out(a11_wr[337]));
			radix2 #(.width(width)) rd_st10_338  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[338]), .rdlo_in(a10_wr[339]),  .coef_in(coef[0]), .rdup_out(a11_wr[338]), .rdlo_out(a11_wr[339]));
			radix2 #(.width(width)) rd_st10_340  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[340]), .rdlo_in(a10_wr[341]),  .coef_in(coef[0]), .rdup_out(a11_wr[340]), .rdlo_out(a11_wr[341]));
			radix2 #(.width(width)) rd_st10_342  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[342]), .rdlo_in(a10_wr[343]),  .coef_in(coef[0]), .rdup_out(a11_wr[342]), .rdlo_out(a11_wr[343]));
			radix2 #(.width(width)) rd_st10_344  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[344]), .rdlo_in(a10_wr[345]),  .coef_in(coef[0]), .rdup_out(a11_wr[344]), .rdlo_out(a11_wr[345]));
			radix2 #(.width(width)) rd_st10_346  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[346]), .rdlo_in(a10_wr[347]),  .coef_in(coef[0]), .rdup_out(a11_wr[346]), .rdlo_out(a11_wr[347]));
			radix2 #(.width(width)) rd_st10_348  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[348]), .rdlo_in(a10_wr[349]),  .coef_in(coef[0]), .rdup_out(a11_wr[348]), .rdlo_out(a11_wr[349]));
			radix2 #(.width(width)) rd_st10_350  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[350]), .rdlo_in(a10_wr[351]),  .coef_in(coef[0]), .rdup_out(a11_wr[350]), .rdlo_out(a11_wr[351]));
			radix2 #(.width(width)) rd_st10_352  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[352]), .rdlo_in(a10_wr[353]),  .coef_in(coef[0]), .rdup_out(a11_wr[352]), .rdlo_out(a11_wr[353]));
			radix2 #(.width(width)) rd_st10_354  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[354]), .rdlo_in(a10_wr[355]),  .coef_in(coef[0]), .rdup_out(a11_wr[354]), .rdlo_out(a11_wr[355]));
			radix2 #(.width(width)) rd_st10_356  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[356]), .rdlo_in(a10_wr[357]),  .coef_in(coef[0]), .rdup_out(a11_wr[356]), .rdlo_out(a11_wr[357]));
			radix2 #(.width(width)) rd_st10_358  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[358]), .rdlo_in(a10_wr[359]),  .coef_in(coef[0]), .rdup_out(a11_wr[358]), .rdlo_out(a11_wr[359]));
			radix2 #(.width(width)) rd_st10_360  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[360]), .rdlo_in(a10_wr[361]),  .coef_in(coef[0]), .rdup_out(a11_wr[360]), .rdlo_out(a11_wr[361]));
			radix2 #(.width(width)) rd_st10_362  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[362]), .rdlo_in(a10_wr[363]),  .coef_in(coef[0]), .rdup_out(a11_wr[362]), .rdlo_out(a11_wr[363]));
			radix2 #(.width(width)) rd_st10_364  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[364]), .rdlo_in(a10_wr[365]),  .coef_in(coef[0]), .rdup_out(a11_wr[364]), .rdlo_out(a11_wr[365]));
			radix2 #(.width(width)) rd_st10_366  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[366]), .rdlo_in(a10_wr[367]),  .coef_in(coef[0]), .rdup_out(a11_wr[366]), .rdlo_out(a11_wr[367]));
			radix2 #(.width(width)) rd_st10_368  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[368]), .rdlo_in(a10_wr[369]),  .coef_in(coef[0]), .rdup_out(a11_wr[368]), .rdlo_out(a11_wr[369]));
			radix2 #(.width(width)) rd_st10_370  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[370]), .rdlo_in(a10_wr[371]),  .coef_in(coef[0]), .rdup_out(a11_wr[370]), .rdlo_out(a11_wr[371]));
			radix2 #(.width(width)) rd_st10_372  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[372]), .rdlo_in(a10_wr[373]),  .coef_in(coef[0]), .rdup_out(a11_wr[372]), .rdlo_out(a11_wr[373]));
			radix2 #(.width(width)) rd_st10_374  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[374]), .rdlo_in(a10_wr[375]),  .coef_in(coef[0]), .rdup_out(a11_wr[374]), .rdlo_out(a11_wr[375]));
			radix2 #(.width(width)) rd_st10_376  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[376]), .rdlo_in(a10_wr[377]),  .coef_in(coef[0]), .rdup_out(a11_wr[376]), .rdlo_out(a11_wr[377]));
			radix2 #(.width(width)) rd_st10_378  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[378]), .rdlo_in(a10_wr[379]),  .coef_in(coef[0]), .rdup_out(a11_wr[378]), .rdlo_out(a11_wr[379]));
			radix2 #(.width(width)) rd_st10_380  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[380]), .rdlo_in(a10_wr[381]),  .coef_in(coef[0]), .rdup_out(a11_wr[380]), .rdlo_out(a11_wr[381]));
			radix2 #(.width(width)) rd_st10_382  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[382]), .rdlo_in(a10_wr[383]),  .coef_in(coef[0]), .rdup_out(a11_wr[382]), .rdlo_out(a11_wr[383]));
			radix2 #(.width(width)) rd_st10_384  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[384]), .rdlo_in(a10_wr[385]),  .coef_in(coef[0]), .rdup_out(a11_wr[384]), .rdlo_out(a11_wr[385]));
			radix2 #(.width(width)) rd_st10_386  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[386]), .rdlo_in(a10_wr[387]),  .coef_in(coef[0]), .rdup_out(a11_wr[386]), .rdlo_out(a11_wr[387]));
			radix2 #(.width(width)) rd_st10_388  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[388]), .rdlo_in(a10_wr[389]),  .coef_in(coef[0]), .rdup_out(a11_wr[388]), .rdlo_out(a11_wr[389]));
			radix2 #(.width(width)) rd_st10_390  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[390]), .rdlo_in(a10_wr[391]),  .coef_in(coef[0]), .rdup_out(a11_wr[390]), .rdlo_out(a11_wr[391]));
			radix2 #(.width(width)) rd_st10_392  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[392]), .rdlo_in(a10_wr[393]),  .coef_in(coef[0]), .rdup_out(a11_wr[392]), .rdlo_out(a11_wr[393]));
			radix2 #(.width(width)) rd_st10_394  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[394]), .rdlo_in(a10_wr[395]),  .coef_in(coef[0]), .rdup_out(a11_wr[394]), .rdlo_out(a11_wr[395]));
			radix2 #(.width(width)) rd_st10_396  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[396]), .rdlo_in(a10_wr[397]),  .coef_in(coef[0]), .rdup_out(a11_wr[396]), .rdlo_out(a11_wr[397]));
			radix2 #(.width(width)) rd_st10_398  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[398]), .rdlo_in(a10_wr[399]),  .coef_in(coef[0]), .rdup_out(a11_wr[398]), .rdlo_out(a11_wr[399]));
			radix2 #(.width(width)) rd_st10_400  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[400]), .rdlo_in(a10_wr[401]),  .coef_in(coef[0]), .rdup_out(a11_wr[400]), .rdlo_out(a11_wr[401]));
			radix2 #(.width(width)) rd_st10_402  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[402]), .rdlo_in(a10_wr[403]),  .coef_in(coef[0]), .rdup_out(a11_wr[402]), .rdlo_out(a11_wr[403]));
			radix2 #(.width(width)) rd_st10_404  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[404]), .rdlo_in(a10_wr[405]),  .coef_in(coef[0]), .rdup_out(a11_wr[404]), .rdlo_out(a11_wr[405]));
			radix2 #(.width(width)) rd_st10_406  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[406]), .rdlo_in(a10_wr[407]),  .coef_in(coef[0]), .rdup_out(a11_wr[406]), .rdlo_out(a11_wr[407]));
			radix2 #(.width(width)) rd_st10_408  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[408]), .rdlo_in(a10_wr[409]),  .coef_in(coef[0]), .rdup_out(a11_wr[408]), .rdlo_out(a11_wr[409]));
			radix2 #(.width(width)) rd_st10_410  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[410]), .rdlo_in(a10_wr[411]),  .coef_in(coef[0]), .rdup_out(a11_wr[410]), .rdlo_out(a11_wr[411]));
			radix2 #(.width(width)) rd_st10_412  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[412]), .rdlo_in(a10_wr[413]),  .coef_in(coef[0]), .rdup_out(a11_wr[412]), .rdlo_out(a11_wr[413]));
			radix2 #(.width(width)) rd_st10_414  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[414]), .rdlo_in(a10_wr[415]),  .coef_in(coef[0]), .rdup_out(a11_wr[414]), .rdlo_out(a11_wr[415]));
			radix2 #(.width(width)) rd_st10_416  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[416]), .rdlo_in(a10_wr[417]),  .coef_in(coef[0]), .rdup_out(a11_wr[416]), .rdlo_out(a11_wr[417]));
			radix2 #(.width(width)) rd_st10_418  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[418]), .rdlo_in(a10_wr[419]),  .coef_in(coef[0]), .rdup_out(a11_wr[418]), .rdlo_out(a11_wr[419]));
			radix2 #(.width(width)) rd_st10_420  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[420]), .rdlo_in(a10_wr[421]),  .coef_in(coef[0]), .rdup_out(a11_wr[420]), .rdlo_out(a11_wr[421]));
			radix2 #(.width(width)) rd_st10_422  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[422]), .rdlo_in(a10_wr[423]),  .coef_in(coef[0]), .rdup_out(a11_wr[422]), .rdlo_out(a11_wr[423]));
			radix2 #(.width(width)) rd_st10_424  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[424]), .rdlo_in(a10_wr[425]),  .coef_in(coef[0]), .rdup_out(a11_wr[424]), .rdlo_out(a11_wr[425]));
			radix2 #(.width(width)) rd_st10_426  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[426]), .rdlo_in(a10_wr[427]),  .coef_in(coef[0]), .rdup_out(a11_wr[426]), .rdlo_out(a11_wr[427]));
			radix2 #(.width(width)) rd_st10_428  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[428]), .rdlo_in(a10_wr[429]),  .coef_in(coef[0]), .rdup_out(a11_wr[428]), .rdlo_out(a11_wr[429]));
			radix2 #(.width(width)) rd_st10_430  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[430]), .rdlo_in(a10_wr[431]),  .coef_in(coef[0]), .rdup_out(a11_wr[430]), .rdlo_out(a11_wr[431]));
			radix2 #(.width(width)) rd_st10_432  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[432]), .rdlo_in(a10_wr[433]),  .coef_in(coef[0]), .rdup_out(a11_wr[432]), .rdlo_out(a11_wr[433]));
			radix2 #(.width(width)) rd_st10_434  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[434]), .rdlo_in(a10_wr[435]),  .coef_in(coef[0]), .rdup_out(a11_wr[434]), .rdlo_out(a11_wr[435]));
			radix2 #(.width(width)) rd_st10_436  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[436]), .rdlo_in(a10_wr[437]),  .coef_in(coef[0]), .rdup_out(a11_wr[436]), .rdlo_out(a11_wr[437]));
			radix2 #(.width(width)) rd_st10_438  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[438]), .rdlo_in(a10_wr[439]),  .coef_in(coef[0]), .rdup_out(a11_wr[438]), .rdlo_out(a11_wr[439]));
			radix2 #(.width(width)) rd_st10_440  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[440]), .rdlo_in(a10_wr[441]),  .coef_in(coef[0]), .rdup_out(a11_wr[440]), .rdlo_out(a11_wr[441]));
			radix2 #(.width(width)) rd_st10_442  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[442]), .rdlo_in(a10_wr[443]),  .coef_in(coef[0]), .rdup_out(a11_wr[442]), .rdlo_out(a11_wr[443]));
			radix2 #(.width(width)) rd_st10_444  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[444]), .rdlo_in(a10_wr[445]),  .coef_in(coef[0]), .rdup_out(a11_wr[444]), .rdlo_out(a11_wr[445]));
			radix2 #(.width(width)) rd_st10_446  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[446]), .rdlo_in(a10_wr[447]),  .coef_in(coef[0]), .rdup_out(a11_wr[446]), .rdlo_out(a11_wr[447]));
			radix2 #(.width(width)) rd_st10_448  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[448]), .rdlo_in(a10_wr[449]),  .coef_in(coef[0]), .rdup_out(a11_wr[448]), .rdlo_out(a11_wr[449]));
			radix2 #(.width(width)) rd_st10_450  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[450]), .rdlo_in(a10_wr[451]),  .coef_in(coef[0]), .rdup_out(a11_wr[450]), .rdlo_out(a11_wr[451]));
			radix2 #(.width(width)) rd_st10_452  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[452]), .rdlo_in(a10_wr[453]),  .coef_in(coef[0]), .rdup_out(a11_wr[452]), .rdlo_out(a11_wr[453]));
			radix2 #(.width(width)) rd_st10_454  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[454]), .rdlo_in(a10_wr[455]),  .coef_in(coef[0]), .rdup_out(a11_wr[454]), .rdlo_out(a11_wr[455]));
			radix2 #(.width(width)) rd_st10_456  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[456]), .rdlo_in(a10_wr[457]),  .coef_in(coef[0]), .rdup_out(a11_wr[456]), .rdlo_out(a11_wr[457]));
			radix2 #(.width(width)) rd_st10_458  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[458]), .rdlo_in(a10_wr[459]),  .coef_in(coef[0]), .rdup_out(a11_wr[458]), .rdlo_out(a11_wr[459]));
			radix2 #(.width(width)) rd_st10_460  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[460]), .rdlo_in(a10_wr[461]),  .coef_in(coef[0]), .rdup_out(a11_wr[460]), .rdlo_out(a11_wr[461]));
			radix2 #(.width(width)) rd_st10_462  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[462]), .rdlo_in(a10_wr[463]),  .coef_in(coef[0]), .rdup_out(a11_wr[462]), .rdlo_out(a11_wr[463]));
			radix2 #(.width(width)) rd_st10_464  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[464]), .rdlo_in(a10_wr[465]),  .coef_in(coef[0]), .rdup_out(a11_wr[464]), .rdlo_out(a11_wr[465]));
			radix2 #(.width(width)) rd_st10_466  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[466]), .rdlo_in(a10_wr[467]),  .coef_in(coef[0]), .rdup_out(a11_wr[466]), .rdlo_out(a11_wr[467]));
			radix2 #(.width(width)) rd_st10_468  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[468]), .rdlo_in(a10_wr[469]),  .coef_in(coef[0]), .rdup_out(a11_wr[468]), .rdlo_out(a11_wr[469]));
			radix2 #(.width(width)) rd_st10_470  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[470]), .rdlo_in(a10_wr[471]),  .coef_in(coef[0]), .rdup_out(a11_wr[470]), .rdlo_out(a11_wr[471]));
			radix2 #(.width(width)) rd_st10_472  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[472]), .rdlo_in(a10_wr[473]),  .coef_in(coef[0]), .rdup_out(a11_wr[472]), .rdlo_out(a11_wr[473]));
			radix2 #(.width(width)) rd_st10_474  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[474]), .rdlo_in(a10_wr[475]),  .coef_in(coef[0]), .rdup_out(a11_wr[474]), .rdlo_out(a11_wr[475]));
			radix2 #(.width(width)) rd_st10_476  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[476]), .rdlo_in(a10_wr[477]),  .coef_in(coef[0]), .rdup_out(a11_wr[476]), .rdlo_out(a11_wr[477]));
			radix2 #(.width(width)) rd_st10_478  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[478]), .rdlo_in(a10_wr[479]),  .coef_in(coef[0]), .rdup_out(a11_wr[478]), .rdlo_out(a11_wr[479]));
			radix2 #(.width(width)) rd_st10_480  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[480]), .rdlo_in(a10_wr[481]),  .coef_in(coef[0]), .rdup_out(a11_wr[480]), .rdlo_out(a11_wr[481]));
			radix2 #(.width(width)) rd_st10_482  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[482]), .rdlo_in(a10_wr[483]),  .coef_in(coef[0]), .rdup_out(a11_wr[482]), .rdlo_out(a11_wr[483]));
			radix2 #(.width(width)) rd_st10_484  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[484]), .rdlo_in(a10_wr[485]),  .coef_in(coef[0]), .rdup_out(a11_wr[484]), .rdlo_out(a11_wr[485]));
			radix2 #(.width(width)) rd_st10_486  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[486]), .rdlo_in(a10_wr[487]),  .coef_in(coef[0]), .rdup_out(a11_wr[486]), .rdlo_out(a11_wr[487]));
			radix2 #(.width(width)) rd_st10_488  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[488]), .rdlo_in(a10_wr[489]),  .coef_in(coef[0]), .rdup_out(a11_wr[488]), .rdlo_out(a11_wr[489]));
			radix2 #(.width(width)) rd_st10_490  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[490]), .rdlo_in(a10_wr[491]),  .coef_in(coef[0]), .rdup_out(a11_wr[490]), .rdlo_out(a11_wr[491]));
			radix2 #(.width(width)) rd_st10_492  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[492]), .rdlo_in(a10_wr[493]),  .coef_in(coef[0]), .rdup_out(a11_wr[492]), .rdlo_out(a11_wr[493]));
			radix2 #(.width(width)) rd_st10_494  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[494]), .rdlo_in(a10_wr[495]),  .coef_in(coef[0]), .rdup_out(a11_wr[494]), .rdlo_out(a11_wr[495]));
			radix2 #(.width(width)) rd_st10_496  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[496]), .rdlo_in(a10_wr[497]),  .coef_in(coef[0]), .rdup_out(a11_wr[496]), .rdlo_out(a11_wr[497]));
			radix2 #(.width(width)) rd_st10_498  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[498]), .rdlo_in(a10_wr[499]),  .coef_in(coef[0]), .rdup_out(a11_wr[498]), .rdlo_out(a11_wr[499]));
			radix2 #(.width(width)) rd_st10_500  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[500]), .rdlo_in(a10_wr[501]),  .coef_in(coef[0]), .rdup_out(a11_wr[500]), .rdlo_out(a11_wr[501]));
			radix2 #(.width(width)) rd_st10_502  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[502]), .rdlo_in(a10_wr[503]),  .coef_in(coef[0]), .rdup_out(a11_wr[502]), .rdlo_out(a11_wr[503]));
			radix2 #(.width(width)) rd_st10_504  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[504]), .rdlo_in(a10_wr[505]),  .coef_in(coef[0]), .rdup_out(a11_wr[504]), .rdlo_out(a11_wr[505]));
			radix2 #(.width(width)) rd_st10_506  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[506]), .rdlo_in(a10_wr[507]),  .coef_in(coef[0]), .rdup_out(a11_wr[506]), .rdlo_out(a11_wr[507]));
			radix2 #(.width(width)) rd_st10_508  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[508]), .rdlo_in(a10_wr[509]),  .coef_in(coef[0]), .rdup_out(a11_wr[508]), .rdlo_out(a11_wr[509]));
			radix2 #(.width(width)) rd_st10_510  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[510]), .rdlo_in(a10_wr[511]),  .coef_in(coef[0]), .rdup_out(a11_wr[510]), .rdlo_out(a11_wr[511]));
			radix2 #(.width(width)) rd_st10_512  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[512]), .rdlo_in(a10_wr[513]),  .coef_in(coef[0]), .rdup_out(a11_wr[512]), .rdlo_out(a11_wr[513]));
			radix2 #(.width(width)) rd_st10_514  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[514]), .rdlo_in(a10_wr[515]),  .coef_in(coef[0]), .rdup_out(a11_wr[514]), .rdlo_out(a11_wr[515]));
			radix2 #(.width(width)) rd_st10_516  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[516]), .rdlo_in(a10_wr[517]),  .coef_in(coef[0]), .rdup_out(a11_wr[516]), .rdlo_out(a11_wr[517]));
			radix2 #(.width(width)) rd_st10_518  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[518]), .rdlo_in(a10_wr[519]),  .coef_in(coef[0]), .rdup_out(a11_wr[518]), .rdlo_out(a11_wr[519]));
			radix2 #(.width(width)) rd_st10_520  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[520]), .rdlo_in(a10_wr[521]),  .coef_in(coef[0]), .rdup_out(a11_wr[520]), .rdlo_out(a11_wr[521]));
			radix2 #(.width(width)) rd_st10_522  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[522]), .rdlo_in(a10_wr[523]),  .coef_in(coef[0]), .rdup_out(a11_wr[522]), .rdlo_out(a11_wr[523]));
			radix2 #(.width(width)) rd_st10_524  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[524]), .rdlo_in(a10_wr[525]),  .coef_in(coef[0]), .rdup_out(a11_wr[524]), .rdlo_out(a11_wr[525]));
			radix2 #(.width(width)) rd_st10_526  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[526]), .rdlo_in(a10_wr[527]),  .coef_in(coef[0]), .rdup_out(a11_wr[526]), .rdlo_out(a11_wr[527]));
			radix2 #(.width(width)) rd_st10_528  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[528]), .rdlo_in(a10_wr[529]),  .coef_in(coef[0]), .rdup_out(a11_wr[528]), .rdlo_out(a11_wr[529]));
			radix2 #(.width(width)) rd_st10_530  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[530]), .rdlo_in(a10_wr[531]),  .coef_in(coef[0]), .rdup_out(a11_wr[530]), .rdlo_out(a11_wr[531]));
			radix2 #(.width(width)) rd_st10_532  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[532]), .rdlo_in(a10_wr[533]),  .coef_in(coef[0]), .rdup_out(a11_wr[532]), .rdlo_out(a11_wr[533]));
			radix2 #(.width(width)) rd_st10_534  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[534]), .rdlo_in(a10_wr[535]),  .coef_in(coef[0]), .rdup_out(a11_wr[534]), .rdlo_out(a11_wr[535]));
			radix2 #(.width(width)) rd_st10_536  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[536]), .rdlo_in(a10_wr[537]),  .coef_in(coef[0]), .rdup_out(a11_wr[536]), .rdlo_out(a11_wr[537]));
			radix2 #(.width(width)) rd_st10_538  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[538]), .rdlo_in(a10_wr[539]),  .coef_in(coef[0]), .rdup_out(a11_wr[538]), .rdlo_out(a11_wr[539]));
			radix2 #(.width(width)) rd_st10_540  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[540]), .rdlo_in(a10_wr[541]),  .coef_in(coef[0]), .rdup_out(a11_wr[540]), .rdlo_out(a11_wr[541]));
			radix2 #(.width(width)) rd_st10_542  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[542]), .rdlo_in(a10_wr[543]),  .coef_in(coef[0]), .rdup_out(a11_wr[542]), .rdlo_out(a11_wr[543]));
			radix2 #(.width(width)) rd_st10_544  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[544]), .rdlo_in(a10_wr[545]),  .coef_in(coef[0]), .rdup_out(a11_wr[544]), .rdlo_out(a11_wr[545]));
			radix2 #(.width(width)) rd_st10_546  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[546]), .rdlo_in(a10_wr[547]),  .coef_in(coef[0]), .rdup_out(a11_wr[546]), .rdlo_out(a11_wr[547]));
			radix2 #(.width(width)) rd_st10_548  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[548]), .rdlo_in(a10_wr[549]),  .coef_in(coef[0]), .rdup_out(a11_wr[548]), .rdlo_out(a11_wr[549]));
			radix2 #(.width(width)) rd_st10_550  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[550]), .rdlo_in(a10_wr[551]),  .coef_in(coef[0]), .rdup_out(a11_wr[550]), .rdlo_out(a11_wr[551]));
			radix2 #(.width(width)) rd_st10_552  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[552]), .rdlo_in(a10_wr[553]),  .coef_in(coef[0]), .rdup_out(a11_wr[552]), .rdlo_out(a11_wr[553]));
			radix2 #(.width(width)) rd_st10_554  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[554]), .rdlo_in(a10_wr[555]),  .coef_in(coef[0]), .rdup_out(a11_wr[554]), .rdlo_out(a11_wr[555]));
			radix2 #(.width(width)) rd_st10_556  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[556]), .rdlo_in(a10_wr[557]),  .coef_in(coef[0]), .rdup_out(a11_wr[556]), .rdlo_out(a11_wr[557]));
			radix2 #(.width(width)) rd_st10_558  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[558]), .rdlo_in(a10_wr[559]),  .coef_in(coef[0]), .rdup_out(a11_wr[558]), .rdlo_out(a11_wr[559]));
			radix2 #(.width(width)) rd_st10_560  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[560]), .rdlo_in(a10_wr[561]),  .coef_in(coef[0]), .rdup_out(a11_wr[560]), .rdlo_out(a11_wr[561]));
			radix2 #(.width(width)) rd_st10_562  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[562]), .rdlo_in(a10_wr[563]),  .coef_in(coef[0]), .rdup_out(a11_wr[562]), .rdlo_out(a11_wr[563]));
			radix2 #(.width(width)) rd_st10_564  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[564]), .rdlo_in(a10_wr[565]),  .coef_in(coef[0]), .rdup_out(a11_wr[564]), .rdlo_out(a11_wr[565]));
			radix2 #(.width(width)) rd_st10_566  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[566]), .rdlo_in(a10_wr[567]),  .coef_in(coef[0]), .rdup_out(a11_wr[566]), .rdlo_out(a11_wr[567]));
			radix2 #(.width(width)) rd_st10_568  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[568]), .rdlo_in(a10_wr[569]),  .coef_in(coef[0]), .rdup_out(a11_wr[568]), .rdlo_out(a11_wr[569]));
			radix2 #(.width(width)) rd_st10_570  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[570]), .rdlo_in(a10_wr[571]),  .coef_in(coef[0]), .rdup_out(a11_wr[570]), .rdlo_out(a11_wr[571]));
			radix2 #(.width(width)) rd_st10_572  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[572]), .rdlo_in(a10_wr[573]),  .coef_in(coef[0]), .rdup_out(a11_wr[572]), .rdlo_out(a11_wr[573]));
			radix2 #(.width(width)) rd_st10_574  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[574]), .rdlo_in(a10_wr[575]),  .coef_in(coef[0]), .rdup_out(a11_wr[574]), .rdlo_out(a11_wr[575]));
			radix2 #(.width(width)) rd_st10_576  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[576]), .rdlo_in(a10_wr[577]),  .coef_in(coef[0]), .rdup_out(a11_wr[576]), .rdlo_out(a11_wr[577]));
			radix2 #(.width(width)) rd_st10_578  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[578]), .rdlo_in(a10_wr[579]),  .coef_in(coef[0]), .rdup_out(a11_wr[578]), .rdlo_out(a11_wr[579]));
			radix2 #(.width(width)) rd_st10_580  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[580]), .rdlo_in(a10_wr[581]),  .coef_in(coef[0]), .rdup_out(a11_wr[580]), .rdlo_out(a11_wr[581]));
			radix2 #(.width(width)) rd_st10_582  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[582]), .rdlo_in(a10_wr[583]),  .coef_in(coef[0]), .rdup_out(a11_wr[582]), .rdlo_out(a11_wr[583]));
			radix2 #(.width(width)) rd_st10_584  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[584]), .rdlo_in(a10_wr[585]),  .coef_in(coef[0]), .rdup_out(a11_wr[584]), .rdlo_out(a11_wr[585]));
			radix2 #(.width(width)) rd_st10_586  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[586]), .rdlo_in(a10_wr[587]),  .coef_in(coef[0]), .rdup_out(a11_wr[586]), .rdlo_out(a11_wr[587]));
			radix2 #(.width(width)) rd_st10_588  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[588]), .rdlo_in(a10_wr[589]),  .coef_in(coef[0]), .rdup_out(a11_wr[588]), .rdlo_out(a11_wr[589]));
			radix2 #(.width(width)) rd_st10_590  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[590]), .rdlo_in(a10_wr[591]),  .coef_in(coef[0]), .rdup_out(a11_wr[590]), .rdlo_out(a11_wr[591]));
			radix2 #(.width(width)) rd_st10_592  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[592]), .rdlo_in(a10_wr[593]),  .coef_in(coef[0]), .rdup_out(a11_wr[592]), .rdlo_out(a11_wr[593]));
			radix2 #(.width(width)) rd_st10_594  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[594]), .rdlo_in(a10_wr[595]),  .coef_in(coef[0]), .rdup_out(a11_wr[594]), .rdlo_out(a11_wr[595]));
			radix2 #(.width(width)) rd_st10_596  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[596]), .rdlo_in(a10_wr[597]),  .coef_in(coef[0]), .rdup_out(a11_wr[596]), .rdlo_out(a11_wr[597]));
			radix2 #(.width(width)) rd_st10_598  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[598]), .rdlo_in(a10_wr[599]),  .coef_in(coef[0]), .rdup_out(a11_wr[598]), .rdlo_out(a11_wr[599]));
			radix2 #(.width(width)) rd_st10_600  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[600]), .rdlo_in(a10_wr[601]),  .coef_in(coef[0]), .rdup_out(a11_wr[600]), .rdlo_out(a11_wr[601]));
			radix2 #(.width(width)) rd_st10_602  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[602]), .rdlo_in(a10_wr[603]),  .coef_in(coef[0]), .rdup_out(a11_wr[602]), .rdlo_out(a11_wr[603]));
			radix2 #(.width(width)) rd_st10_604  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[604]), .rdlo_in(a10_wr[605]),  .coef_in(coef[0]), .rdup_out(a11_wr[604]), .rdlo_out(a11_wr[605]));
			radix2 #(.width(width)) rd_st10_606  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[606]), .rdlo_in(a10_wr[607]),  .coef_in(coef[0]), .rdup_out(a11_wr[606]), .rdlo_out(a11_wr[607]));
			radix2 #(.width(width)) rd_st10_608  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[608]), .rdlo_in(a10_wr[609]),  .coef_in(coef[0]), .rdup_out(a11_wr[608]), .rdlo_out(a11_wr[609]));
			radix2 #(.width(width)) rd_st10_610  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[610]), .rdlo_in(a10_wr[611]),  .coef_in(coef[0]), .rdup_out(a11_wr[610]), .rdlo_out(a11_wr[611]));
			radix2 #(.width(width)) rd_st10_612  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[612]), .rdlo_in(a10_wr[613]),  .coef_in(coef[0]), .rdup_out(a11_wr[612]), .rdlo_out(a11_wr[613]));
			radix2 #(.width(width)) rd_st10_614  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[614]), .rdlo_in(a10_wr[615]),  .coef_in(coef[0]), .rdup_out(a11_wr[614]), .rdlo_out(a11_wr[615]));
			radix2 #(.width(width)) rd_st10_616  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[616]), .rdlo_in(a10_wr[617]),  .coef_in(coef[0]), .rdup_out(a11_wr[616]), .rdlo_out(a11_wr[617]));
			radix2 #(.width(width)) rd_st10_618  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[618]), .rdlo_in(a10_wr[619]),  .coef_in(coef[0]), .rdup_out(a11_wr[618]), .rdlo_out(a11_wr[619]));
			radix2 #(.width(width)) rd_st10_620  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[620]), .rdlo_in(a10_wr[621]),  .coef_in(coef[0]), .rdup_out(a11_wr[620]), .rdlo_out(a11_wr[621]));
			radix2 #(.width(width)) rd_st10_622  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[622]), .rdlo_in(a10_wr[623]),  .coef_in(coef[0]), .rdup_out(a11_wr[622]), .rdlo_out(a11_wr[623]));
			radix2 #(.width(width)) rd_st10_624  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[624]), .rdlo_in(a10_wr[625]),  .coef_in(coef[0]), .rdup_out(a11_wr[624]), .rdlo_out(a11_wr[625]));
			radix2 #(.width(width)) rd_st10_626  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[626]), .rdlo_in(a10_wr[627]),  .coef_in(coef[0]), .rdup_out(a11_wr[626]), .rdlo_out(a11_wr[627]));
			radix2 #(.width(width)) rd_st10_628  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[628]), .rdlo_in(a10_wr[629]),  .coef_in(coef[0]), .rdup_out(a11_wr[628]), .rdlo_out(a11_wr[629]));
			radix2 #(.width(width)) rd_st10_630  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[630]), .rdlo_in(a10_wr[631]),  .coef_in(coef[0]), .rdup_out(a11_wr[630]), .rdlo_out(a11_wr[631]));
			radix2 #(.width(width)) rd_st10_632  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[632]), .rdlo_in(a10_wr[633]),  .coef_in(coef[0]), .rdup_out(a11_wr[632]), .rdlo_out(a11_wr[633]));
			radix2 #(.width(width)) rd_st10_634  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[634]), .rdlo_in(a10_wr[635]),  .coef_in(coef[0]), .rdup_out(a11_wr[634]), .rdlo_out(a11_wr[635]));
			radix2 #(.width(width)) rd_st10_636  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[636]), .rdlo_in(a10_wr[637]),  .coef_in(coef[0]), .rdup_out(a11_wr[636]), .rdlo_out(a11_wr[637]));
			radix2 #(.width(width)) rd_st10_638  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[638]), .rdlo_in(a10_wr[639]),  .coef_in(coef[0]), .rdup_out(a11_wr[638]), .rdlo_out(a11_wr[639]));
			radix2 #(.width(width)) rd_st10_640  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[640]), .rdlo_in(a10_wr[641]),  .coef_in(coef[0]), .rdup_out(a11_wr[640]), .rdlo_out(a11_wr[641]));
			radix2 #(.width(width)) rd_st10_642  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[642]), .rdlo_in(a10_wr[643]),  .coef_in(coef[0]), .rdup_out(a11_wr[642]), .rdlo_out(a11_wr[643]));
			radix2 #(.width(width)) rd_st10_644  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[644]), .rdlo_in(a10_wr[645]),  .coef_in(coef[0]), .rdup_out(a11_wr[644]), .rdlo_out(a11_wr[645]));
			radix2 #(.width(width)) rd_st10_646  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[646]), .rdlo_in(a10_wr[647]),  .coef_in(coef[0]), .rdup_out(a11_wr[646]), .rdlo_out(a11_wr[647]));
			radix2 #(.width(width)) rd_st10_648  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[648]), .rdlo_in(a10_wr[649]),  .coef_in(coef[0]), .rdup_out(a11_wr[648]), .rdlo_out(a11_wr[649]));
			radix2 #(.width(width)) rd_st10_650  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[650]), .rdlo_in(a10_wr[651]),  .coef_in(coef[0]), .rdup_out(a11_wr[650]), .rdlo_out(a11_wr[651]));
			radix2 #(.width(width)) rd_st10_652  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[652]), .rdlo_in(a10_wr[653]),  .coef_in(coef[0]), .rdup_out(a11_wr[652]), .rdlo_out(a11_wr[653]));
			radix2 #(.width(width)) rd_st10_654  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[654]), .rdlo_in(a10_wr[655]),  .coef_in(coef[0]), .rdup_out(a11_wr[654]), .rdlo_out(a11_wr[655]));
			radix2 #(.width(width)) rd_st10_656  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[656]), .rdlo_in(a10_wr[657]),  .coef_in(coef[0]), .rdup_out(a11_wr[656]), .rdlo_out(a11_wr[657]));
			radix2 #(.width(width)) rd_st10_658  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[658]), .rdlo_in(a10_wr[659]),  .coef_in(coef[0]), .rdup_out(a11_wr[658]), .rdlo_out(a11_wr[659]));
			radix2 #(.width(width)) rd_st10_660  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[660]), .rdlo_in(a10_wr[661]),  .coef_in(coef[0]), .rdup_out(a11_wr[660]), .rdlo_out(a11_wr[661]));
			radix2 #(.width(width)) rd_st10_662  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[662]), .rdlo_in(a10_wr[663]),  .coef_in(coef[0]), .rdup_out(a11_wr[662]), .rdlo_out(a11_wr[663]));
			radix2 #(.width(width)) rd_st10_664  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[664]), .rdlo_in(a10_wr[665]),  .coef_in(coef[0]), .rdup_out(a11_wr[664]), .rdlo_out(a11_wr[665]));
			radix2 #(.width(width)) rd_st10_666  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[666]), .rdlo_in(a10_wr[667]),  .coef_in(coef[0]), .rdup_out(a11_wr[666]), .rdlo_out(a11_wr[667]));
			radix2 #(.width(width)) rd_st10_668  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[668]), .rdlo_in(a10_wr[669]),  .coef_in(coef[0]), .rdup_out(a11_wr[668]), .rdlo_out(a11_wr[669]));
			radix2 #(.width(width)) rd_st10_670  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[670]), .rdlo_in(a10_wr[671]),  .coef_in(coef[0]), .rdup_out(a11_wr[670]), .rdlo_out(a11_wr[671]));
			radix2 #(.width(width)) rd_st10_672  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[672]), .rdlo_in(a10_wr[673]),  .coef_in(coef[0]), .rdup_out(a11_wr[672]), .rdlo_out(a11_wr[673]));
			radix2 #(.width(width)) rd_st10_674  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[674]), .rdlo_in(a10_wr[675]),  .coef_in(coef[0]), .rdup_out(a11_wr[674]), .rdlo_out(a11_wr[675]));
			radix2 #(.width(width)) rd_st10_676  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[676]), .rdlo_in(a10_wr[677]),  .coef_in(coef[0]), .rdup_out(a11_wr[676]), .rdlo_out(a11_wr[677]));
			radix2 #(.width(width)) rd_st10_678  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[678]), .rdlo_in(a10_wr[679]),  .coef_in(coef[0]), .rdup_out(a11_wr[678]), .rdlo_out(a11_wr[679]));
			radix2 #(.width(width)) rd_st10_680  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[680]), .rdlo_in(a10_wr[681]),  .coef_in(coef[0]), .rdup_out(a11_wr[680]), .rdlo_out(a11_wr[681]));
			radix2 #(.width(width)) rd_st10_682  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[682]), .rdlo_in(a10_wr[683]),  .coef_in(coef[0]), .rdup_out(a11_wr[682]), .rdlo_out(a11_wr[683]));
			radix2 #(.width(width)) rd_st10_684  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[684]), .rdlo_in(a10_wr[685]),  .coef_in(coef[0]), .rdup_out(a11_wr[684]), .rdlo_out(a11_wr[685]));
			radix2 #(.width(width)) rd_st10_686  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[686]), .rdlo_in(a10_wr[687]),  .coef_in(coef[0]), .rdup_out(a11_wr[686]), .rdlo_out(a11_wr[687]));
			radix2 #(.width(width)) rd_st10_688  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[688]), .rdlo_in(a10_wr[689]),  .coef_in(coef[0]), .rdup_out(a11_wr[688]), .rdlo_out(a11_wr[689]));
			radix2 #(.width(width)) rd_st10_690  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[690]), .rdlo_in(a10_wr[691]),  .coef_in(coef[0]), .rdup_out(a11_wr[690]), .rdlo_out(a11_wr[691]));
			radix2 #(.width(width)) rd_st10_692  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[692]), .rdlo_in(a10_wr[693]),  .coef_in(coef[0]), .rdup_out(a11_wr[692]), .rdlo_out(a11_wr[693]));
			radix2 #(.width(width)) rd_st10_694  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[694]), .rdlo_in(a10_wr[695]),  .coef_in(coef[0]), .rdup_out(a11_wr[694]), .rdlo_out(a11_wr[695]));
			radix2 #(.width(width)) rd_st10_696  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[696]), .rdlo_in(a10_wr[697]),  .coef_in(coef[0]), .rdup_out(a11_wr[696]), .rdlo_out(a11_wr[697]));
			radix2 #(.width(width)) rd_st10_698  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[698]), .rdlo_in(a10_wr[699]),  .coef_in(coef[0]), .rdup_out(a11_wr[698]), .rdlo_out(a11_wr[699]));
			radix2 #(.width(width)) rd_st10_700  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[700]), .rdlo_in(a10_wr[701]),  .coef_in(coef[0]), .rdup_out(a11_wr[700]), .rdlo_out(a11_wr[701]));
			radix2 #(.width(width)) rd_st10_702  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[702]), .rdlo_in(a10_wr[703]),  .coef_in(coef[0]), .rdup_out(a11_wr[702]), .rdlo_out(a11_wr[703]));
			radix2 #(.width(width)) rd_st10_704  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[704]), .rdlo_in(a10_wr[705]),  .coef_in(coef[0]), .rdup_out(a11_wr[704]), .rdlo_out(a11_wr[705]));
			radix2 #(.width(width)) rd_st10_706  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[706]), .rdlo_in(a10_wr[707]),  .coef_in(coef[0]), .rdup_out(a11_wr[706]), .rdlo_out(a11_wr[707]));
			radix2 #(.width(width)) rd_st10_708  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[708]), .rdlo_in(a10_wr[709]),  .coef_in(coef[0]), .rdup_out(a11_wr[708]), .rdlo_out(a11_wr[709]));
			radix2 #(.width(width)) rd_st10_710  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[710]), .rdlo_in(a10_wr[711]),  .coef_in(coef[0]), .rdup_out(a11_wr[710]), .rdlo_out(a11_wr[711]));
			radix2 #(.width(width)) rd_st10_712  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[712]), .rdlo_in(a10_wr[713]),  .coef_in(coef[0]), .rdup_out(a11_wr[712]), .rdlo_out(a11_wr[713]));
			radix2 #(.width(width)) rd_st10_714  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[714]), .rdlo_in(a10_wr[715]),  .coef_in(coef[0]), .rdup_out(a11_wr[714]), .rdlo_out(a11_wr[715]));
			radix2 #(.width(width)) rd_st10_716  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[716]), .rdlo_in(a10_wr[717]),  .coef_in(coef[0]), .rdup_out(a11_wr[716]), .rdlo_out(a11_wr[717]));
			radix2 #(.width(width)) rd_st10_718  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[718]), .rdlo_in(a10_wr[719]),  .coef_in(coef[0]), .rdup_out(a11_wr[718]), .rdlo_out(a11_wr[719]));
			radix2 #(.width(width)) rd_st10_720  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[720]), .rdlo_in(a10_wr[721]),  .coef_in(coef[0]), .rdup_out(a11_wr[720]), .rdlo_out(a11_wr[721]));
			radix2 #(.width(width)) rd_st10_722  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[722]), .rdlo_in(a10_wr[723]),  .coef_in(coef[0]), .rdup_out(a11_wr[722]), .rdlo_out(a11_wr[723]));
			radix2 #(.width(width)) rd_st10_724  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[724]), .rdlo_in(a10_wr[725]),  .coef_in(coef[0]), .rdup_out(a11_wr[724]), .rdlo_out(a11_wr[725]));
			radix2 #(.width(width)) rd_st10_726  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[726]), .rdlo_in(a10_wr[727]),  .coef_in(coef[0]), .rdup_out(a11_wr[726]), .rdlo_out(a11_wr[727]));
			radix2 #(.width(width)) rd_st10_728  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[728]), .rdlo_in(a10_wr[729]),  .coef_in(coef[0]), .rdup_out(a11_wr[728]), .rdlo_out(a11_wr[729]));
			radix2 #(.width(width)) rd_st10_730  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[730]), .rdlo_in(a10_wr[731]),  .coef_in(coef[0]), .rdup_out(a11_wr[730]), .rdlo_out(a11_wr[731]));
			radix2 #(.width(width)) rd_st10_732  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[732]), .rdlo_in(a10_wr[733]),  .coef_in(coef[0]), .rdup_out(a11_wr[732]), .rdlo_out(a11_wr[733]));
			radix2 #(.width(width)) rd_st10_734  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[734]), .rdlo_in(a10_wr[735]),  .coef_in(coef[0]), .rdup_out(a11_wr[734]), .rdlo_out(a11_wr[735]));
			radix2 #(.width(width)) rd_st10_736  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[736]), .rdlo_in(a10_wr[737]),  .coef_in(coef[0]), .rdup_out(a11_wr[736]), .rdlo_out(a11_wr[737]));
			radix2 #(.width(width)) rd_st10_738  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[738]), .rdlo_in(a10_wr[739]),  .coef_in(coef[0]), .rdup_out(a11_wr[738]), .rdlo_out(a11_wr[739]));
			radix2 #(.width(width)) rd_st10_740  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[740]), .rdlo_in(a10_wr[741]),  .coef_in(coef[0]), .rdup_out(a11_wr[740]), .rdlo_out(a11_wr[741]));
			radix2 #(.width(width)) rd_st10_742  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[742]), .rdlo_in(a10_wr[743]),  .coef_in(coef[0]), .rdup_out(a11_wr[742]), .rdlo_out(a11_wr[743]));
			radix2 #(.width(width)) rd_st10_744  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[744]), .rdlo_in(a10_wr[745]),  .coef_in(coef[0]), .rdup_out(a11_wr[744]), .rdlo_out(a11_wr[745]));
			radix2 #(.width(width)) rd_st10_746  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[746]), .rdlo_in(a10_wr[747]),  .coef_in(coef[0]), .rdup_out(a11_wr[746]), .rdlo_out(a11_wr[747]));
			radix2 #(.width(width)) rd_st10_748  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[748]), .rdlo_in(a10_wr[749]),  .coef_in(coef[0]), .rdup_out(a11_wr[748]), .rdlo_out(a11_wr[749]));
			radix2 #(.width(width)) rd_st10_750  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[750]), .rdlo_in(a10_wr[751]),  .coef_in(coef[0]), .rdup_out(a11_wr[750]), .rdlo_out(a11_wr[751]));
			radix2 #(.width(width)) rd_st10_752  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[752]), .rdlo_in(a10_wr[753]),  .coef_in(coef[0]), .rdup_out(a11_wr[752]), .rdlo_out(a11_wr[753]));
			radix2 #(.width(width)) rd_st10_754  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[754]), .rdlo_in(a10_wr[755]),  .coef_in(coef[0]), .rdup_out(a11_wr[754]), .rdlo_out(a11_wr[755]));
			radix2 #(.width(width)) rd_st10_756  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[756]), .rdlo_in(a10_wr[757]),  .coef_in(coef[0]), .rdup_out(a11_wr[756]), .rdlo_out(a11_wr[757]));
			radix2 #(.width(width)) rd_st10_758  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[758]), .rdlo_in(a10_wr[759]),  .coef_in(coef[0]), .rdup_out(a11_wr[758]), .rdlo_out(a11_wr[759]));
			radix2 #(.width(width)) rd_st10_760  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[760]), .rdlo_in(a10_wr[761]),  .coef_in(coef[0]), .rdup_out(a11_wr[760]), .rdlo_out(a11_wr[761]));
			radix2 #(.width(width)) rd_st10_762  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[762]), .rdlo_in(a10_wr[763]),  .coef_in(coef[0]), .rdup_out(a11_wr[762]), .rdlo_out(a11_wr[763]));
			radix2 #(.width(width)) rd_st10_764  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[764]), .rdlo_in(a10_wr[765]),  .coef_in(coef[0]), .rdup_out(a11_wr[764]), .rdlo_out(a11_wr[765]));
			radix2 #(.width(width)) rd_st10_766  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[766]), .rdlo_in(a10_wr[767]),  .coef_in(coef[0]), .rdup_out(a11_wr[766]), .rdlo_out(a11_wr[767]));
			radix2 #(.width(width)) rd_st10_768  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[768]), .rdlo_in(a10_wr[769]),  .coef_in(coef[0]), .rdup_out(a11_wr[768]), .rdlo_out(a11_wr[769]));
			radix2 #(.width(width)) rd_st10_770  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[770]), .rdlo_in(a10_wr[771]),  .coef_in(coef[0]), .rdup_out(a11_wr[770]), .rdlo_out(a11_wr[771]));
			radix2 #(.width(width)) rd_st10_772  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[772]), .rdlo_in(a10_wr[773]),  .coef_in(coef[0]), .rdup_out(a11_wr[772]), .rdlo_out(a11_wr[773]));
			radix2 #(.width(width)) rd_st10_774  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[774]), .rdlo_in(a10_wr[775]),  .coef_in(coef[0]), .rdup_out(a11_wr[774]), .rdlo_out(a11_wr[775]));
			radix2 #(.width(width)) rd_st10_776  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[776]), .rdlo_in(a10_wr[777]),  .coef_in(coef[0]), .rdup_out(a11_wr[776]), .rdlo_out(a11_wr[777]));
			radix2 #(.width(width)) rd_st10_778  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[778]), .rdlo_in(a10_wr[779]),  .coef_in(coef[0]), .rdup_out(a11_wr[778]), .rdlo_out(a11_wr[779]));
			radix2 #(.width(width)) rd_st10_780  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[780]), .rdlo_in(a10_wr[781]),  .coef_in(coef[0]), .rdup_out(a11_wr[780]), .rdlo_out(a11_wr[781]));
			radix2 #(.width(width)) rd_st10_782  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[782]), .rdlo_in(a10_wr[783]),  .coef_in(coef[0]), .rdup_out(a11_wr[782]), .rdlo_out(a11_wr[783]));
			radix2 #(.width(width)) rd_st10_784  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[784]), .rdlo_in(a10_wr[785]),  .coef_in(coef[0]), .rdup_out(a11_wr[784]), .rdlo_out(a11_wr[785]));
			radix2 #(.width(width)) rd_st10_786  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[786]), .rdlo_in(a10_wr[787]),  .coef_in(coef[0]), .rdup_out(a11_wr[786]), .rdlo_out(a11_wr[787]));
			radix2 #(.width(width)) rd_st10_788  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[788]), .rdlo_in(a10_wr[789]),  .coef_in(coef[0]), .rdup_out(a11_wr[788]), .rdlo_out(a11_wr[789]));
			radix2 #(.width(width)) rd_st10_790  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[790]), .rdlo_in(a10_wr[791]),  .coef_in(coef[0]), .rdup_out(a11_wr[790]), .rdlo_out(a11_wr[791]));
			radix2 #(.width(width)) rd_st10_792  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[792]), .rdlo_in(a10_wr[793]),  .coef_in(coef[0]), .rdup_out(a11_wr[792]), .rdlo_out(a11_wr[793]));
			radix2 #(.width(width)) rd_st10_794  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[794]), .rdlo_in(a10_wr[795]),  .coef_in(coef[0]), .rdup_out(a11_wr[794]), .rdlo_out(a11_wr[795]));
			radix2 #(.width(width)) rd_st10_796  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[796]), .rdlo_in(a10_wr[797]),  .coef_in(coef[0]), .rdup_out(a11_wr[796]), .rdlo_out(a11_wr[797]));
			radix2 #(.width(width)) rd_st10_798  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[798]), .rdlo_in(a10_wr[799]),  .coef_in(coef[0]), .rdup_out(a11_wr[798]), .rdlo_out(a11_wr[799]));
			radix2 #(.width(width)) rd_st10_800  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[800]), .rdlo_in(a10_wr[801]),  .coef_in(coef[0]), .rdup_out(a11_wr[800]), .rdlo_out(a11_wr[801]));
			radix2 #(.width(width)) rd_st10_802  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[802]), .rdlo_in(a10_wr[803]),  .coef_in(coef[0]), .rdup_out(a11_wr[802]), .rdlo_out(a11_wr[803]));
			radix2 #(.width(width)) rd_st10_804  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[804]), .rdlo_in(a10_wr[805]),  .coef_in(coef[0]), .rdup_out(a11_wr[804]), .rdlo_out(a11_wr[805]));
			radix2 #(.width(width)) rd_st10_806  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[806]), .rdlo_in(a10_wr[807]),  .coef_in(coef[0]), .rdup_out(a11_wr[806]), .rdlo_out(a11_wr[807]));
			radix2 #(.width(width)) rd_st10_808  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[808]), .rdlo_in(a10_wr[809]),  .coef_in(coef[0]), .rdup_out(a11_wr[808]), .rdlo_out(a11_wr[809]));
			radix2 #(.width(width)) rd_st10_810  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[810]), .rdlo_in(a10_wr[811]),  .coef_in(coef[0]), .rdup_out(a11_wr[810]), .rdlo_out(a11_wr[811]));
			radix2 #(.width(width)) rd_st10_812  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[812]), .rdlo_in(a10_wr[813]),  .coef_in(coef[0]), .rdup_out(a11_wr[812]), .rdlo_out(a11_wr[813]));
			radix2 #(.width(width)) rd_st10_814  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[814]), .rdlo_in(a10_wr[815]),  .coef_in(coef[0]), .rdup_out(a11_wr[814]), .rdlo_out(a11_wr[815]));
			radix2 #(.width(width)) rd_st10_816  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[816]), .rdlo_in(a10_wr[817]),  .coef_in(coef[0]), .rdup_out(a11_wr[816]), .rdlo_out(a11_wr[817]));
			radix2 #(.width(width)) rd_st10_818  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[818]), .rdlo_in(a10_wr[819]),  .coef_in(coef[0]), .rdup_out(a11_wr[818]), .rdlo_out(a11_wr[819]));
			radix2 #(.width(width)) rd_st10_820  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[820]), .rdlo_in(a10_wr[821]),  .coef_in(coef[0]), .rdup_out(a11_wr[820]), .rdlo_out(a11_wr[821]));
			radix2 #(.width(width)) rd_st10_822  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[822]), .rdlo_in(a10_wr[823]),  .coef_in(coef[0]), .rdup_out(a11_wr[822]), .rdlo_out(a11_wr[823]));
			radix2 #(.width(width)) rd_st10_824  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[824]), .rdlo_in(a10_wr[825]),  .coef_in(coef[0]), .rdup_out(a11_wr[824]), .rdlo_out(a11_wr[825]));
			radix2 #(.width(width)) rd_st10_826  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[826]), .rdlo_in(a10_wr[827]),  .coef_in(coef[0]), .rdup_out(a11_wr[826]), .rdlo_out(a11_wr[827]));
			radix2 #(.width(width)) rd_st10_828  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[828]), .rdlo_in(a10_wr[829]),  .coef_in(coef[0]), .rdup_out(a11_wr[828]), .rdlo_out(a11_wr[829]));
			radix2 #(.width(width)) rd_st10_830  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[830]), .rdlo_in(a10_wr[831]),  .coef_in(coef[0]), .rdup_out(a11_wr[830]), .rdlo_out(a11_wr[831]));
			radix2 #(.width(width)) rd_st10_832  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[832]), .rdlo_in(a10_wr[833]),  .coef_in(coef[0]), .rdup_out(a11_wr[832]), .rdlo_out(a11_wr[833]));
			radix2 #(.width(width)) rd_st10_834  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[834]), .rdlo_in(a10_wr[835]),  .coef_in(coef[0]), .rdup_out(a11_wr[834]), .rdlo_out(a11_wr[835]));
			radix2 #(.width(width)) rd_st10_836  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[836]), .rdlo_in(a10_wr[837]),  .coef_in(coef[0]), .rdup_out(a11_wr[836]), .rdlo_out(a11_wr[837]));
			radix2 #(.width(width)) rd_st10_838  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[838]), .rdlo_in(a10_wr[839]),  .coef_in(coef[0]), .rdup_out(a11_wr[838]), .rdlo_out(a11_wr[839]));
			radix2 #(.width(width)) rd_st10_840  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[840]), .rdlo_in(a10_wr[841]),  .coef_in(coef[0]), .rdup_out(a11_wr[840]), .rdlo_out(a11_wr[841]));
			radix2 #(.width(width)) rd_st10_842  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[842]), .rdlo_in(a10_wr[843]),  .coef_in(coef[0]), .rdup_out(a11_wr[842]), .rdlo_out(a11_wr[843]));
			radix2 #(.width(width)) rd_st10_844  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[844]), .rdlo_in(a10_wr[845]),  .coef_in(coef[0]), .rdup_out(a11_wr[844]), .rdlo_out(a11_wr[845]));
			radix2 #(.width(width)) rd_st10_846  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[846]), .rdlo_in(a10_wr[847]),  .coef_in(coef[0]), .rdup_out(a11_wr[846]), .rdlo_out(a11_wr[847]));
			radix2 #(.width(width)) rd_st10_848  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[848]), .rdlo_in(a10_wr[849]),  .coef_in(coef[0]), .rdup_out(a11_wr[848]), .rdlo_out(a11_wr[849]));
			radix2 #(.width(width)) rd_st10_850  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[850]), .rdlo_in(a10_wr[851]),  .coef_in(coef[0]), .rdup_out(a11_wr[850]), .rdlo_out(a11_wr[851]));
			radix2 #(.width(width)) rd_st10_852  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[852]), .rdlo_in(a10_wr[853]),  .coef_in(coef[0]), .rdup_out(a11_wr[852]), .rdlo_out(a11_wr[853]));
			radix2 #(.width(width)) rd_st10_854  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[854]), .rdlo_in(a10_wr[855]),  .coef_in(coef[0]), .rdup_out(a11_wr[854]), .rdlo_out(a11_wr[855]));
			radix2 #(.width(width)) rd_st10_856  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[856]), .rdlo_in(a10_wr[857]),  .coef_in(coef[0]), .rdup_out(a11_wr[856]), .rdlo_out(a11_wr[857]));
			radix2 #(.width(width)) rd_st10_858  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[858]), .rdlo_in(a10_wr[859]),  .coef_in(coef[0]), .rdup_out(a11_wr[858]), .rdlo_out(a11_wr[859]));
			radix2 #(.width(width)) rd_st10_860  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[860]), .rdlo_in(a10_wr[861]),  .coef_in(coef[0]), .rdup_out(a11_wr[860]), .rdlo_out(a11_wr[861]));
			radix2 #(.width(width)) rd_st10_862  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[862]), .rdlo_in(a10_wr[863]),  .coef_in(coef[0]), .rdup_out(a11_wr[862]), .rdlo_out(a11_wr[863]));
			radix2 #(.width(width)) rd_st10_864  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[864]), .rdlo_in(a10_wr[865]),  .coef_in(coef[0]), .rdup_out(a11_wr[864]), .rdlo_out(a11_wr[865]));
			radix2 #(.width(width)) rd_st10_866  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[866]), .rdlo_in(a10_wr[867]),  .coef_in(coef[0]), .rdup_out(a11_wr[866]), .rdlo_out(a11_wr[867]));
			radix2 #(.width(width)) rd_st10_868  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[868]), .rdlo_in(a10_wr[869]),  .coef_in(coef[0]), .rdup_out(a11_wr[868]), .rdlo_out(a11_wr[869]));
			radix2 #(.width(width)) rd_st10_870  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[870]), .rdlo_in(a10_wr[871]),  .coef_in(coef[0]), .rdup_out(a11_wr[870]), .rdlo_out(a11_wr[871]));
			radix2 #(.width(width)) rd_st10_872  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[872]), .rdlo_in(a10_wr[873]),  .coef_in(coef[0]), .rdup_out(a11_wr[872]), .rdlo_out(a11_wr[873]));
			radix2 #(.width(width)) rd_st10_874  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[874]), .rdlo_in(a10_wr[875]),  .coef_in(coef[0]), .rdup_out(a11_wr[874]), .rdlo_out(a11_wr[875]));
			radix2 #(.width(width)) rd_st10_876  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[876]), .rdlo_in(a10_wr[877]),  .coef_in(coef[0]), .rdup_out(a11_wr[876]), .rdlo_out(a11_wr[877]));
			radix2 #(.width(width)) rd_st10_878  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[878]), .rdlo_in(a10_wr[879]),  .coef_in(coef[0]), .rdup_out(a11_wr[878]), .rdlo_out(a11_wr[879]));
			radix2 #(.width(width)) rd_st10_880  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[880]), .rdlo_in(a10_wr[881]),  .coef_in(coef[0]), .rdup_out(a11_wr[880]), .rdlo_out(a11_wr[881]));
			radix2 #(.width(width)) rd_st10_882  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[882]), .rdlo_in(a10_wr[883]),  .coef_in(coef[0]), .rdup_out(a11_wr[882]), .rdlo_out(a11_wr[883]));
			radix2 #(.width(width)) rd_st10_884  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[884]), .rdlo_in(a10_wr[885]),  .coef_in(coef[0]), .rdup_out(a11_wr[884]), .rdlo_out(a11_wr[885]));
			radix2 #(.width(width)) rd_st10_886  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[886]), .rdlo_in(a10_wr[887]),  .coef_in(coef[0]), .rdup_out(a11_wr[886]), .rdlo_out(a11_wr[887]));
			radix2 #(.width(width)) rd_st10_888  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[888]), .rdlo_in(a10_wr[889]),  .coef_in(coef[0]), .rdup_out(a11_wr[888]), .rdlo_out(a11_wr[889]));
			radix2 #(.width(width)) rd_st10_890  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[890]), .rdlo_in(a10_wr[891]),  .coef_in(coef[0]), .rdup_out(a11_wr[890]), .rdlo_out(a11_wr[891]));
			radix2 #(.width(width)) rd_st10_892  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[892]), .rdlo_in(a10_wr[893]),  .coef_in(coef[0]), .rdup_out(a11_wr[892]), .rdlo_out(a11_wr[893]));
			radix2 #(.width(width)) rd_st10_894  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[894]), .rdlo_in(a10_wr[895]),  .coef_in(coef[0]), .rdup_out(a11_wr[894]), .rdlo_out(a11_wr[895]));
			radix2 #(.width(width)) rd_st10_896  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[896]), .rdlo_in(a10_wr[897]),  .coef_in(coef[0]), .rdup_out(a11_wr[896]), .rdlo_out(a11_wr[897]));
			radix2 #(.width(width)) rd_st10_898  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[898]), .rdlo_in(a10_wr[899]),  .coef_in(coef[0]), .rdup_out(a11_wr[898]), .rdlo_out(a11_wr[899]));
			radix2 #(.width(width)) rd_st10_900  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[900]), .rdlo_in(a10_wr[901]),  .coef_in(coef[0]), .rdup_out(a11_wr[900]), .rdlo_out(a11_wr[901]));
			radix2 #(.width(width)) rd_st10_902  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[902]), .rdlo_in(a10_wr[903]),  .coef_in(coef[0]), .rdup_out(a11_wr[902]), .rdlo_out(a11_wr[903]));
			radix2 #(.width(width)) rd_st10_904  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[904]), .rdlo_in(a10_wr[905]),  .coef_in(coef[0]), .rdup_out(a11_wr[904]), .rdlo_out(a11_wr[905]));
			radix2 #(.width(width)) rd_st10_906  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[906]), .rdlo_in(a10_wr[907]),  .coef_in(coef[0]), .rdup_out(a11_wr[906]), .rdlo_out(a11_wr[907]));
			radix2 #(.width(width)) rd_st10_908  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[908]), .rdlo_in(a10_wr[909]),  .coef_in(coef[0]), .rdup_out(a11_wr[908]), .rdlo_out(a11_wr[909]));
			radix2 #(.width(width)) rd_st10_910  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[910]), .rdlo_in(a10_wr[911]),  .coef_in(coef[0]), .rdup_out(a11_wr[910]), .rdlo_out(a11_wr[911]));
			radix2 #(.width(width)) rd_st10_912  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[912]), .rdlo_in(a10_wr[913]),  .coef_in(coef[0]), .rdup_out(a11_wr[912]), .rdlo_out(a11_wr[913]));
			radix2 #(.width(width)) rd_st10_914  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[914]), .rdlo_in(a10_wr[915]),  .coef_in(coef[0]), .rdup_out(a11_wr[914]), .rdlo_out(a11_wr[915]));
			radix2 #(.width(width)) rd_st10_916  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[916]), .rdlo_in(a10_wr[917]),  .coef_in(coef[0]), .rdup_out(a11_wr[916]), .rdlo_out(a11_wr[917]));
			radix2 #(.width(width)) rd_st10_918  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[918]), .rdlo_in(a10_wr[919]),  .coef_in(coef[0]), .rdup_out(a11_wr[918]), .rdlo_out(a11_wr[919]));
			radix2 #(.width(width)) rd_st10_920  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[920]), .rdlo_in(a10_wr[921]),  .coef_in(coef[0]), .rdup_out(a11_wr[920]), .rdlo_out(a11_wr[921]));
			radix2 #(.width(width)) rd_st10_922  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[922]), .rdlo_in(a10_wr[923]),  .coef_in(coef[0]), .rdup_out(a11_wr[922]), .rdlo_out(a11_wr[923]));
			radix2 #(.width(width)) rd_st10_924  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[924]), .rdlo_in(a10_wr[925]),  .coef_in(coef[0]), .rdup_out(a11_wr[924]), .rdlo_out(a11_wr[925]));
			radix2 #(.width(width)) rd_st10_926  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[926]), .rdlo_in(a10_wr[927]),  .coef_in(coef[0]), .rdup_out(a11_wr[926]), .rdlo_out(a11_wr[927]));
			radix2 #(.width(width)) rd_st10_928  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[928]), .rdlo_in(a10_wr[929]),  .coef_in(coef[0]), .rdup_out(a11_wr[928]), .rdlo_out(a11_wr[929]));
			radix2 #(.width(width)) rd_st10_930  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[930]), .rdlo_in(a10_wr[931]),  .coef_in(coef[0]), .rdup_out(a11_wr[930]), .rdlo_out(a11_wr[931]));
			radix2 #(.width(width)) rd_st10_932  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[932]), .rdlo_in(a10_wr[933]),  .coef_in(coef[0]), .rdup_out(a11_wr[932]), .rdlo_out(a11_wr[933]));
			radix2 #(.width(width)) rd_st10_934  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[934]), .rdlo_in(a10_wr[935]),  .coef_in(coef[0]), .rdup_out(a11_wr[934]), .rdlo_out(a11_wr[935]));
			radix2 #(.width(width)) rd_st10_936  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[936]), .rdlo_in(a10_wr[937]),  .coef_in(coef[0]), .rdup_out(a11_wr[936]), .rdlo_out(a11_wr[937]));
			radix2 #(.width(width)) rd_st10_938  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[938]), .rdlo_in(a10_wr[939]),  .coef_in(coef[0]), .rdup_out(a11_wr[938]), .rdlo_out(a11_wr[939]));
			radix2 #(.width(width)) rd_st10_940  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[940]), .rdlo_in(a10_wr[941]),  .coef_in(coef[0]), .rdup_out(a11_wr[940]), .rdlo_out(a11_wr[941]));
			radix2 #(.width(width)) rd_st10_942  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[942]), .rdlo_in(a10_wr[943]),  .coef_in(coef[0]), .rdup_out(a11_wr[942]), .rdlo_out(a11_wr[943]));
			radix2 #(.width(width)) rd_st10_944  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[944]), .rdlo_in(a10_wr[945]),  .coef_in(coef[0]), .rdup_out(a11_wr[944]), .rdlo_out(a11_wr[945]));
			radix2 #(.width(width)) rd_st10_946  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[946]), .rdlo_in(a10_wr[947]),  .coef_in(coef[0]), .rdup_out(a11_wr[946]), .rdlo_out(a11_wr[947]));
			radix2 #(.width(width)) rd_st10_948  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[948]), .rdlo_in(a10_wr[949]),  .coef_in(coef[0]), .rdup_out(a11_wr[948]), .rdlo_out(a11_wr[949]));
			radix2 #(.width(width)) rd_st10_950  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[950]), .rdlo_in(a10_wr[951]),  .coef_in(coef[0]), .rdup_out(a11_wr[950]), .rdlo_out(a11_wr[951]));
			radix2 #(.width(width)) rd_st10_952  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[952]), .rdlo_in(a10_wr[953]),  .coef_in(coef[0]), .rdup_out(a11_wr[952]), .rdlo_out(a11_wr[953]));
			radix2 #(.width(width)) rd_st10_954  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[954]), .rdlo_in(a10_wr[955]),  .coef_in(coef[0]), .rdup_out(a11_wr[954]), .rdlo_out(a11_wr[955]));
			radix2 #(.width(width)) rd_st10_956  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[956]), .rdlo_in(a10_wr[957]),  .coef_in(coef[0]), .rdup_out(a11_wr[956]), .rdlo_out(a11_wr[957]));
			radix2 #(.width(width)) rd_st10_958  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[958]), .rdlo_in(a10_wr[959]),  .coef_in(coef[0]), .rdup_out(a11_wr[958]), .rdlo_out(a11_wr[959]));
			radix2 #(.width(width)) rd_st10_960  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[960]), .rdlo_in(a10_wr[961]),  .coef_in(coef[0]), .rdup_out(a11_wr[960]), .rdlo_out(a11_wr[961]));
			radix2 #(.width(width)) rd_st10_962  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[962]), .rdlo_in(a10_wr[963]),  .coef_in(coef[0]), .rdup_out(a11_wr[962]), .rdlo_out(a11_wr[963]));
			radix2 #(.width(width)) rd_st10_964  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[964]), .rdlo_in(a10_wr[965]),  .coef_in(coef[0]), .rdup_out(a11_wr[964]), .rdlo_out(a11_wr[965]));
			radix2 #(.width(width)) rd_st10_966  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[966]), .rdlo_in(a10_wr[967]),  .coef_in(coef[0]), .rdup_out(a11_wr[966]), .rdlo_out(a11_wr[967]));
			radix2 #(.width(width)) rd_st10_968  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[968]), .rdlo_in(a10_wr[969]),  .coef_in(coef[0]), .rdup_out(a11_wr[968]), .rdlo_out(a11_wr[969]));
			radix2 #(.width(width)) rd_st10_970  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[970]), .rdlo_in(a10_wr[971]),  .coef_in(coef[0]), .rdup_out(a11_wr[970]), .rdlo_out(a11_wr[971]));
			radix2 #(.width(width)) rd_st10_972  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[972]), .rdlo_in(a10_wr[973]),  .coef_in(coef[0]), .rdup_out(a11_wr[972]), .rdlo_out(a11_wr[973]));
			radix2 #(.width(width)) rd_st10_974  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[974]), .rdlo_in(a10_wr[975]),  .coef_in(coef[0]), .rdup_out(a11_wr[974]), .rdlo_out(a11_wr[975]));
			radix2 #(.width(width)) rd_st10_976  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[976]), .rdlo_in(a10_wr[977]),  .coef_in(coef[0]), .rdup_out(a11_wr[976]), .rdlo_out(a11_wr[977]));
			radix2 #(.width(width)) rd_st10_978  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[978]), .rdlo_in(a10_wr[979]),  .coef_in(coef[0]), .rdup_out(a11_wr[978]), .rdlo_out(a11_wr[979]));
			radix2 #(.width(width)) rd_st10_980  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[980]), .rdlo_in(a10_wr[981]),  .coef_in(coef[0]), .rdup_out(a11_wr[980]), .rdlo_out(a11_wr[981]));
			radix2 #(.width(width)) rd_st10_982  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[982]), .rdlo_in(a10_wr[983]),  .coef_in(coef[0]), .rdup_out(a11_wr[982]), .rdlo_out(a11_wr[983]));
			radix2 #(.width(width)) rd_st10_984  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[984]), .rdlo_in(a10_wr[985]),  .coef_in(coef[0]), .rdup_out(a11_wr[984]), .rdlo_out(a11_wr[985]));
			radix2 #(.width(width)) rd_st10_986  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[986]), .rdlo_in(a10_wr[987]),  .coef_in(coef[0]), .rdup_out(a11_wr[986]), .rdlo_out(a11_wr[987]));
			radix2 #(.width(width)) rd_st10_988  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[988]), .rdlo_in(a10_wr[989]),  .coef_in(coef[0]), .rdup_out(a11_wr[988]), .rdlo_out(a11_wr[989]));
			radix2 #(.width(width)) rd_st10_990  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[990]), .rdlo_in(a10_wr[991]),  .coef_in(coef[0]), .rdup_out(a11_wr[990]), .rdlo_out(a11_wr[991]));
			radix2 #(.width(width)) rd_st10_992  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[992]), .rdlo_in(a10_wr[993]),  .coef_in(coef[0]), .rdup_out(a11_wr[992]), .rdlo_out(a11_wr[993]));
			radix2 #(.width(width)) rd_st10_994  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[994]), .rdlo_in(a10_wr[995]),  .coef_in(coef[0]), .rdup_out(a11_wr[994]), .rdlo_out(a11_wr[995]));
			radix2 #(.width(width)) rd_st10_996  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[996]), .rdlo_in(a10_wr[997]),  .coef_in(coef[0]), .rdup_out(a11_wr[996]), .rdlo_out(a11_wr[997]));
			radix2 #(.width(width)) rd_st10_998  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[998]), .rdlo_in(a10_wr[999]),  .coef_in(coef[0]), .rdup_out(a11_wr[998]), .rdlo_out(a11_wr[999]));
			radix2 #(.width(width)) rd_st10_1000  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1000]), .rdlo_in(a10_wr[1001]),  .coef_in(coef[0]), .rdup_out(a11_wr[1000]), .rdlo_out(a11_wr[1001]));
			radix2 #(.width(width)) rd_st10_1002  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1002]), .rdlo_in(a10_wr[1003]),  .coef_in(coef[0]), .rdup_out(a11_wr[1002]), .rdlo_out(a11_wr[1003]));
			radix2 #(.width(width)) rd_st10_1004  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1004]), .rdlo_in(a10_wr[1005]),  .coef_in(coef[0]), .rdup_out(a11_wr[1004]), .rdlo_out(a11_wr[1005]));
			radix2 #(.width(width)) rd_st10_1006  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1006]), .rdlo_in(a10_wr[1007]),  .coef_in(coef[0]), .rdup_out(a11_wr[1006]), .rdlo_out(a11_wr[1007]));
			radix2 #(.width(width)) rd_st10_1008  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1008]), .rdlo_in(a10_wr[1009]),  .coef_in(coef[0]), .rdup_out(a11_wr[1008]), .rdlo_out(a11_wr[1009]));
			radix2 #(.width(width)) rd_st10_1010  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1010]), .rdlo_in(a10_wr[1011]),  .coef_in(coef[0]), .rdup_out(a11_wr[1010]), .rdlo_out(a11_wr[1011]));
			radix2 #(.width(width)) rd_st10_1012  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1012]), .rdlo_in(a10_wr[1013]),  .coef_in(coef[0]), .rdup_out(a11_wr[1012]), .rdlo_out(a11_wr[1013]));
			radix2 #(.width(width)) rd_st10_1014  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1014]), .rdlo_in(a10_wr[1015]),  .coef_in(coef[0]), .rdup_out(a11_wr[1014]), .rdlo_out(a11_wr[1015]));
			radix2 #(.width(width)) rd_st10_1016  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1016]), .rdlo_in(a10_wr[1017]),  .coef_in(coef[0]), .rdup_out(a11_wr[1016]), .rdlo_out(a11_wr[1017]));
			radix2 #(.width(width)) rd_st10_1018  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1018]), .rdlo_in(a10_wr[1019]),  .coef_in(coef[0]), .rdup_out(a11_wr[1018]), .rdlo_out(a11_wr[1019]));
			radix2 #(.width(width)) rd_st10_1020  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1020]), .rdlo_in(a10_wr[1021]),  .coef_in(coef[0]), .rdup_out(a11_wr[1020]), .rdlo_out(a11_wr[1021]));
			radix2 #(.width(width)) rd_st10_1022  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1022]), .rdlo_in(a10_wr[1023]),  .coef_in(coef[0]), .rdup_out(a11_wr[1022]), .rdlo_out(a11_wr[1023]));
			radix2 #(.width(width)) rd_st10_1024  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1024]), .rdlo_in(a10_wr[1025]),  .coef_in(coef[0]), .rdup_out(a11_wr[1024]), .rdlo_out(a11_wr[1025]));
			radix2 #(.width(width)) rd_st10_1026  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1026]), .rdlo_in(a10_wr[1027]),  .coef_in(coef[0]), .rdup_out(a11_wr[1026]), .rdlo_out(a11_wr[1027]));
			radix2 #(.width(width)) rd_st10_1028  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1028]), .rdlo_in(a10_wr[1029]),  .coef_in(coef[0]), .rdup_out(a11_wr[1028]), .rdlo_out(a11_wr[1029]));
			radix2 #(.width(width)) rd_st10_1030  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1030]), .rdlo_in(a10_wr[1031]),  .coef_in(coef[0]), .rdup_out(a11_wr[1030]), .rdlo_out(a11_wr[1031]));
			radix2 #(.width(width)) rd_st10_1032  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1032]), .rdlo_in(a10_wr[1033]),  .coef_in(coef[0]), .rdup_out(a11_wr[1032]), .rdlo_out(a11_wr[1033]));
			radix2 #(.width(width)) rd_st10_1034  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1034]), .rdlo_in(a10_wr[1035]),  .coef_in(coef[0]), .rdup_out(a11_wr[1034]), .rdlo_out(a11_wr[1035]));
			radix2 #(.width(width)) rd_st10_1036  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1036]), .rdlo_in(a10_wr[1037]),  .coef_in(coef[0]), .rdup_out(a11_wr[1036]), .rdlo_out(a11_wr[1037]));
			radix2 #(.width(width)) rd_st10_1038  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1038]), .rdlo_in(a10_wr[1039]),  .coef_in(coef[0]), .rdup_out(a11_wr[1038]), .rdlo_out(a11_wr[1039]));
			radix2 #(.width(width)) rd_st10_1040  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1040]), .rdlo_in(a10_wr[1041]),  .coef_in(coef[0]), .rdup_out(a11_wr[1040]), .rdlo_out(a11_wr[1041]));
			radix2 #(.width(width)) rd_st10_1042  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1042]), .rdlo_in(a10_wr[1043]),  .coef_in(coef[0]), .rdup_out(a11_wr[1042]), .rdlo_out(a11_wr[1043]));
			radix2 #(.width(width)) rd_st10_1044  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1044]), .rdlo_in(a10_wr[1045]),  .coef_in(coef[0]), .rdup_out(a11_wr[1044]), .rdlo_out(a11_wr[1045]));
			radix2 #(.width(width)) rd_st10_1046  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1046]), .rdlo_in(a10_wr[1047]),  .coef_in(coef[0]), .rdup_out(a11_wr[1046]), .rdlo_out(a11_wr[1047]));
			radix2 #(.width(width)) rd_st10_1048  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1048]), .rdlo_in(a10_wr[1049]),  .coef_in(coef[0]), .rdup_out(a11_wr[1048]), .rdlo_out(a11_wr[1049]));
			radix2 #(.width(width)) rd_st10_1050  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1050]), .rdlo_in(a10_wr[1051]),  .coef_in(coef[0]), .rdup_out(a11_wr[1050]), .rdlo_out(a11_wr[1051]));
			radix2 #(.width(width)) rd_st10_1052  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1052]), .rdlo_in(a10_wr[1053]),  .coef_in(coef[0]), .rdup_out(a11_wr[1052]), .rdlo_out(a11_wr[1053]));
			radix2 #(.width(width)) rd_st10_1054  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1054]), .rdlo_in(a10_wr[1055]),  .coef_in(coef[0]), .rdup_out(a11_wr[1054]), .rdlo_out(a11_wr[1055]));
			radix2 #(.width(width)) rd_st10_1056  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1056]), .rdlo_in(a10_wr[1057]),  .coef_in(coef[0]), .rdup_out(a11_wr[1056]), .rdlo_out(a11_wr[1057]));
			radix2 #(.width(width)) rd_st10_1058  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1058]), .rdlo_in(a10_wr[1059]),  .coef_in(coef[0]), .rdup_out(a11_wr[1058]), .rdlo_out(a11_wr[1059]));
			radix2 #(.width(width)) rd_st10_1060  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1060]), .rdlo_in(a10_wr[1061]),  .coef_in(coef[0]), .rdup_out(a11_wr[1060]), .rdlo_out(a11_wr[1061]));
			radix2 #(.width(width)) rd_st10_1062  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1062]), .rdlo_in(a10_wr[1063]),  .coef_in(coef[0]), .rdup_out(a11_wr[1062]), .rdlo_out(a11_wr[1063]));
			radix2 #(.width(width)) rd_st10_1064  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1064]), .rdlo_in(a10_wr[1065]),  .coef_in(coef[0]), .rdup_out(a11_wr[1064]), .rdlo_out(a11_wr[1065]));
			radix2 #(.width(width)) rd_st10_1066  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1066]), .rdlo_in(a10_wr[1067]),  .coef_in(coef[0]), .rdup_out(a11_wr[1066]), .rdlo_out(a11_wr[1067]));
			radix2 #(.width(width)) rd_st10_1068  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1068]), .rdlo_in(a10_wr[1069]),  .coef_in(coef[0]), .rdup_out(a11_wr[1068]), .rdlo_out(a11_wr[1069]));
			radix2 #(.width(width)) rd_st10_1070  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1070]), .rdlo_in(a10_wr[1071]),  .coef_in(coef[0]), .rdup_out(a11_wr[1070]), .rdlo_out(a11_wr[1071]));
			radix2 #(.width(width)) rd_st10_1072  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1072]), .rdlo_in(a10_wr[1073]),  .coef_in(coef[0]), .rdup_out(a11_wr[1072]), .rdlo_out(a11_wr[1073]));
			radix2 #(.width(width)) rd_st10_1074  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1074]), .rdlo_in(a10_wr[1075]),  .coef_in(coef[0]), .rdup_out(a11_wr[1074]), .rdlo_out(a11_wr[1075]));
			radix2 #(.width(width)) rd_st10_1076  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1076]), .rdlo_in(a10_wr[1077]),  .coef_in(coef[0]), .rdup_out(a11_wr[1076]), .rdlo_out(a11_wr[1077]));
			radix2 #(.width(width)) rd_st10_1078  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1078]), .rdlo_in(a10_wr[1079]),  .coef_in(coef[0]), .rdup_out(a11_wr[1078]), .rdlo_out(a11_wr[1079]));
			radix2 #(.width(width)) rd_st10_1080  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1080]), .rdlo_in(a10_wr[1081]),  .coef_in(coef[0]), .rdup_out(a11_wr[1080]), .rdlo_out(a11_wr[1081]));
			radix2 #(.width(width)) rd_st10_1082  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1082]), .rdlo_in(a10_wr[1083]),  .coef_in(coef[0]), .rdup_out(a11_wr[1082]), .rdlo_out(a11_wr[1083]));
			radix2 #(.width(width)) rd_st10_1084  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1084]), .rdlo_in(a10_wr[1085]),  .coef_in(coef[0]), .rdup_out(a11_wr[1084]), .rdlo_out(a11_wr[1085]));
			radix2 #(.width(width)) rd_st10_1086  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1086]), .rdlo_in(a10_wr[1087]),  .coef_in(coef[0]), .rdup_out(a11_wr[1086]), .rdlo_out(a11_wr[1087]));
			radix2 #(.width(width)) rd_st10_1088  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1088]), .rdlo_in(a10_wr[1089]),  .coef_in(coef[0]), .rdup_out(a11_wr[1088]), .rdlo_out(a11_wr[1089]));
			radix2 #(.width(width)) rd_st10_1090  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1090]), .rdlo_in(a10_wr[1091]),  .coef_in(coef[0]), .rdup_out(a11_wr[1090]), .rdlo_out(a11_wr[1091]));
			radix2 #(.width(width)) rd_st10_1092  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1092]), .rdlo_in(a10_wr[1093]),  .coef_in(coef[0]), .rdup_out(a11_wr[1092]), .rdlo_out(a11_wr[1093]));
			radix2 #(.width(width)) rd_st10_1094  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1094]), .rdlo_in(a10_wr[1095]),  .coef_in(coef[0]), .rdup_out(a11_wr[1094]), .rdlo_out(a11_wr[1095]));
			radix2 #(.width(width)) rd_st10_1096  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1096]), .rdlo_in(a10_wr[1097]),  .coef_in(coef[0]), .rdup_out(a11_wr[1096]), .rdlo_out(a11_wr[1097]));
			radix2 #(.width(width)) rd_st10_1098  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1098]), .rdlo_in(a10_wr[1099]),  .coef_in(coef[0]), .rdup_out(a11_wr[1098]), .rdlo_out(a11_wr[1099]));
			radix2 #(.width(width)) rd_st10_1100  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1100]), .rdlo_in(a10_wr[1101]),  .coef_in(coef[0]), .rdup_out(a11_wr[1100]), .rdlo_out(a11_wr[1101]));
			radix2 #(.width(width)) rd_st10_1102  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1102]), .rdlo_in(a10_wr[1103]),  .coef_in(coef[0]), .rdup_out(a11_wr[1102]), .rdlo_out(a11_wr[1103]));
			radix2 #(.width(width)) rd_st10_1104  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1104]), .rdlo_in(a10_wr[1105]),  .coef_in(coef[0]), .rdup_out(a11_wr[1104]), .rdlo_out(a11_wr[1105]));
			radix2 #(.width(width)) rd_st10_1106  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1106]), .rdlo_in(a10_wr[1107]),  .coef_in(coef[0]), .rdup_out(a11_wr[1106]), .rdlo_out(a11_wr[1107]));
			radix2 #(.width(width)) rd_st10_1108  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1108]), .rdlo_in(a10_wr[1109]),  .coef_in(coef[0]), .rdup_out(a11_wr[1108]), .rdlo_out(a11_wr[1109]));
			radix2 #(.width(width)) rd_st10_1110  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1110]), .rdlo_in(a10_wr[1111]),  .coef_in(coef[0]), .rdup_out(a11_wr[1110]), .rdlo_out(a11_wr[1111]));
			radix2 #(.width(width)) rd_st10_1112  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1112]), .rdlo_in(a10_wr[1113]),  .coef_in(coef[0]), .rdup_out(a11_wr[1112]), .rdlo_out(a11_wr[1113]));
			radix2 #(.width(width)) rd_st10_1114  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1114]), .rdlo_in(a10_wr[1115]),  .coef_in(coef[0]), .rdup_out(a11_wr[1114]), .rdlo_out(a11_wr[1115]));
			radix2 #(.width(width)) rd_st10_1116  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1116]), .rdlo_in(a10_wr[1117]),  .coef_in(coef[0]), .rdup_out(a11_wr[1116]), .rdlo_out(a11_wr[1117]));
			radix2 #(.width(width)) rd_st10_1118  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1118]), .rdlo_in(a10_wr[1119]),  .coef_in(coef[0]), .rdup_out(a11_wr[1118]), .rdlo_out(a11_wr[1119]));
			radix2 #(.width(width)) rd_st10_1120  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1120]), .rdlo_in(a10_wr[1121]),  .coef_in(coef[0]), .rdup_out(a11_wr[1120]), .rdlo_out(a11_wr[1121]));
			radix2 #(.width(width)) rd_st10_1122  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1122]), .rdlo_in(a10_wr[1123]),  .coef_in(coef[0]), .rdup_out(a11_wr[1122]), .rdlo_out(a11_wr[1123]));
			radix2 #(.width(width)) rd_st10_1124  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1124]), .rdlo_in(a10_wr[1125]),  .coef_in(coef[0]), .rdup_out(a11_wr[1124]), .rdlo_out(a11_wr[1125]));
			radix2 #(.width(width)) rd_st10_1126  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1126]), .rdlo_in(a10_wr[1127]),  .coef_in(coef[0]), .rdup_out(a11_wr[1126]), .rdlo_out(a11_wr[1127]));
			radix2 #(.width(width)) rd_st10_1128  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1128]), .rdlo_in(a10_wr[1129]),  .coef_in(coef[0]), .rdup_out(a11_wr[1128]), .rdlo_out(a11_wr[1129]));
			radix2 #(.width(width)) rd_st10_1130  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1130]), .rdlo_in(a10_wr[1131]),  .coef_in(coef[0]), .rdup_out(a11_wr[1130]), .rdlo_out(a11_wr[1131]));
			radix2 #(.width(width)) rd_st10_1132  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1132]), .rdlo_in(a10_wr[1133]),  .coef_in(coef[0]), .rdup_out(a11_wr[1132]), .rdlo_out(a11_wr[1133]));
			radix2 #(.width(width)) rd_st10_1134  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1134]), .rdlo_in(a10_wr[1135]),  .coef_in(coef[0]), .rdup_out(a11_wr[1134]), .rdlo_out(a11_wr[1135]));
			radix2 #(.width(width)) rd_st10_1136  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1136]), .rdlo_in(a10_wr[1137]),  .coef_in(coef[0]), .rdup_out(a11_wr[1136]), .rdlo_out(a11_wr[1137]));
			radix2 #(.width(width)) rd_st10_1138  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1138]), .rdlo_in(a10_wr[1139]),  .coef_in(coef[0]), .rdup_out(a11_wr[1138]), .rdlo_out(a11_wr[1139]));
			radix2 #(.width(width)) rd_st10_1140  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1140]), .rdlo_in(a10_wr[1141]),  .coef_in(coef[0]), .rdup_out(a11_wr[1140]), .rdlo_out(a11_wr[1141]));
			radix2 #(.width(width)) rd_st10_1142  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1142]), .rdlo_in(a10_wr[1143]),  .coef_in(coef[0]), .rdup_out(a11_wr[1142]), .rdlo_out(a11_wr[1143]));
			radix2 #(.width(width)) rd_st10_1144  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1144]), .rdlo_in(a10_wr[1145]),  .coef_in(coef[0]), .rdup_out(a11_wr[1144]), .rdlo_out(a11_wr[1145]));
			radix2 #(.width(width)) rd_st10_1146  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1146]), .rdlo_in(a10_wr[1147]),  .coef_in(coef[0]), .rdup_out(a11_wr[1146]), .rdlo_out(a11_wr[1147]));
			radix2 #(.width(width)) rd_st10_1148  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1148]), .rdlo_in(a10_wr[1149]),  .coef_in(coef[0]), .rdup_out(a11_wr[1148]), .rdlo_out(a11_wr[1149]));
			radix2 #(.width(width)) rd_st10_1150  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1150]), .rdlo_in(a10_wr[1151]),  .coef_in(coef[0]), .rdup_out(a11_wr[1150]), .rdlo_out(a11_wr[1151]));
			radix2 #(.width(width)) rd_st10_1152  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1152]), .rdlo_in(a10_wr[1153]),  .coef_in(coef[0]), .rdup_out(a11_wr[1152]), .rdlo_out(a11_wr[1153]));
			radix2 #(.width(width)) rd_st10_1154  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1154]), .rdlo_in(a10_wr[1155]),  .coef_in(coef[0]), .rdup_out(a11_wr[1154]), .rdlo_out(a11_wr[1155]));
			radix2 #(.width(width)) rd_st10_1156  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1156]), .rdlo_in(a10_wr[1157]),  .coef_in(coef[0]), .rdup_out(a11_wr[1156]), .rdlo_out(a11_wr[1157]));
			radix2 #(.width(width)) rd_st10_1158  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1158]), .rdlo_in(a10_wr[1159]),  .coef_in(coef[0]), .rdup_out(a11_wr[1158]), .rdlo_out(a11_wr[1159]));
			radix2 #(.width(width)) rd_st10_1160  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1160]), .rdlo_in(a10_wr[1161]),  .coef_in(coef[0]), .rdup_out(a11_wr[1160]), .rdlo_out(a11_wr[1161]));
			radix2 #(.width(width)) rd_st10_1162  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1162]), .rdlo_in(a10_wr[1163]),  .coef_in(coef[0]), .rdup_out(a11_wr[1162]), .rdlo_out(a11_wr[1163]));
			radix2 #(.width(width)) rd_st10_1164  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1164]), .rdlo_in(a10_wr[1165]),  .coef_in(coef[0]), .rdup_out(a11_wr[1164]), .rdlo_out(a11_wr[1165]));
			radix2 #(.width(width)) rd_st10_1166  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1166]), .rdlo_in(a10_wr[1167]),  .coef_in(coef[0]), .rdup_out(a11_wr[1166]), .rdlo_out(a11_wr[1167]));
			radix2 #(.width(width)) rd_st10_1168  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1168]), .rdlo_in(a10_wr[1169]),  .coef_in(coef[0]), .rdup_out(a11_wr[1168]), .rdlo_out(a11_wr[1169]));
			radix2 #(.width(width)) rd_st10_1170  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1170]), .rdlo_in(a10_wr[1171]),  .coef_in(coef[0]), .rdup_out(a11_wr[1170]), .rdlo_out(a11_wr[1171]));
			radix2 #(.width(width)) rd_st10_1172  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1172]), .rdlo_in(a10_wr[1173]),  .coef_in(coef[0]), .rdup_out(a11_wr[1172]), .rdlo_out(a11_wr[1173]));
			radix2 #(.width(width)) rd_st10_1174  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1174]), .rdlo_in(a10_wr[1175]),  .coef_in(coef[0]), .rdup_out(a11_wr[1174]), .rdlo_out(a11_wr[1175]));
			radix2 #(.width(width)) rd_st10_1176  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1176]), .rdlo_in(a10_wr[1177]),  .coef_in(coef[0]), .rdup_out(a11_wr[1176]), .rdlo_out(a11_wr[1177]));
			radix2 #(.width(width)) rd_st10_1178  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1178]), .rdlo_in(a10_wr[1179]),  .coef_in(coef[0]), .rdup_out(a11_wr[1178]), .rdlo_out(a11_wr[1179]));
			radix2 #(.width(width)) rd_st10_1180  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1180]), .rdlo_in(a10_wr[1181]),  .coef_in(coef[0]), .rdup_out(a11_wr[1180]), .rdlo_out(a11_wr[1181]));
			radix2 #(.width(width)) rd_st10_1182  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1182]), .rdlo_in(a10_wr[1183]),  .coef_in(coef[0]), .rdup_out(a11_wr[1182]), .rdlo_out(a11_wr[1183]));
			radix2 #(.width(width)) rd_st10_1184  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1184]), .rdlo_in(a10_wr[1185]),  .coef_in(coef[0]), .rdup_out(a11_wr[1184]), .rdlo_out(a11_wr[1185]));
			radix2 #(.width(width)) rd_st10_1186  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1186]), .rdlo_in(a10_wr[1187]),  .coef_in(coef[0]), .rdup_out(a11_wr[1186]), .rdlo_out(a11_wr[1187]));
			radix2 #(.width(width)) rd_st10_1188  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1188]), .rdlo_in(a10_wr[1189]),  .coef_in(coef[0]), .rdup_out(a11_wr[1188]), .rdlo_out(a11_wr[1189]));
			radix2 #(.width(width)) rd_st10_1190  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1190]), .rdlo_in(a10_wr[1191]),  .coef_in(coef[0]), .rdup_out(a11_wr[1190]), .rdlo_out(a11_wr[1191]));
			radix2 #(.width(width)) rd_st10_1192  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1192]), .rdlo_in(a10_wr[1193]),  .coef_in(coef[0]), .rdup_out(a11_wr[1192]), .rdlo_out(a11_wr[1193]));
			radix2 #(.width(width)) rd_st10_1194  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1194]), .rdlo_in(a10_wr[1195]),  .coef_in(coef[0]), .rdup_out(a11_wr[1194]), .rdlo_out(a11_wr[1195]));
			radix2 #(.width(width)) rd_st10_1196  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1196]), .rdlo_in(a10_wr[1197]),  .coef_in(coef[0]), .rdup_out(a11_wr[1196]), .rdlo_out(a11_wr[1197]));
			radix2 #(.width(width)) rd_st10_1198  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1198]), .rdlo_in(a10_wr[1199]),  .coef_in(coef[0]), .rdup_out(a11_wr[1198]), .rdlo_out(a11_wr[1199]));
			radix2 #(.width(width)) rd_st10_1200  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1200]), .rdlo_in(a10_wr[1201]),  .coef_in(coef[0]), .rdup_out(a11_wr[1200]), .rdlo_out(a11_wr[1201]));
			radix2 #(.width(width)) rd_st10_1202  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1202]), .rdlo_in(a10_wr[1203]),  .coef_in(coef[0]), .rdup_out(a11_wr[1202]), .rdlo_out(a11_wr[1203]));
			radix2 #(.width(width)) rd_st10_1204  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1204]), .rdlo_in(a10_wr[1205]),  .coef_in(coef[0]), .rdup_out(a11_wr[1204]), .rdlo_out(a11_wr[1205]));
			radix2 #(.width(width)) rd_st10_1206  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1206]), .rdlo_in(a10_wr[1207]),  .coef_in(coef[0]), .rdup_out(a11_wr[1206]), .rdlo_out(a11_wr[1207]));
			radix2 #(.width(width)) rd_st10_1208  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1208]), .rdlo_in(a10_wr[1209]),  .coef_in(coef[0]), .rdup_out(a11_wr[1208]), .rdlo_out(a11_wr[1209]));
			radix2 #(.width(width)) rd_st10_1210  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1210]), .rdlo_in(a10_wr[1211]),  .coef_in(coef[0]), .rdup_out(a11_wr[1210]), .rdlo_out(a11_wr[1211]));
			radix2 #(.width(width)) rd_st10_1212  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1212]), .rdlo_in(a10_wr[1213]),  .coef_in(coef[0]), .rdup_out(a11_wr[1212]), .rdlo_out(a11_wr[1213]));
			radix2 #(.width(width)) rd_st10_1214  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1214]), .rdlo_in(a10_wr[1215]),  .coef_in(coef[0]), .rdup_out(a11_wr[1214]), .rdlo_out(a11_wr[1215]));
			radix2 #(.width(width)) rd_st10_1216  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1216]), .rdlo_in(a10_wr[1217]),  .coef_in(coef[0]), .rdup_out(a11_wr[1216]), .rdlo_out(a11_wr[1217]));
			radix2 #(.width(width)) rd_st10_1218  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1218]), .rdlo_in(a10_wr[1219]),  .coef_in(coef[0]), .rdup_out(a11_wr[1218]), .rdlo_out(a11_wr[1219]));
			radix2 #(.width(width)) rd_st10_1220  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1220]), .rdlo_in(a10_wr[1221]),  .coef_in(coef[0]), .rdup_out(a11_wr[1220]), .rdlo_out(a11_wr[1221]));
			radix2 #(.width(width)) rd_st10_1222  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1222]), .rdlo_in(a10_wr[1223]),  .coef_in(coef[0]), .rdup_out(a11_wr[1222]), .rdlo_out(a11_wr[1223]));
			radix2 #(.width(width)) rd_st10_1224  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1224]), .rdlo_in(a10_wr[1225]),  .coef_in(coef[0]), .rdup_out(a11_wr[1224]), .rdlo_out(a11_wr[1225]));
			radix2 #(.width(width)) rd_st10_1226  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1226]), .rdlo_in(a10_wr[1227]),  .coef_in(coef[0]), .rdup_out(a11_wr[1226]), .rdlo_out(a11_wr[1227]));
			radix2 #(.width(width)) rd_st10_1228  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1228]), .rdlo_in(a10_wr[1229]),  .coef_in(coef[0]), .rdup_out(a11_wr[1228]), .rdlo_out(a11_wr[1229]));
			radix2 #(.width(width)) rd_st10_1230  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1230]), .rdlo_in(a10_wr[1231]),  .coef_in(coef[0]), .rdup_out(a11_wr[1230]), .rdlo_out(a11_wr[1231]));
			radix2 #(.width(width)) rd_st10_1232  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1232]), .rdlo_in(a10_wr[1233]),  .coef_in(coef[0]), .rdup_out(a11_wr[1232]), .rdlo_out(a11_wr[1233]));
			radix2 #(.width(width)) rd_st10_1234  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1234]), .rdlo_in(a10_wr[1235]),  .coef_in(coef[0]), .rdup_out(a11_wr[1234]), .rdlo_out(a11_wr[1235]));
			radix2 #(.width(width)) rd_st10_1236  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1236]), .rdlo_in(a10_wr[1237]),  .coef_in(coef[0]), .rdup_out(a11_wr[1236]), .rdlo_out(a11_wr[1237]));
			radix2 #(.width(width)) rd_st10_1238  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1238]), .rdlo_in(a10_wr[1239]),  .coef_in(coef[0]), .rdup_out(a11_wr[1238]), .rdlo_out(a11_wr[1239]));
			radix2 #(.width(width)) rd_st10_1240  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1240]), .rdlo_in(a10_wr[1241]),  .coef_in(coef[0]), .rdup_out(a11_wr[1240]), .rdlo_out(a11_wr[1241]));
			radix2 #(.width(width)) rd_st10_1242  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1242]), .rdlo_in(a10_wr[1243]),  .coef_in(coef[0]), .rdup_out(a11_wr[1242]), .rdlo_out(a11_wr[1243]));
			radix2 #(.width(width)) rd_st10_1244  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1244]), .rdlo_in(a10_wr[1245]),  .coef_in(coef[0]), .rdup_out(a11_wr[1244]), .rdlo_out(a11_wr[1245]));
			radix2 #(.width(width)) rd_st10_1246  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1246]), .rdlo_in(a10_wr[1247]),  .coef_in(coef[0]), .rdup_out(a11_wr[1246]), .rdlo_out(a11_wr[1247]));
			radix2 #(.width(width)) rd_st10_1248  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1248]), .rdlo_in(a10_wr[1249]),  .coef_in(coef[0]), .rdup_out(a11_wr[1248]), .rdlo_out(a11_wr[1249]));
			radix2 #(.width(width)) rd_st10_1250  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1250]), .rdlo_in(a10_wr[1251]),  .coef_in(coef[0]), .rdup_out(a11_wr[1250]), .rdlo_out(a11_wr[1251]));
			radix2 #(.width(width)) rd_st10_1252  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1252]), .rdlo_in(a10_wr[1253]),  .coef_in(coef[0]), .rdup_out(a11_wr[1252]), .rdlo_out(a11_wr[1253]));
			radix2 #(.width(width)) rd_st10_1254  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1254]), .rdlo_in(a10_wr[1255]),  .coef_in(coef[0]), .rdup_out(a11_wr[1254]), .rdlo_out(a11_wr[1255]));
			radix2 #(.width(width)) rd_st10_1256  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1256]), .rdlo_in(a10_wr[1257]),  .coef_in(coef[0]), .rdup_out(a11_wr[1256]), .rdlo_out(a11_wr[1257]));
			radix2 #(.width(width)) rd_st10_1258  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1258]), .rdlo_in(a10_wr[1259]),  .coef_in(coef[0]), .rdup_out(a11_wr[1258]), .rdlo_out(a11_wr[1259]));
			radix2 #(.width(width)) rd_st10_1260  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1260]), .rdlo_in(a10_wr[1261]),  .coef_in(coef[0]), .rdup_out(a11_wr[1260]), .rdlo_out(a11_wr[1261]));
			radix2 #(.width(width)) rd_st10_1262  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1262]), .rdlo_in(a10_wr[1263]),  .coef_in(coef[0]), .rdup_out(a11_wr[1262]), .rdlo_out(a11_wr[1263]));
			radix2 #(.width(width)) rd_st10_1264  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1264]), .rdlo_in(a10_wr[1265]),  .coef_in(coef[0]), .rdup_out(a11_wr[1264]), .rdlo_out(a11_wr[1265]));
			radix2 #(.width(width)) rd_st10_1266  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1266]), .rdlo_in(a10_wr[1267]),  .coef_in(coef[0]), .rdup_out(a11_wr[1266]), .rdlo_out(a11_wr[1267]));
			radix2 #(.width(width)) rd_st10_1268  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1268]), .rdlo_in(a10_wr[1269]),  .coef_in(coef[0]), .rdup_out(a11_wr[1268]), .rdlo_out(a11_wr[1269]));
			radix2 #(.width(width)) rd_st10_1270  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1270]), .rdlo_in(a10_wr[1271]),  .coef_in(coef[0]), .rdup_out(a11_wr[1270]), .rdlo_out(a11_wr[1271]));
			radix2 #(.width(width)) rd_st10_1272  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1272]), .rdlo_in(a10_wr[1273]),  .coef_in(coef[0]), .rdup_out(a11_wr[1272]), .rdlo_out(a11_wr[1273]));
			radix2 #(.width(width)) rd_st10_1274  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1274]), .rdlo_in(a10_wr[1275]),  .coef_in(coef[0]), .rdup_out(a11_wr[1274]), .rdlo_out(a11_wr[1275]));
			radix2 #(.width(width)) rd_st10_1276  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1276]), .rdlo_in(a10_wr[1277]),  .coef_in(coef[0]), .rdup_out(a11_wr[1276]), .rdlo_out(a11_wr[1277]));
			radix2 #(.width(width)) rd_st10_1278  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1278]), .rdlo_in(a10_wr[1279]),  .coef_in(coef[0]), .rdup_out(a11_wr[1278]), .rdlo_out(a11_wr[1279]));
			radix2 #(.width(width)) rd_st10_1280  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1280]), .rdlo_in(a10_wr[1281]),  .coef_in(coef[0]), .rdup_out(a11_wr[1280]), .rdlo_out(a11_wr[1281]));
			radix2 #(.width(width)) rd_st10_1282  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1282]), .rdlo_in(a10_wr[1283]),  .coef_in(coef[0]), .rdup_out(a11_wr[1282]), .rdlo_out(a11_wr[1283]));
			radix2 #(.width(width)) rd_st10_1284  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1284]), .rdlo_in(a10_wr[1285]),  .coef_in(coef[0]), .rdup_out(a11_wr[1284]), .rdlo_out(a11_wr[1285]));
			radix2 #(.width(width)) rd_st10_1286  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1286]), .rdlo_in(a10_wr[1287]),  .coef_in(coef[0]), .rdup_out(a11_wr[1286]), .rdlo_out(a11_wr[1287]));
			radix2 #(.width(width)) rd_st10_1288  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1288]), .rdlo_in(a10_wr[1289]),  .coef_in(coef[0]), .rdup_out(a11_wr[1288]), .rdlo_out(a11_wr[1289]));
			radix2 #(.width(width)) rd_st10_1290  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1290]), .rdlo_in(a10_wr[1291]),  .coef_in(coef[0]), .rdup_out(a11_wr[1290]), .rdlo_out(a11_wr[1291]));
			radix2 #(.width(width)) rd_st10_1292  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1292]), .rdlo_in(a10_wr[1293]),  .coef_in(coef[0]), .rdup_out(a11_wr[1292]), .rdlo_out(a11_wr[1293]));
			radix2 #(.width(width)) rd_st10_1294  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1294]), .rdlo_in(a10_wr[1295]),  .coef_in(coef[0]), .rdup_out(a11_wr[1294]), .rdlo_out(a11_wr[1295]));
			radix2 #(.width(width)) rd_st10_1296  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1296]), .rdlo_in(a10_wr[1297]),  .coef_in(coef[0]), .rdup_out(a11_wr[1296]), .rdlo_out(a11_wr[1297]));
			radix2 #(.width(width)) rd_st10_1298  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1298]), .rdlo_in(a10_wr[1299]),  .coef_in(coef[0]), .rdup_out(a11_wr[1298]), .rdlo_out(a11_wr[1299]));
			radix2 #(.width(width)) rd_st10_1300  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1300]), .rdlo_in(a10_wr[1301]),  .coef_in(coef[0]), .rdup_out(a11_wr[1300]), .rdlo_out(a11_wr[1301]));
			radix2 #(.width(width)) rd_st10_1302  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1302]), .rdlo_in(a10_wr[1303]),  .coef_in(coef[0]), .rdup_out(a11_wr[1302]), .rdlo_out(a11_wr[1303]));
			radix2 #(.width(width)) rd_st10_1304  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1304]), .rdlo_in(a10_wr[1305]),  .coef_in(coef[0]), .rdup_out(a11_wr[1304]), .rdlo_out(a11_wr[1305]));
			radix2 #(.width(width)) rd_st10_1306  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1306]), .rdlo_in(a10_wr[1307]),  .coef_in(coef[0]), .rdup_out(a11_wr[1306]), .rdlo_out(a11_wr[1307]));
			radix2 #(.width(width)) rd_st10_1308  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1308]), .rdlo_in(a10_wr[1309]),  .coef_in(coef[0]), .rdup_out(a11_wr[1308]), .rdlo_out(a11_wr[1309]));
			radix2 #(.width(width)) rd_st10_1310  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1310]), .rdlo_in(a10_wr[1311]),  .coef_in(coef[0]), .rdup_out(a11_wr[1310]), .rdlo_out(a11_wr[1311]));
			radix2 #(.width(width)) rd_st10_1312  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1312]), .rdlo_in(a10_wr[1313]),  .coef_in(coef[0]), .rdup_out(a11_wr[1312]), .rdlo_out(a11_wr[1313]));
			radix2 #(.width(width)) rd_st10_1314  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1314]), .rdlo_in(a10_wr[1315]),  .coef_in(coef[0]), .rdup_out(a11_wr[1314]), .rdlo_out(a11_wr[1315]));
			radix2 #(.width(width)) rd_st10_1316  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1316]), .rdlo_in(a10_wr[1317]),  .coef_in(coef[0]), .rdup_out(a11_wr[1316]), .rdlo_out(a11_wr[1317]));
			radix2 #(.width(width)) rd_st10_1318  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1318]), .rdlo_in(a10_wr[1319]),  .coef_in(coef[0]), .rdup_out(a11_wr[1318]), .rdlo_out(a11_wr[1319]));
			radix2 #(.width(width)) rd_st10_1320  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1320]), .rdlo_in(a10_wr[1321]),  .coef_in(coef[0]), .rdup_out(a11_wr[1320]), .rdlo_out(a11_wr[1321]));
			radix2 #(.width(width)) rd_st10_1322  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1322]), .rdlo_in(a10_wr[1323]),  .coef_in(coef[0]), .rdup_out(a11_wr[1322]), .rdlo_out(a11_wr[1323]));
			radix2 #(.width(width)) rd_st10_1324  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1324]), .rdlo_in(a10_wr[1325]),  .coef_in(coef[0]), .rdup_out(a11_wr[1324]), .rdlo_out(a11_wr[1325]));
			radix2 #(.width(width)) rd_st10_1326  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1326]), .rdlo_in(a10_wr[1327]),  .coef_in(coef[0]), .rdup_out(a11_wr[1326]), .rdlo_out(a11_wr[1327]));
			radix2 #(.width(width)) rd_st10_1328  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1328]), .rdlo_in(a10_wr[1329]),  .coef_in(coef[0]), .rdup_out(a11_wr[1328]), .rdlo_out(a11_wr[1329]));
			radix2 #(.width(width)) rd_st10_1330  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1330]), .rdlo_in(a10_wr[1331]),  .coef_in(coef[0]), .rdup_out(a11_wr[1330]), .rdlo_out(a11_wr[1331]));
			radix2 #(.width(width)) rd_st10_1332  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1332]), .rdlo_in(a10_wr[1333]),  .coef_in(coef[0]), .rdup_out(a11_wr[1332]), .rdlo_out(a11_wr[1333]));
			radix2 #(.width(width)) rd_st10_1334  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1334]), .rdlo_in(a10_wr[1335]),  .coef_in(coef[0]), .rdup_out(a11_wr[1334]), .rdlo_out(a11_wr[1335]));
			radix2 #(.width(width)) rd_st10_1336  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1336]), .rdlo_in(a10_wr[1337]),  .coef_in(coef[0]), .rdup_out(a11_wr[1336]), .rdlo_out(a11_wr[1337]));
			radix2 #(.width(width)) rd_st10_1338  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1338]), .rdlo_in(a10_wr[1339]),  .coef_in(coef[0]), .rdup_out(a11_wr[1338]), .rdlo_out(a11_wr[1339]));
			radix2 #(.width(width)) rd_st10_1340  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1340]), .rdlo_in(a10_wr[1341]),  .coef_in(coef[0]), .rdup_out(a11_wr[1340]), .rdlo_out(a11_wr[1341]));
			radix2 #(.width(width)) rd_st10_1342  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1342]), .rdlo_in(a10_wr[1343]),  .coef_in(coef[0]), .rdup_out(a11_wr[1342]), .rdlo_out(a11_wr[1343]));
			radix2 #(.width(width)) rd_st10_1344  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1344]), .rdlo_in(a10_wr[1345]),  .coef_in(coef[0]), .rdup_out(a11_wr[1344]), .rdlo_out(a11_wr[1345]));
			radix2 #(.width(width)) rd_st10_1346  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1346]), .rdlo_in(a10_wr[1347]),  .coef_in(coef[0]), .rdup_out(a11_wr[1346]), .rdlo_out(a11_wr[1347]));
			radix2 #(.width(width)) rd_st10_1348  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1348]), .rdlo_in(a10_wr[1349]),  .coef_in(coef[0]), .rdup_out(a11_wr[1348]), .rdlo_out(a11_wr[1349]));
			radix2 #(.width(width)) rd_st10_1350  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1350]), .rdlo_in(a10_wr[1351]),  .coef_in(coef[0]), .rdup_out(a11_wr[1350]), .rdlo_out(a11_wr[1351]));
			radix2 #(.width(width)) rd_st10_1352  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1352]), .rdlo_in(a10_wr[1353]),  .coef_in(coef[0]), .rdup_out(a11_wr[1352]), .rdlo_out(a11_wr[1353]));
			radix2 #(.width(width)) rd_st10_1354  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1354]), .rdlo_in(a10_wr[1355]),  .coef_in(coef[0]), .rdup_out(a11_wr[1354]), .rdlo_out(a11_wr[1355]));
			radix2 #(.width(width)) rd_st10_1356  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1356]), .rdlo_in(a10_wr[1357]),  .coef_in(coef[0]), .rdup_out(a11_wr[1356]), .rdlo_out(a11_wr[1357]));
			radix2 #(.width(width)) rd_st10_1358  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1358]), .rdlo_in(a10_wr[1359]),  .coef_in(coef[0]), .rdup_out(a11_wr[1358]), .rdlo_out(a11_wr[1359]));
			radix2 #(.width(width)) rd_st10_1360  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1360]), .rdlo_in(a10_wr[1361]),  .coef_in(coef[0]), .rdup_out(a11_wr[1360]), .rdlo_out(a11_wr[1361]));
			radix2 #(.width(width)) rd_st10_1362  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1362]), .rdlo_in(a10_wr[1363]),  .coef_in(coef[0]), .rdup_out(a11_wr[1362]), .rdlo_out(a11_wr[1363]));
			radix2 #(.width(width)) rd_st10_1364  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1364]), .rdlo_in(a10_wr[1365]),  .coef_in(coef[0]), .rdup_out(a11_wr[1364]), .rdlo_out(a11_wr[1365]));
			radix2 #(.width(width)) rd_st10_1366  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1366]), .rdlo_in(a10_wr[1367]),  .coef_in(coef[0]), .rdup_out(a11_wr[1366]), .rdlo_out(a11_wr[1367]));
			radix2 #(.width(width)) rd_st10_1368  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1368]), .rdlo_in(a10_wr[1369]),  .coef_in(coef[0]), .rdup_out(a11_wr[1368]), .rdlo_out(a11_wr[1369]));
			radix2 #(.width(width)) rd_st10_1370  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1370]), .rdlo_in(a10_wr[1371]),  .coef_in(coef[0]), .rdup_out(a11_wr[1370]), .rdlo_out(a11_wr[1371]));
			radix2 #(.width(width)) rd_st10_1372  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1372]), .rdlo_in(a10_wr[1373]),  .coef_in(coef[0]), .rdup_out(a11_wr[1372]), .rdlo_out(a11_wr[1373]));
			radix2 #(.width(width)) rd_st10_1374  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1374]), .rdlo_in(a10_wr[1375]),  .coef_in(coef[0]), .rdup_out(a11_wr[1374]), .rdlo_out(a11_wr[1375]));
			radix2 #(.width(width)) rd_st10_1376  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1376]), .rdlo_in(a10_wr[1377]),  .coef_in(coef[0]), .rdup_out(a11_wr[1376]), .rdlo_out(a11_wr[1377]));
			radix2 #(.width(width)) rd_st10_1378  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1378]), .rdlo_in(a10_wr[1379]),  .coef_in(coef[0]), .rdup_out(a11_wr[1378]), .rdlo_out(a11_wr[1379]));
			radix2 #(.width(width)) rd_st10_1380  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1380]), .rdlo_in(a10_wr[1381]),  .coef_in(coef[0]), .rdup_out(a11_wr[1380]), .rdlo_out(a11_wr[1381]));
			radix2 #(.width(width)) rd_st10_1382  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1382]), .rdlo_in(a10_wr[1383]),  .coef_in(coef[0]), .rdup_out(a11_wr[1382]), .rdlo_out(a11_wr[1383]));
			radix2 #(.width(width)) rd_st10_1384  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1384]), .rdlo_in(a10_wr[1385]),  .coef_in(coef[0]), .rdup_out(a11_wr[1384]), .rdlo_out(a11_wr[1385]));
			radix2 #(.width(width)) rd_st10_1386  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1386]), .rdlo_in(a10_wr[1387]),  .coef_in(coef[0]), .rdup_out(a11_wr[1386]), .rdlo_out(a11_wr[1387]));
			radix2 #(.width(width)) rd_st10_1388  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1388]), .rdlo_in(a10_wr[1389]),  .coef_in(coef[0]), .rdup_out(a11_wr[1388]), .rdlo_out(a11_wr[1389]));
			radix2 #(.width(width)) rd_st10_1390  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1390]), .rdlo_in(a10_wr[1391]),  .coef_in(coef[0]), .rdup_out(a11_wr[1390]), .rdlo_out(a11_wr[1391]));
			radix2 #(.width(width)) rd_st10_1392  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1392]), .rdlo_in(a10_wr[1393]),  .coef_in(coef[0]), .rdup_out(a11_wr[1392]), .rdlo_out(a11_wr[1393]));
			radix2 #(.width(width)) rd_st10_1394  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1394]), .rdlo_in(a10_wr[1395]),  .coef_in(coef[0]), .rdup_out(a11_wr[1394]), .rdlo_out(a11_wr[1395]));
			radix2 #(.width(width)) rd_st10_1396  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1396]), .rdlo_in(a10_wr[1397]),  .coef_in(coef[0]), .rdup_out(a11_wr[1396]), .rdlo_out(a11_wr[1397]));
			radix2 #(.width(width)) rd_st10_1398  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1398]), .rdlo_in(a10_wr[1399]),  .coef_in(coef[0]), .rdup_out(a11_wr[1398]), .rdlo_out(a11_wr[1399]));
			radix2 #(.width(width)) rd_st10_1400  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1400]), .rdlo_in(a10_wr[1401]),  .coef_in(coef[0]), .rdup_out(a11_wr[1400]), .rdlo_out(a11_wr[1401]));
			radix2 #(.width(width)) rd_st10_1402  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1402]), .rdlo_in(a10_wr[1403]),  .coef_in(coef[0]), .rdup_out(a11_wr[1402]), .rdlo_out(a11_wr[1403]));
			radix2 #(.width(width)) rd_st10_1404  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1404]), .rdlo_in(a10_wr[1405]),  .coef_in(coef[0]), .rdup_out(a11_wr[1404]), .rdlo_out(a11_wr[1405]));
			radix2 #(.width(width)) rd_st10_1406  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1406]), .rdlo_in(a10_wr[1407]),  .coef_in(coef[0]), .rdup_out(a11_wr[1406]), .rdlo_out(a11_wr[1407]));
			radix2 #(.width(width)) rd_st10_1408  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1408]), .rdlo_in(a10_wr[1409]),  .coef_in(coef[0]), .rdup_out(a11_wr[1408]), .rdlo_out(a11_wr[1409]));
			radix2 #(.width(width)) rd_st10_1410  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1410]), .rdlo_in(a10_wr[1411]),  .coef_in(coef[0]), .rdup_out(a11_wr[1410]), .rdlo_out(a11_wr[1411]));
			radix2 #(.width(width)) rd_st10_1412  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1412]), .rdlo_in(a10_wr[1413]),  .coef_in(coef[0]), .rdup_out(a11_wr[1412]), .rdlo_out(a11_wr[1413]));
			radix2 #(.width(width)) rd_st10_1414  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1414]), .rdlo_in(a10_wr[1415]),  .coef_in(coef[0]), .rdup_out(a11_wr[1414]), .rdlo_out(a11_wr[1415]));
			radix2 #(.width(width)) rd_st10_1416  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1416]), .rdlo_in(a10_wr[1417]),  .coef_in(coef[0]), .rdup_out(a11_wr[1416]), .rdlo_out(a11_wr[1417]));
			radix2 #(.width(width)) rd_st10_1418  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1418]), .rdlo_in(a10_wr[1419]),  .coef_in(coef[0]), .rdup_out(a11_wr[1418]), .rdlo_out(a11_wr[1419]));
			radix2 #(.width(width)) rd_st10_1420  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1420]), .rdlo_in(a10_wr[1421]),  .coef_in(coef[0]), .rdup_out(a11_wr[1420]), .rdlo_out(a11_wr[1421]));
			radix2 #(.width(width)) rd_st10_1422  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1422]), .rdlo_in(a10_wr[1423]),  .coef_in(coef[0]), .rdup_out(a11_wr[1422]), .rdlo_out(a11_wr[1423]));
			radix2 #(.width(width)) rd_st10_1424  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1424]), .rdlo_in(a10_wr[1425]),  .coef_in(coef[0]), .rdup_out(a11_wr[1424]), .rdlo_out(a11_wr[1425]));
			radix2 #(.width(width)) rd_st10_1426  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1426]), .rdlo_in(a10_wr[1427]),  .coef_in(coef[0]), .rdup_out(a11_wr[1426]), .rdlo_out(a11_wr[1427]));
			radix2 #(.width(width)) rd_st10_1428  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1428]), .rdlo_in(a10_wr[1429]),  .coef_in(coef[0]), .rdup_out(a11_wr[1428]), .rdlo_out(a11_wr[1429]));
			radix2 #(.width(width)) rd_st10_1430  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1430]), .rdlo_in(a10_wr[1431]),  .coef_in(coef[0]), .rdup_out(a11_wr[1430]), .rdlo_out(a11_wr[1431]));
			radix2 #(.width(width)) rd_st10_1432  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1432]), .rdlo_in(a10_wr[1433]),  .coef_in(coef[0]), .rdup_out(a11_wr[1432]), .rdlo_out(a11_wr[1433]));
			radix2 #(.width(width)) rd_st10_1434  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1434]), .rdlo_in(a10_wr[1435]),  .coef_in(coef[0]), .rdup_out(a11_wr[1434]), .rdlo_out(a11_wr[1435]));
			radix2 #(.width(width)) rd_st10_1436  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1436]), .rdlo_in(a10_wr[1437]),  .coef_in(coef[0]), .rdup_out(a11_wr[1436]), .rdlo_out(a11_wr[1437]));
			radix2 #(.width(width)) rd_st10_1438  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1438]), .rdlo_in(a10_wr[1439]),  .coef_in(coef[0]), .rdup_out(a11_wr[1438]), .rdlo_out(a11_wr[1439]));
			radix2 #(.width(width)) rd_st10_1440  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1440]), .rdlo_in(a10_wr[1441]),  .coef_in(coef[0]), .rdup_out(a11_wr[1440]), .rdlo_out(a11_wr[1441]));
			radix2 #(.width(width)) rd_st10_1442  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1442]), .rdlo_in(a10_wr[1443]),  .coef_in(coef[0]), .rdup_out(a11_wr[1442]), .rdlo_out(a11_wr[1443]));
			radix2 #(.width(width)) rd_st10_1444  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1444]), .rdlo_in(a10_wr[1445]),  .coef_in(coef[0]), .rdup_out(a11_wr[1444]), .rdlo_out(a11_wr[1445]));
			radix2 #(.width(width)) rd_st10_1446  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1446]), .rdlo_in(a10_wr[1447]),  .coef_in(coef[0]), .rdup_out(a11_wr[1446]), .rdlo_out(a11_wr[1447]));
			radix2 #(.width(width)) rd_st10_1448  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1448]), .rdlo_in(a10_wr[1449]),  .coef_in(coef[0]), .rdup_out(a11_wr[1448]), .rdlo_out(a11_wr[1449]));
			radix2 #(.width(width)) rd_st10_1450  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1450]), .rdlo_in(a10_wr[1451]),  .coef_in(coef[0]), .rdup_out(a11_wr[1450]), .rdlo_out(a11_wr[1451]));
			radix2 #(.width(width)) rd_st10_1452  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1452]), .rdlo_in(a10_wr[1453]),  .coef_in(coef[0]), .rdup_out(a11_wr[1452]), .rdlo_out(a11_wr[1453]));
			radix2 #(.width(width)) rd_st10_1454  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1454]), .rdlo_in(a10_wr[1455]),  .coef_in(coef[0]), .rdup_out(a11_wr[1454]), .rdlo_out(a11_wr[1455]));
			radix2 #(.width(width)) rd_st10_1456  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1456]), .rdlo_in(a10_wr[1457]),  .coef_in(coef[0]), .rdup_out(a11_wr[1456]), .rdlo_out(a11_wr[1457]));
			radix2 #(.width(width)) rd_st10_1458  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1458]), .rdlo_in(a10_wr[1459]),  .coef_in(coef[0]), .rdup_out(a11_wr[1458]), .rdlo_out(a11_wr[1459]));
			radix2 #(.width(width)) rd_st10_1460  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1460]), .rdlo_in(a10_wr[1461]),  .coef_in(coef[0]), .rdup_out(a11_wr[1460]), .rdlo_out(a11_wr[1461]));
			radix2 #(.width(width)) rd_st10_1462  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1462]), .rdlo_in(a10_wr[1463]),  .coef_in(coef[0]), .rdup_out(a11_wr[1462]), .rdlo_out(a11_wr[1463]));
			radix2 #(.width(width)) rd_st10_1464  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1464]), .rdlo_in(a10_wr[1465]),  .coef_in(coef[0]), .rdup_out(a11_wr[1464]), .rdlo_out(a11_wr[1465]));
			radix2 #(.width(width)) rd_st10_1466  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1466]), .rdlo_in(a10_wr[1467]),  .coef_in(coef[0]), .rdup_out(a11_wr[1466]), .rdlo_out(a11_wr[1467]));
			radix2 #(.width(width)) rd_st10_1468  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1468]), .rdlo_in(a10_wr[1469]),  .coef_in(coef[0]), .rdup_out(a11_wr[1468]), .rdlo_out(a11_wr[1469]));
			radix2 #(.width(width)) rd_st10_1470  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1470]), .rdlo_in(a10_wr[1471]),  .coef_in(coef[0]), .rdup_out(a11_wr[1470]), .rdlo_out(a11_wr[1471]));
			radix2 #(.width(width)) rd_st10_1472  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1472]), .rdlo_in(a10_wr[1473]),  .coef_in(coef[0]), .rdup_out(a11_wr[1472]), .rdlo_out(a11_wr[1473]));
			radix2 #(.width(width)) rd_st10_1474  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1474]), .rdlo_in(a10_wr[1475]),  .coef_in(coef[0]), .rdup_out(a11_wr[1474]), .rdlo_out(a11_wr[1475]));
			radix2 #(.width(width)) rd_st10_1476  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1476]), .rdlo_in(a10_wr[1477]),  .coef_in(coef[0]), .rdup_out(a11_wr[1476]), .rdlo_out(a11_wr[1477]));
			radix2 #(.width(width)) rd_st10_1478  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1478]), .rdlo_in(a10_wr[1479]),  .coef_in(coef[0]), .rdup_out(a11_wr[1478]), .rdlo_out(a11_wr[1479]));
			radix2 #(.width(width)) rd_st10_1480  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1480]), .rdlo_in(a10_wr[1481]),  .coef_in(coef[0]), .rdup_out(a11_wr[1480]), .rdlo_out(a11_wr[1481]));
			radix2 #(.width(width)) rd_st10_1482  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1482]), .rdlo_in(a10_wr[1483]),  .coef_in(coef[0]), .rdup_out(a11_wr[1482]), .rdlo_out(a11_wr[1483]));
			radix2 #(.width(width)) rd_st10_1484  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1484]), .rdlo_in(a10_wr[1485]),  .coef_in(coef[0]), .rdup_out(a11_wr[1484]), .rdlo_out(a11_wr[1485]));
			radix2 #(.width(width)) rd_st10_1486  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1486]), .rdlo_in(a10_wr[1487]),  .coef_in(coef[0]), .rdup_out(a11_wr[1486]), .rdlo_out(a11_wr[1487]));
			radix2 #(.width(width)) rd_st10_1488  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1488]), .rdlo_in(a10_wr[1489]),  .coef_in(coef[0]), .rdup_out(a11_wr[1488]), .rdlo_out(a11_wr[1489]));
			radix2 #(.width(width)) rd_st10_1490  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1490]), .rdlo_in(a10_wr[1491]),  .coef_in(coef[0]), .rdup_out(a11_wr[1490]), .rdlo_out(a11_wr[1491]));
			radix2 #(.width(width)) rd_st10_1492  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1492]), .rdlo_in(a10_wr[1493]),  .coef_in(coef[0]), .rdup_out(a11_wr[1492]), .rdlo_out(a11_wr[1493]));
			radix2 #(.width(width)) rd_st10_1494  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1494]), .rdlo_in(a10_wr[1495]),  .coef_in(coef[0]), .rdup_out(a11_wr[1494]), .rdlo_out(a11_wr[1495]));
			radix2 #(.width(width)) rd_st10_1496  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1496]), .rdlo_in(a10_wr[1497]),  .coef_in(coef[0]), .rdup_out(a11_wr[1496]), .rdlo_out(a11_wr[1497]));
			radix2 #(.width(width)) rd_st10_1498  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1498]), .rdlo_in(a10_wr[1499]),  .coef_in(coef[0]), .rdup_out(a11_wr[1498]), .rdlo_out(a11_wr[1499]));
			radix2 #(.width(width)) rd_st10_1500  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1500]), .rdlo_in(a10_wr[1501]),  .coef_in(coef[0]), .rdup_out(a11_wr[1500]), .rdlo_out(a11_wr[1501]));
			radix2 #(.width(width)) rd_st10_1502  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1502]), .rdlo_in(a10_wr[1503]),  .coef_in(coef[0]), .rdup_out(a11_wr[1502]), .rdlo_out(a11_wr[1503]));
			radix2 #(.width(width)) rd_st10_1504  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1504]), .rdlo_in(a10_wr[1505]),  .coef_in(coef[0]), .rdup_out(a11_wr[1504]), .rdlo_out(a11_wr[1505]));
			radix2 #(.width(width)) rd_st10_1506  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1506]), .rdlo_in(a10_wr[1507]),  .coef_in(coef[0]), .rdup_out(a11_wr[1506]), .rdlo_out(a11_wr[1507]));
			radix2 #(.width(width)) rd_st10_1508  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1508]), .rdlo_in(a10_wr[1509]),  .coef_in(coef[0]), .rdup_out(a11_wr[1508]), .rdlo_out(a11_wr[1509]));
			radix2 #(.width(width)) rd_st10_1510  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1510]), .rdlo_in(a10_wr[1511]),  .coef_in(coef[0]), .rdup_out(a11_wr[1510]), .rdlo_out(a11_wr[1511]));
			radix2 #(.width(width)) rd_st10_1512  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1512]), .rdlo_in(a10_wr[1513]),  .coef_in(coef[0]), .rdup_out(a11_wr[1512]), .rdlo_out(a11_wr[1513]));
			radix2 #(.width(width)) rd_st10_1514  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1514]), .rdlo_in(a10_wr[1515]),  .coef_in(coef[0]), .rdup_out(a11_wr[1514]), .rdlo_out(a11_wr[1515]));
			radix2 #(.width(width)) rd_st10_1516  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1516]), .rdlo_in(a10_wr[1517]),  .coef_in(coef[0]), .rdup_out(a11_wr[1516]), .rdlo_out(a11_wr[1517]));
			radix2 #(.width(width)) rd_st10_1518  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1518]), .rdlo_in(a10_wr[1519]),  .coef_in(coef[0]), .rdup_out(a11_wr[1518]), .rdlo_out(a11_wr[1519]));
			radix2 #(.width(width)) rd_st10_1520  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1520]), .rdlo_in(a10_wr[1521]),  .coef_in(coef[0]), .rdup_out(a11_wr[1520]), .rdlo_out(a11_wr[1521]));
			radix2 #(.width(width)) rd_st10_1522  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1522]), .rdlo_in(a10_wr[1523]),  .coef_in(coef[0]), .rdup_out(a11_wr[1522]), .rdlo_out(a11_wr[1523]));
			radix2 #(.width(width)) rd_st10_1524  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1524]), .rdlo_in(a10_wr[1525]),  .coef_in(coef[0]), .rdup_out(a11_wr[1524]), .rdlo_out(a11_wr[1525]));
			radix2 #(.width(width)) rd_st10_1526  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1526]), .rdlo_in(a10_wr[1527]),  .coef_in(coef[0]), .rdup_out(a11_wr[1526]), .rdlo_out(a11_wr[1527]));
			radix2 #(.width(width)) rd_st10_1528  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1528]), .rdlo_in(a10_wr[1529]),  .coef_in(coef[0]), .rdup_out(a11_wr[1528]), .rdlo_out(a11_wr[1529]));
			radix2 #(.width(width)) rd_st10_1530  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1530]), .rdlo_in(a10_wr[1531]),  .coef_in(coef[0]), .rdup_out(a11_wr[1530]), .rdlo_out(a11_wr[1531]));
			radix2 #(.width(width)) rd_st10_1532  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1532]), .rdlo_in(a10_wr[1533]),  .coef_in(coef[0]), .rdup_out(a11_wr[1532]), .rdlo_out(a11_wr[1533]));
			radix2 #(.width(width)) rd_st10_1534  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1534]), .rdlo_in(a10_wr[1535]),  .coef_in(coef[0]), .rdup_out(a11_wr[1534]), .rdlo_out(a11_wr[1535]));
			radix2 #(.width(width)) rd_st10_1536  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1536]), .rdlo_in(a10_wr[1537]),  .coef_in(coef[0]), .rdup_out(a11_wr[1536]), .rdlo_out(a11_wr[1537]));
			radix2 #(.width(width)) rd_st10_1538  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1538]), .rdlo_in(a10_wr[1539]),  .coef_in(coef[0]), .rdup_out(a11_wr[1538]), .rdlo_out(a11_wr[1539]));
			radix2 #(.width(width)) rd_st10_1540  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1540]), .rdlo_in(a10_wr[1541]),  .coef_in(coef[0]), .rdup_out(a11_wr[1540]), .rdlo_out(a11_wr[1541]));
			radix2 #(.width(width)) rd_st10_1542  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1542]), .rdlo_in(a10_wr[1543]),  .coef_in(coef[0]), .rdup_out(a11_wr[1542]), .rdlo_out(a11_wr[1543]));
			radix2 #(.width(width)) rd_st10_1544  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1544]), .rdlo_in(a10_wr[1545]),  .coef_in(coef[0]), .rdup_out(a11_wr[1544]), .rdlo_out(a11_wr[1545]));
			radix2 #(.width(width)) rd_st10_1546  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1546]), .rdlo_in(a10_wr[1547]),  .coef_in(coef[0]), .rdup_out(a11_wr[1546]), .rdlo_out(a11_wr[1547]));
			radix2 #(.width(width)) rd_st10_1548  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1548]), .rdlo_in(a10_wr[1549]),  .coef_in(coef[0]), .rdup_out(a11_wr[1548]), .rdlo_out(a11_wr[1549]));
			radix2 #(.width(width)) rd_st10_1550  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1550]), .rdlo_in(a10_wr[1551]),  .coef_in(coef[0]), .rdup_out(a11_wr[1550]), .rdlo_out(a11_wr[1551]));
			radix2 #(.width(width)) rd_st10_1552  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1552]), .rdlo_in(a10_wr[1553]),  .coef_in(coef[0]), .rdup_out(a11_wr[1552]), .rdlo_out(a11_wr[1553]));
			radix2 #(.width(width)) rd_st10_1554  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1554]), .rdlo_in(a10_wr[1555]),  .coef_in(coef[0]), .rdup_out(a11_wr[1554]), .rdlo_out(a11_wr[1555]));
			radix2 #(.width(width)) rd_st10_1556  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1556]), .rdlo_in(a10_wr[1557]),  .coef_in(coef[0]), .rdup_out(a11_wr[1556]), .rdlo_out(a11_wr[1557]));
			radix2 #(.width(width)) rd_st10_1558  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1558]), .rdlo_in(a10_wr[1559]),  .coef_in(coef[0]), .rdup_out(a11_wr[1558]), .rdlo_out(a11_wr[1559]));
			radix2 #(.width(width)) rd_st10_1560  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1560]), .rdlo_in(a10_wr[1561]),  .coef_in(coef[0]), .rdup_out(a11_wr[1560]), .rdlo_out(a11_wr[1561]));
			radix2 #(.width(width)) rd_st10_1562  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1562]), .rdlo_in(a10_wr[1563]),  .coef_in(coef[0]), .rdup_out(a11_wr[1562]), .rdlo_out(a11_wr[1563]));
			radix2 #(.width(width)) rd_st10_1564  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1564]), .rdlo_in(a10_wr[1565]),  .coef_in(coef[0]), .rdup_out(a11_wr[1564]), .rdlo_out(a11_wr[1565]));
			radix2 #(.width(width)) rd_st10_1566  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1566]), .rdlo_in(a10_wr[1567]),  .coef_in(coef[0]), .rdup_out(a11_wr[1566]), .rdlo_out(a11_wr[1567]));
			radix2 #(.width(width)) rd_st10_1568  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1568]), .rdlo_in(a10_wr[1569]),  .coef_in(coef[0]), .rdup_out(a11_wr[1568]), .rdlo_out(a11_wr[1569]));
			radix2 #(.width(width)) rd_st10_1570  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1570]), .rdlo_in(a10_wr[1571]),  .coef_in(coef[0]), .rdup_out(a11_wr[1570]), .rdlo_out(a11_wr[1571]));
			radix2 #(.width(width)) rd_st10_1572  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1572]), .rdlo_in(a10_wr[1573]),  .coef_in(coef[0]), .rdup_out(a11_wr[1572]), .rdlo_out(a11_wr[1573]));
			radix2 #(.width(width)) rd_st10_1574  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1574]), .rdlo_in(a10_wr[1575]),  .coef_in(coef[0]), .rdup_out(a11_wr[1574]), .rdlo_out(a11_wr[1575]));
			radix2 #(.width(width)) rd_st10_1576  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1576]), .rdlo_in(a10_wr[1577]),  .coef_in(coef[0]), .rdup_out(a11_wr[1576]), .rdlo_out(a11_wr[1577]));
			radix2 #(.width(width)) rd_st10_1578  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1578]), .rdlo_in(a10_wr[1579]),  .coef_in(coef[0]), .rdup_out(a11_wr[1578]), .rdlo_out(a11_wr[1579]));
			radix2 #(.width(width)) rd_st10_1580  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1580]), .rdlo_in(a10_wr[1581]),  .coef_in(coef[0]), .rdup_out(a11_wr[1580]), .rdlo_out(a11_wr[1581]));
			radix2 #(.width(width)) rd_st10_1582  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1582]), .rdlo_in(a10_wr[1583]),  .coef_in(coef[0]), .rdup_out(a11_wr[1582]), .rdlo_out(a11_wr[1583]));
			radix2 #(.width(width)) rd_st10_1584  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1584]), .rdlo_in(a10_wr[1585]),  .coef_in(coef[0]), .rdup_out(a11_wr[1584]), .rdlo_out(a11_wr[1585]));
			radix2 #(.width(width)) rd_st10_1586  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1586]), .rdlo_in(a10_wr[1587]),  .coef_in(coef[0]), .rdup_out(a11_wr[1586]), .rdlo_out(a11_wr[1587]));
			radix2 #(.width(width)) rd_st10_1588  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1588]), .rdlo_in(a10_wr[1589]),  .coef_in(coef[0]), .rdup_out(a11_wr[1588]), .rdlo_out(a11_wr[1589]));
			radix2 #(.width(width)) rd_st10_1590  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1590]), .rdlo_in(a10_wr[1591]),  .coef_in(coef[0]), .rdup_out(a11_wr[1590]), .rdlo_out(a11_wr[1591]));
			radix2 #(.width(width)) rd_st10_1592  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1592]), .rdlo_in(a10_wr[1593]),  .coef_in(coef[0]), .rdup_out(a11_wr[1592]), .rdlo_out(a11_wr[1593]));
			radix2 #(.width(width)) rd_st10_1594  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1594]), .rdlo_in(a10_wr[1595]),  .coef_in(coef[0]), .rdup_out(a11_wr[1594]), .rdlo_out(a11_wr[1595]));
			radix2 #(.width(width)) rd_st10_1596  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1596]), .rdlo_in(a10_wr[1597]),  .coef_in(coef[0]), .rdup_out(a11_wr[1596]), .rdlo_out(a11_wr[1597]));
			radix2 #(.width(width)) rd_st10_1598  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1598]), .rdlo_in(a10_wr[1599]),  .coef_in(coef[0]), .rdup_out(a11_wr[1598]), .rdlo_out(a11_wr[1599]));
			radix2 #(.width(width)) rd_st10_1600  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1600]), .rdlo_in(a10_wr[1601]),  .coef_in(coef[0]), .rdup_out(a11_wr[1600]), .rdlo_out(a11_wr[1601]));
			radix2 #(.width(width)) rd_st10_1602  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1602]), .rdlo_in(a10_wr[1603]),  .coef_in(coef[0]), .rdup_out(a11_wr[1602]), .rdlo_out(a11_wr[1603]));
			radix2 #(.width(width)) rd_st10_1604  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1604]), .rdlo_in(a10_wr[1605]),  .coef_in(coef[0]), .rdup_out(a11_wr[1604]), .rdlo_out(a11_wr[1605]));
			radix2 #(.width(width)) rd_st10_1606  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1606]), .rdlo_in(a10_wr[1607]),  .coef_in(coef[0]), .rdup_out(a11_wr[1606]), .rdlo_out(a11_wr[1607]));
			radix2 #(.width(width)) rd_st10_1608  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1608]), .rdlo_in(a10_wr[1609]),  .coef_in(coef[0]), .rdup_out(a11_wr[1608]), .rdlo_out(a11_wr[1609]));
			radix2 #(.width(width)) rd_st10_1610  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1610]), .rdlo_in(a10_wr[1611]),  .coef_in(coef[0]), .rdup_out(a11_wr[1610]), .rdlo_out(a11_wr[1611]));
			radix2 #(.width(width)) rd_st10_1612  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1612]), .rdlo_in(a10_wr[1613]),  .coef_in(coef[0]), .rdup_out(a11_wr[1612]), .rdlo_out(a11_wr[1613]));
			radix2 #(.width(width)) rd_st10_1614  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1614]), .rdlo_in(a10_wr[1615]),  .coef_in(coef[0]), .rdup_out(a11_wr[1614]), .rdlo_out(a11_wr[1615]));
			radix2 #(.width(width)) rd_st10_1616  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1616]), .rdlo_in(a10_wr[1617]),  .coef_in(coef[0]), .rdup_out(a11_wr[1616]), .rdlo_out(a11_wr[1617]));
			radix2 #(.width(width)) rd_st10_1618  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1618]), .rdlo_in(a10_wr[1619]),  .coef_in(coef[0]), .rdup_out(a11_wr[1618]), .rdlo_out(a11_wr[1619]));
			radix2 #(.width(width)) rd_st10_1620  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1620]), .rdlo_in(a10_wr[1621]),  .coef_in(coef[0]), .rdup_out(a11_wr[1620]), .rdlo_out(a11_wr[1621]));
			radix2 #(.width(width)) rd_st10_1622  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1622]), .rdlo_in(a10_wr[1623]),  .coef_in(coef[0]), .rdup_out(a11_wr[1622]), .rdlo_out(a11_wr[1623]));
			radix2 #(.width(width)) rd_st10_1624  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1624]), .rdlo_in(a10_wr[1625]),  .coef_in(coef[0]), .rdup_out(a11_wr[1624]), .rdlo_out(a11_wr[1625]));
			radix2 #(.width(width)) rd_st10_1626  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1626]), .rdlo_in(a10_wr[1627]),  .coef_in(coef[0]), .rdup_out(a11_wr[1626]), .rdlo_out(a11_wr[1627]));
			radix2 #(.width(width)) rd_st10_1628  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1628]), .rdlo_in(a10_wr[1629]),  .coef_in(coef[0]), .rdup_out(a11_wr[1628]), .rdlo_out(a11_wr[1629]));
			radix2 #(.width(width)) rd_st10_1630  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1630]), .rdlo_in(a10_wr[1631]),  .coef_in(coef[0]), .rdup_out(a11_wr[1630]), .rdlo_out(a11_wr[1631]));
			radix2 #(.width(width)) rd_st10_1632  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1632]), .rdlo_in(a10_wr[1633]),  .coef_in(coef[0]), .rdup_out(a11_wr[1632]), .rdlo_out(a11_wr[1633]));
			radix2 #(.width(width)) rd_st10_1634  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1634]), .rdlo_in(a10_wr[1635]),  .coef_in(coef[0]), .rdup_out(a11_wr[1634]), .rdlo_out(a11_wr[1635]));
			radix2 #(.width(width)) rd_st10_1636  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1636]), .rdlo_in(a10_wr[1637]),  .coef_in(coef[0]), .rdup_out(a11_wr[1636]), .rdlo_out(a11_wr[1637]));
			radix2 #(.width(width)) rd_st10_1638  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1638]), .rdlo_in(a10_wr[1639]),  .coef_in(coef[0]), .rdup_out(a11_wr[1638]), .rdlo_out(a11_wr[1639]));
			radix2 #(.width(width)) rd_st10_1640  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1640]), .rdlo_in(a10_wr[1641]),  .coef_in(coef[0]), .rdup_out(a11_wr[1640]), .rdlo_out(a11_wr[1641]));
			radix2 #(.width(width)) rd_st10_1642  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1642]), .rdlo_in(a10_wr[1643]),  .coef_in(coef[0]), .rdup_out(a11_wr[1642]), .rdlo_out(a11_wr[1643]));
			radix2 #(.width(width)) rd_st10_1644  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1644]), .rdlo_in(a10_wr[1645]),  .coef_in(coef[0]), .rdup_out(a11_wr[1644]), .rdlo_out(a11_wr[1645]));
			radix2 #(.width(width)) rd_st10_1646  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1646]), .rdlo_in(a10_wr[1647]),  .coef_in(coef[0]), .rdup_out(a11_wr[1646]), .rdlo_out(a11_wr[1647]));
			radix2 #(.width(width)) rd_st10_1648  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1648]), .rdlo_in(a10_wr[1649]),  .coef_in(coef[0]), .rdup_out(a11_wr[1648]), .rdlo_out(a11_wr[1649]));
			radix2 #(.width(width)) rd_st10_1650  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1650]), .rdlo_in(a10_wr[1651]),  .coef_in(coef[0]), .rdup_out(a11_wr[1650]), .rdlo_out(a11_wr[1651]));
			radix2 #(.width(width)) rd_st10_1652  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1652]), .rdlo_in(a10_wr[1653]),  .coef_in(coef[0]), .rdup_out(a11_wr[1652]), .rdlo_out(a11_wr[1653]));
			radix2 #(.width(width)) rd_st10_1654  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1654]), .rdlo_in(a10_wr[1655]),  .coef_in(coef[0]), .rdup_out(a11_wr[1654]), .rdlo_out(a11_wr[1655]));
			radix2 #(.width(width)) rd_st10_1656  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1656]), .rdlo_in(a10_wr[1657]),  .coef_in(coef[0]), .rdup_out(a11_wr[1656]), .rdlo_out(a11_wr[1657]));
			radix2 #(.width(width)) rd_st10_1658  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1658]), .rdlo_in(a10_wr[1659]),  .coef_in(coef[0]), .rdup_out(a11_wr[1658]), .rdlo_out(a11_wr[1659]));
			radix2 #(.width(width)) rd_st10_1660  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1660]), .rdlo_in(a10_wr[1661]),  .coef_in(coef[0]), .rdup_out(a11_wr[1660]), .rdlo_out(a11_wr[1661]));
			radix2 #(.width(width)) rd_st10_1662  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1662]), .rdlo_in(a10_wr[1663]),  .coef_in(coef[0]), .rdup_out(a11_wr[1662]), .rdlo_out(a11_wr[1663]));
			radix2 #(.width(width)) rd_st10_1664  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1664]), .rdlo_in(a10_wr[1665]),  .coef_in(coef[0]), .rdup_out(a11_wr[1664]), .rdlo_out(a11_wr[1665]));
			radix2 #(.width(width)) rd_st10_1666  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1666]), .rdlo_in(a10_wr[1667]),  .coef_in(coef[0]), .rdup_out(a11_wr[1666]), .rdlo_out(a11_wr[1667]));
			radix2 #(.width(width)) rd_st10_1668  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1668]), .rdlo_in(a10_wr[1669]),  .coef_in(coef[0]), .rdup_out(a11_wr[1668]), .rdlo_out(a11_wr[1669]));
			radix2 #(.width(width)) rd_st10_1670  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1670]), .rdlo_in(a10_wr[1671]),  .coef_in(coef[0]), .rdup_out(a11_wr[1670]), .rdlo_out(a11_wr[1671]));
			radix2 #(.width(width)) rd_st10_1672  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1672]), .rdlo_in(a10_wr[1673]),  .coef_in(coef[0]), .rdup_out(a11_wr[1672]), .rdlo_out(a11_wr[1673]));
			radix2 #(.width(width)) rd_st10_1674  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1674]), .rdlo_in(a10_wr[1675]),  .coef_in(coef[0]), .rdup_out(a11_wr[1674]), .rdlo_out(a11_wr[1675]));
			radix2 #(.width(width)) rd_st10_1676  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1676]), .rdlo_in(a10_wr[1677]),  .coef_in(coef[0]), .rdup_out(a11_wr[1676]), .rdlo_out(a11_wr[1677]));
			radix2 #(.width(width)) rd_st10_1678  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1678]), .rdlo_in(a10_wr[1679]),  .coef_in(coef[0]), .rdup_out(a11_wr[1678]), .rdlo_out(a11_wr[1679]));
			radix2 #(.width(width)) rd_st10_1680  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1680]), .rdlo_in(a10_wr[1681]),  .coef_in(coef[0]), .rdup_out(a11_wr[1680]), .rdlo_out(a11_wr[1681]));
			radix2 #(.width(width)) rd_st10_1682  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1682]), .rdlo_in(a10_wr[1683]),  .coef_in(coef[0]), .rdup_out(a11_wr[1682]), .rdlo_out(a11_wr[1683]));
			radix2 #(.width(width)) rd_st10_1684  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1684]), .rdlo_in(a10_wr[1685]),  .coef_in(coef[0]), .rdup_out(a11_wr[1684]), .rdlo_out(a11_wr[1685]));
			radix2 #(.width(width)) rd_st10_1686  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1686]), .rdlo_in(a10_wr[1687]),  .coef_in(coef[0]), .rdup_out(a11_wr[1686]), .rdlo_out(a11_wr[1687]));
			radix2 #(.width(width)) rd_st10_1688  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1688]), .rdlo_in(a10_wr[1689]),  .coef_in(coef[0]), .rdup_out(a11_wr[1688]), .rdlo_out(a11_wr[1689]));
			radix2 #(.width(width)) rd_st10_1690  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1690]), .rdlo_in(a10_wr[1691]),  .coef_in(coef[0]), .rdup_out(a11_wr[1690]), .rdlo_out(a11_wr[1691]));
			radix2 #(.width(width)) rd_st10_1692  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1692]), .rdlo_in(a10_wr[1693]),  .coef_in(coef[0]), .rdup_out(a11_wr[1692]), .rdlo_out(a11_wr[1693]));
			radix2 #(.width(width)) rd_st10_1694  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1694]), .rdlo_in(a10_wr[1695]),  .coef_in(coef[0]), .rdup_out(a11_wr[1694]), .rdlo_out(a11_wr[1695]));
			radix2 #(.width(width)) rd_st10_1696  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1696]), .rdlo_in(a10_wr[1697]),  .coef_in(coef[0]), .rdup_out(a11_wr[1696]), .rdlo_out(a11_wr[1697]));
			radix2 #(.width(width)) rd_st10_1698  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1698]), .rdlo_in(a10_wr[1699]),  .coef_in(coef[0]), .rdup_out(a11_wr[1698]), .rdlo_out(a11_wr[1699]));
			radix2 #(.width(width)) rd_st10_1700  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1700]), .rdlo_in(a10_wr[1701]),  .coef_in(coef[0]), .rdup_out(a11_wr[1700]), .rdlo_out(a11_wr[1701]));
			radix2 #(.width(width)) rd_st10_1702  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1702]), .rdlo_in(a10_wr[1703]),  .coef_in(coef[0]), .rdup_out(a11_wr[1702]), .rdlo_out(a11_wr[1703]));
			radix2 #(.width(width)) rd_st10_1704  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1704]), .rdlo_in(a10_wr[1705]),  .coef_in(coef[0]), .rdup_out(a11_wr[1704]), .rdlo_out(a11_wr[1705]));
			radix2 #(.width(width)) rd_st10_1706  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1706]), .rdlo_in(a10_wr[1707]),  .coef_in(coef[0]), .rdup_out(a11_wr[1706]), .rdlo_out(a11_wr[1707]));
			radix2 #(.width(width)) rd_st10_1708  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1708]), .rdlo_in(a10_wr[1709]),  .coef_in(coef[0]), .rdup_out(a11_wr[1708]), .rdlo_out(a11_wr[1709]));
			radix2 #(.width(width)) rd_st10_1710  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1710]), .rdlo_in(a10_wr[1711]),  .coef_in(coef[0]), .rdup_out(a11_wr[1710]), .rdlo_out(a11_wr[1711]));
			radix2 #(.width(width)) rd_st10_1712  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1712]), .rdlo_in(a10_wr[1713]),  .coef_in(coef[0]), .rdup_out(a11_wr[1712]), .rdlo_out(a11_wr[1713]));
			radix2 #(.width(width)) rd_st10_1714  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1714]), .rdlo_in(a10_wr[1715]),  .coef_in(coef[0]), .rdup_out(a11_wr[1714]), .rdlo_out(a11_wr[1715]));
			radix2 #(.width(width)) rd_st10_1716  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1716]), .rdlo_in(a10_wr[1717]),  .coef_in(coef[0]), .rdup_out(a11_wr[1716]), .rdlo_out(a11_wr[1717]));
			radix2 #(.width(width)) rd_st10_1718  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1718]), .rdlo_in(a10_wr[1719]),  .coef_in(coef[0]), .rdup_out(a11_wr[1718]), .rdlo_out(a11_wr[1719]));
			radix2 #(.width(width)) rd_st10_1720  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1720]), .rdlo_in(a10_wr[1721]),  .coef_in(coef[0]), .rdup_out(a11_wr[1720]), .rdlo_out(a11_wr[1721]));
			radix2 #(.width(width)) rd_st10_1722  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1722]), .rdlo_in(a10_wr[1723]),  .coef_in(coef[0]), .rdup_out(a11_wr[1722]), .rdlo_out(a11_wr[1723]));
			radix2 #(.width(width)) rd_st10_1724  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1724]), .rdlo_in(a10_wr[1725]),  .coef_in(coef[0]), .rdup_out(a11_wr[1724]), .rdlo_out(a11_wr[1725]));
			radix2 #(.width(width)) rd_st10_1726  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1726]), .rdlo_in(a10_wr[1727]),  .coef_in(coef[0]), .rdup_out(a11_wr[1726]), .rdlo_out(a11_wr[1727]));
			radix2 #(.width(width)) rd_st10_1728  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1728]), .rdlo_in(a10_wr[1729]),  .coef_in(coef[0]), .rdup_out(a11_wr[1728]), .rdlo_out(a11_wr[1729]));
			radix2 #(.width(width)) rd_st10_1730  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1730]), .rdlo_in(a10_wr[1731]),  .coef_in(coef[0]), .rdup_out(a11_wr[1730]), .rdlo_out(a11_wr[1731]));
			radix2 #(.width(width)) rd_st10_1732  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1732]), .rdlo_in(a10_wr[1733]),  .coef_in(coef[0]), .rdup_out(a11_wr[1732]), .rdlo_out(a11_wr[1733]));
			radix2 #(.width(width)) rd_st10_1734  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1734]), .rdlo_in(a10_wr[1735]),  .coef_in(coef[0]), .rdup_out(a11_wr[1734]), .rdlo_out(a11_wr[1735]));
			radix2 #(.width(width)) rd_st10_1736  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1736]), .rdlo_in(a10_wr[1737]),  .coef_in(coef[0]), .rdup_out(a11_wr[1736]), .rdlo_out(a11_wr[1737]));
			radix2 #(.width(width)) rd_st10_1738  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1738]), .rdlo_in(a10_wr[1739]),  .coef_in(coef[0]), .rdup_out(a11_wr[1738]), .rdlo_out(a11_wr[1739]));
			radix2 #(.width(width)) rd_st10_1740  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1740]), .rdlo_in(a10_wr[1741]),  .coef_in(coef[0]), .rdup_out(a11_wr[1740]), .rdlo_out(a11_wr[1741]));
			radix2 #(.width(width)) rd_st10_1742  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1742]), .rdlo_in(a10_wr[1743]),  .coef_in(coef[0]), .rdup_out(a11_wr[1742]), .rdlo_out(a11_wr[1743]));
			radix2 #(.width(width)) rd_st10_1744  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1744]), .rdlo_in(a10_wr[1745]),  .coef_in(coef[0]), .rdup_out(a11_wr[1744]), .rdlo_out(a11_wr[1745]));
			radix2 #(.width(width)) rd_st10_1746  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1746]), .rdlo_in(a10_wr[1747]),  .coef_in(coef[0]), .rdup_out(a11_wr[1746]), .rdlo_out(a11_wr[1747]));
			radix2 #(.width(width)) rd_st10_1748  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1748]), .rdlo_in(a10_wr[1749]),  .coef_in(coef[0]), .rdup_out(a11_wr[1748]), .rdlo_out(a11_wr[1749]));
			radix2 #(.width(width)) rd_st10_1750  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1750]), .rdlo_in(a10_wr[1751]),  .coef_in(coef[0]), .rdup_out(a11_wr[1750]), .rdlo_out(a11_wr[1751]));
			radix2 #(.width(width)) rd_st10_1752  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1752]), .rdlo_in(a10_wr[1753]),  .coef_in(coef[0]), .rdup_out(a11_wr[1752]), .rdlo_out(a11_wr[1753]));
			radix2 #(.width(width)) rd_st10_1754  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1754]), .rdlo_in(a10_wr[1755]),  .coef_in(coef[0]), .rdup_out(a11_wr[1754]), .rdlo_out(a11_wr[1755]));
			radix2 #(.width(width)) rd_st10_1756  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1756]), .rdlo_in(a10_wr[1757]),  .coef_in(coef[0]), .rdup_out(a11_wr[1756]), .rdlo_out(a11_wr[1757]));
			radix2 #(.width(width)) rd_st10_1758  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1758]), .rdlo_in(a10_wr[1759]),  .coef_in(coef[0]), .rdup_out(a11_wr[1758]), .rdlo_out(a11_wr[1759]));
			radix2 #(.width(width)) rd_st10_1760  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1760]), .rdlo_in(a10_wr[1761]),  .coef_in(coef[0]), .rdup_out(a11_wr[1760]), .rdlo_out(a11_wr[1761]));
			radix2 #(.width(width)) rd_st10_1762  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1762]), .rdlo_in(a10_wr[1763]),  .coef_in(coef[0]), .rdup_out(a11_wr[1762]), .rdlo_out(a11_wr[1763]));
			radix2 #(.width(width)) rd_st10_1764  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1764]), .rdlo_in(a10_wr[1765]),  .coef_in(coef[0]), .rdup_out(a11_wr[1764]), .rdlo_out(a11_wr[1765]));
			radix2 #(.width(width)) rd_st10_1766  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1766]), .rdlo_in(a10_wr[1767]),  .coef_in(coef[0]), .rdup_out(a11_wr[1766]), .rdlo_out(a11_wr[1767]));
			radix2 #(.width(width)) rd_st10_1768  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1768]), .rdlo_in(a10_wr[1769]),  .coef_in(coef[0]), .rdup_out(a11_wr[1768]), .rdlo_out(a11_wr[1769]));
			radix2 #(.width(width)) rd_st10_1770  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1770]), .rdlo_in(a10_wr[1771]),  .coef_in(coef[0]), .rdup_out(a11_wr[1770]), .rdlo_out(a11_wr[1771]));
			radix2 #(.width(width)) rd_st10_1772  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1772]), .rdlo_in(a10_wr[1773]),  .coef_in(coef[0]), .rdup_out(a11_wr[1772]), .rdlo_out(a11_wr[1773]));
			radix2 #(.width(width)) rd_st10_1774  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1774]), .rdlo_in(a10_wr[1775]),  .coef_in(coef[0]), .rdup_out(a11_wr[1774]), .rdlo_out(a11_wr[1775]));
			radix2 #(.width(width)) rd_st10_1776  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1776]), .rdlo_in(a10_wr[1777]),  .coef_in(coef[0]), .rdup_out(a11_wr[1776]), .rdlo_out(a11_wr[1777]));
			radix2 #(.width(width)) rd_st10_1778  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1778]), .rdlo_in(a10_wr[1779]),  .coef_in(coef[0]), .rdup_out(a11_wr[1778]), .rdlo_out(a11_wr[1779]));
			radix2 #(.width(width)) rd_st10_1780  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1780]), .rdlo_in(a10_wr[1781]),  .coef_in(coef[0]), .rdup_out(a11_wr[1780]), .rdlo_out(a11_wr[1781]));
			radix2 #(.width(width)) rd_st10_1782  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1782]), .rdlo_in(a10_wr[1783]),  .coef_in(coef[0]), .rdup_out(a11_wr[1782]), .rdlo_out(a11_wr[1783]));
			radix2 #(.width(width)) rd_st10_1784  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1784]), .rdlo_in(a10_wr[1785]),  .coef_in(coef[0]), .rdup_out(a11_wr[1784]), .rdlo_out(a11_wr[1785]));
			radix2 #(.width(width)) rd_st10_1786  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1786]), .rdlo_in(a10_wr[1787]),  .coef_in(coef[0]), .rdup_out(a11_wr[1786]), .rdlo_out(a11_wr[1787]));
			radix2 #(.width(width)) rd_st10_1788  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1788]), .rdlo_in(a10_wr[1789]),  .coef_in(coef[0]), .rdup_out(a11_wr[1788]), .rdlo_out(a11_wr[1789]));
			radix2 #(.width(width)) rd_st10_1790  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1790]), .rdlo_in(a10_wr[1791]),  .coef_in(coef[0]), .rdup_out(a11_wr[1790]), .rdlo_out(a11_wr[1791]));
			radix2 #(.width(width)) rd_st10_1792  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1792]), .rdlo_in(a10_wr[1793]),  .coef_in(coef[0]), .rdup_out(a11_wr[1792]), .rdlo_out(a11_wr[1793]));
			radix2 #(.width(width)) rd_st10_1794  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1794]), .rdlo_in(a10_wr[1795]),  .coef_in(coef[0]), .rdup_out(a11_wr[1794]), .rdlo_out(a11_wr[1795]));
			radix2 #(.width(width)) rd_st10_1796  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1796]), .rdlo_in(a10_wr[1797]),  .coef_in(coef[0]), .rdup_out(a11_wr[1796]), .rdlo_out(a11_wr[1797]));
			radix2 #(.width(width)) rd_st10_1798  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1798]), .rdlo_in(a10_wr[1799]),  .coef_in(coef[0]), .rdup_out(a11_wr[1798]), .rdlo_out(a11_wr[1799]));
			radix2 #(.width(width)) rd_st10_1800  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1800]), .rdlo_in(a10_wr[1801]),  .coef_in(coef[0]), .rdup_out(a11_wr[1800]), .rdlo_out(a11_wr[1801]));
			radix2 #(.width(width)) rd_st10_1802  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1802]), .rdlo_in(a10_wr[1803]),  .coef_in(coef[0]), .rdup_out(a11_wr[1802]), .rdlo_out(a11_wr[1803]));
			radix2 #(.width(width)) rd_st10_1804  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1804]), .rdlo_in(a10_wr[1805]),  .coef_in(coef[0]), .rdup_out(a11_wr[1804]), .rdlo_out(a11_wr[1805]));
			radix2 #(.width(width)) rd_st10_1806  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1806]), .rdlo_in(a10_wr[1807]),  .coef_in(coef[0]), .rdup_out(a11_wr[1806]), .rdlo_out(a11_wr[1807]));
			radix2 #(.width(width)) rd_st10_1808  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1808]), .rdlo_in(a10_wr[1809]),  .coef_in(coef[0]), .rdup_out(a11_wr[1808]), .rdlo_out(a11_wr[1809]));
			radix2 #(.width(width)) rd_st10_1810  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1810]), .rdlo_in(a10_wr[1811]),  .coef_in(coef[0]), .rdup_out(a11_wr[1810]), .rdlo_out(a11_wr[1811]));
			radix2 #(.width(width)) rd_st10_1812  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1812]), .rdlo_in(a10_wr[1813]),  .coef_in(coef[0]), .rdup_out(a11_wr[1812]), .rdlo_out(a11_wr[1813]));
			radix2 #(.width(width)) rd_st10_1814  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1814]), .rdlo_in(a10_wr[1815]),  .coef_in(coef[0]), .rdup_out(a11_wr[1814]), .rdlo_out(a11_wr[1815]));
			radix2 #(.width(width)) rd_st10_1816  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1816]), .rdlo_in(a10_wr[1817]),  .coef_in(coef[0]), .rdup_out(a11_wr[1816]), .rdlo_out(a11_wr[1817]));
			radix2 #(.width(width)) rd_st10_1818  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1818]), .rdlo_in(a10_wr[1819]),  .coef_in(coef[0]), .rdup_out(a11_wr[1818]), .rdlo_out(a11_wr[1819]));
			radix2 #(.width(width)) rd_st10_1820  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1820]), .rdlo_in(a10_wr[1821]),  .coef_in(coef[0]), .rdup_out(a11_wr[1820]), .rdlo_out(a11_wr[1821]));
			radix2 #(.width(width)) rd_st10_1822  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1822]), .rdlo_in(a10_wr[1823]),  .coef_in(coef[0]), .rdup_out(a11_wr[1822]), .rdlo_out(a11_wr[1823]));
			radix2 #(.width(width)) rd_st10_1824  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1824]), .rdlo_in(a10_wr[1825]),  .coef_in(coef[0]), .rdup_out(a11_wr[1824]), .rdlo_out(a11_wr[1825]));
			radix2 #(.width(width)) rd_st10_1826  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1826]), .rdlo_in(a10_wr[1827]),  .coef_in(coef[0]), .rdup_out(a11_wr[1826]), .rdlo_out(a11_wr[1827]));
			radix2 #(.width(width)) rd_st10_1828  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1828]), .rdlo_in(a10_wr[1829]),  .coef_in(coef[0]), .rdup_out(a11_wr[1828]), .rdlo_out(a11_wr[1829]));
			radix2 #(.width(width)) rd_st10_1830  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1830]), .rdlo_in(a10_wr[1831]),  .coef_in(coef[0]), .rdup_out(a11_wr[1830]), .rdlo_out(a11_wr[1831]));
			radix2 #(.width(width)) rd_st10_1832  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1832]), .rdlo_in(a10_wr[1833]),  .coef_in(coef[0]), .rdup_out(a11_wr[1832]), .rdlo_out(a11_wr[1833]));
			radix2 #(.width(width)) rd_st10_1834  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1834]), .rdlo_in(a10_wr[1835]),  .coef_in(coef[0]), .rdup_out(a11_wr[1834]), .rdlo_out(a11_wr[1835]));
			radix2 #(.width(width)) rd_st10_1836  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1836]), .rdlo_in(a10_wr[1837]),  .coef_in(coef[0]), .rdup_out(a11_wr[1836]), .rdlo_out(a11_wr[1837]));
			radix2 #(.width(width)) rd_st10_1838  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1838]), .rdlo_in(a10_wr[1839]),  .coef_in(coef[0]), .rdup_out(a11_wr[1838]), .rdlo_out(a11_wr[1839]));
			radix2 #(.width(width)) rd_st10_1840  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1840]), .rdlo_in(a10_wr[1841]),  .coef_in(coef[0]), .rdup_out(a11_wr[1840]), .rdlo_out(a11_wr[1841]));
			radix2 #(.width(width)) rd_st10_1842  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1842]), .rdlo_in(a10_wr[1843]),  .coef_in(coef[0]), .rdup_out(a11_wr[1842]), .rdlo_out(a11_wr[1843]));
			radix2 #(.width(width)) rd_st10_1844  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1844]), .rdlo_in(a10_wr[1845]),  .coef_in(coef[0]), .rdup_out(a11_wr[1844]), .rdlo_out(a11_wr[1845]));
			radix2 #(.width(width)) rd_st10_1846  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1846]), .rdlo_in(a10_wr[1847]),  .coef_in(coef[0]), .rdup_out(a11_wr[1846]), .rdlo_out(a11_wr[1847]));
			radix2 #(.width(width)) rd_st10_1848  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1848]), .rdlo_in(a10_wr[1849]),  .coef_in(coef[0]), .rdup_out(a11_wr[1848]), .rdlo_out(a11_wr[1849]));
			radix2 #(.width(width)) rd_st10_1850  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1850]), .rdlo_in(a10_wr[1851]),  .coef_in(coef[0]), .rdup_out(a11_wr[1850]), .rdlo_out(a11_wr[1851]));
			radix2 #(.width(width)) rd_st10_1852  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1852]), .rdlo_in(a10_wr[1853]),  .coef_in(coef[0]), .rdup_out(a11_wr[1852]), .rdlo_out(a11_wr[1853]));
			radix2 #(.width(width)) rd_st10_1854  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1854]), .rdlo_in(a10_wr[1855]),  .coef_in(coef[0]), .rdup_out(a11_wr[1854]), .rdlo_out(a11_wr[1855]));
			radix2 #(.width(width)) rd_st10_1856  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1856]), .rdlo_in(a10_wr[1857]),  .coef_in(coef[0]), .rdup_out(a11_wr[1856]), .rdlo_out(a11_wr[1857]));
			radix2 #(.width(width)) rd_st10_1858  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1858]), .rdlo_in(a10_wr[1859]),  .coef_in(coef[0]), .rdup_out(a11_wr[1858]), .rdlo_out(a11_wr[1859]));
			radix2 #(.width(width)) rd_st10_1860  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1860]), .rdlo_in(a10_wr[1861]),  .coef_in(coef[0]), .rdup_out(a11_wr[1860]), .rdlo_out(a11_wr[1861]));
			radix2 #(.width(width)) rd_st10_1862  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1862]), .rdlo_in(a10_wr[1863]),  .coef_in(coef[0]), .rdup_out(a11_wr[1862]), .rdlo_out(a11_wr[1863]));
			radix2 #(.width(width)) rd_st10_1864  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1864]), .rdlo_in(a10_wr[1865]),  .coef_in(coef[0]), .rdup_out(a11_wr[1864]), .rdlo_out(a11_wr[1865]));
			radix2 #(.width(width)) rd_st10_1866  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1866]), .rdlo_in(a10_wr[1867]),  .coef_in(coef[0]), .rdup_out(a11_wr[1866]), .rdlo_out(a11_wr[1867]));
			radix2 #(.width(width)) rd_st10_1868  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1868]), .rdlo_in(a10_wr[1869]),  .coef_in(coef[0]), .rdup_out(a11_wr[1868]), .rdlo_out(a11_wr[1869]));
			radix2 #(.width(width)) rd_st10_1870  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1870]), .rdlo_in(a10_wr[1871]),  .coef_in(coef[0]), .rdup_out(a11_wr[1870]), .rdlo_out(a11_wr[1871]));
			radix2 #(.width(width)) rd_st10_1872  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1872]), .rdlo_in(a10_wr[1873]),  .coef_in(coef[0]), .rdup_out(a11_wr[1872]), .rdlo_out(a11_wr[1873]));
			radix2 #(.width(width)) rd_st10_1874  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1874]), .rdlo_in(a10_wr[1875]),  .coef_in(coef[0]), .rdup_out(a11_wr[1874]), .rdlo_out(a11_wr[1875]));
			radix2 #(.width(width)) rd_st10_1876  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1876]), .rdlo_in(a10_wr[1877]),  .coef_in(coef[0]), .rdup_out(a11_wr[1876]), .rdlo_out(a11_wr[1877]));
			radix2 #(.width(width)) rd_st10_1878  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1878]), .rdlo_in(a10_wr[1879]),  .coef_in(coef[0]), .rdup_out(a11_wr[1878]), .rdlo_out(a11_wr[1879]));
			radix2 #(.width(width)) rd_st10_1880  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1880]), .rdlo_in(a10_wr[1881]),  .coef_in(coef[0]), .rdup_out(a11_wr[1880]), .rdlo_out(a11_wr[1881]));
			radix2 #(.width(width)) rd_st10_1882  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1882]), .rdlo_in(a10_wr[1883]),  .coef_in(coef[0]), .rdup_out(a11_wr[1882]), .rdlo_out(a11_wr[1883]));
			radix2 #(.width(width)) rd_st10_1884  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1884]), .rdlo_in(a10_wr[1885]),  .coef_in(coef[0]), .rdup_out(a11_wr[1884]), .rdlo_out(a11_wr[1885]));
			radix2 #(.width(width)) rd_st10_1886  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1886]), .rdlo_in(a10_wr[1887]),  .coef_in(coef[0]), .rdup_out(a11_wr[1886]), .rdlo_out(a11_wr[1887]));
			radix2 #(.width(width)) rd_st10_1888  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1888]), .rdlo_in(a10_wr[1889]),  .coef_in(coef[0]), .rdup_out(a11_wr[1888]), .rdlo_out(a11_wr[1889]));
			radix2 #(.width(width)) rd_st10_1890  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1890]), .rdlo_in(a10_wr[1891]),  .coef_in(coef[0]), .rdup_out(a11_wr[1890]), .rdlo_out(a11_wr[1891]));
			radix2 #(.width(width)) rd_st10_1892  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1892]), .rdlo_in(a10_wr[1893]),  .coef_in(coef[0]), .rdup_out(a11_wr[1892]), .rdlo_out(a11_wr[1893]));
			radix2 #(.width(width)) rd_st10_1894  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1894]), .rdlo_in(a10_wr[1895]),  .coef_in(coef[0]), .rdup_out(a11_wr[1894]), .rdlo_out(a11_wr[1895]));
			radix2 #(.width(width)) rd_st10_1896  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1896]), .rdlo_in(a10_wr[1897]),  .coef_in(coef[0]), .rdup_out(a11_wr[1896]), .rdlo_out(a11_wr[1897]));
			radix2 #(.width(width)) rd_st10_1898  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1898]), .rdlo_in(a10_wr[1899]),  .coef_in(coef[0]), .rdup_out(a11_wr[1898]), .rdlo_out(a11_wr[1899]));
			radix2 #(.width(width)) rd_st10_1900  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1900]), .rdlo_in(a10_wr[1901]),  .coef_in(coef[0]), .rdup_out(a11_wr[1900]), .rdlo_out(a11_wr[1901]));
			radix2 #(.width(width)) rd_st10_1902  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1902]), .rdlo_in(a10_wr[1903]),  .coef_in(coef[0]), .rdup_out(a11_wr[1902]), .rdlo_out(a11_wr[1903]));
			radix2 #(.width(width)) rd_st10_1904  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1904]), .rdlo_in(a10_wr[1905]),  .coef_in(coef[0]), .rdup_out(a11_wr[1904]), .rdlo_out(a11_wr[1905]));
			radix2 #(.width(width)) rd_st10_1906  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1906]), .rdlo_in(a10_wr[1907]),  .coef_in(coef[0]), .rdup_out(a11_wr[1906]), .rdlo_out(a11_wr[1907]));
			radix2 #(.width(width)) rd_st10_1908  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1908]), .rdlo_in(a10_wr[1909]),  .coef_in(coef[0]), .rdup_out(a11_wr[1908]), .rdlo_out(a11_wr[1909]));
			radix2 #(.width(width)) rd_st10_1910  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1910]), .rdlo_in(a10_wr[1911]),  .coef_in(coef[0]), .rdup_out(a11_wr[1910]), .rdlo_out(a11_wr[1911]));
			radix2 #(.width(width)) rd_st10_1912  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1912]), .rdlo_in(a10_wr[1913]),  .coef_in(coef[0]), .rdup_out(a11_wr[1912]), .rdlo_out(a11_wr[1913]));
			radix2 #(.width(width)) rd_st10_1914  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1914]), .rdlo_in(a10_wr[1915]),  .coef_in(coef[0]), .rdup_out(a11_wr[1914]), .rdlo_out(a11_wr[1915]));
			radix2 #(.width(width)) rd_st10_1916  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1916]), .rdlo_in(a10_wr[1917]),  .coef_in(coef[0]), .rdup_out(a11_wr[1916]), .rdlo_out(a11_wr[1917]));
			radix2 #(.width(width)) rd_st10_1918  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1918]), .rdlo_in(a10_wr[1919]),  .coef_in(coef[0]), .rdup_out(a11_wr[1918]), .rdlo_out(a11_wr[1919]));
			radix2 #(.width(width)) rd_st10_1920  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1920]), .rdlo_in(a10_wr[1921]),  .coef_in(coef[0]), .rdup_out(a11_wr[1920]), .rdlo_out(a11_wr[1921]));
			radix2 #(.width(width)) rd_st10_1922  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1922]), .rdlo_in(a10_wr[1923]),  .coef_in(coef[0]), .rdup_out(a11_wr[1922]), .rdlo_out(a11_wr[1923]));
			radix2 #(.width(width)) rd_st10_1924  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1924]), .rdlo_in(a10_wr[1925]),  .coef_in(coef[0]), .rdup_out(a11_wr[1924]), .rdlo_out(a11_wr[1925]));
			radix2 #(.width(width)) rd_st10_1926  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1926]), .rdlo_in(a10_wr[1927]),  .coef_in(coef[0]), .rdup_out(a11_wr[1926]), .rdlo_out(a11_wr[1927]));
			radix2 #(.width(width)) rd_st10_1928  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1928]), .rdlo_in(a10_wr[1929]),  .coef_in(coef[0]), .rdup_out(a11_wr[1928]), .rdlo_out(a11_wr[1929]));
			radix2 #(.width(width)) rd_st10_1930  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1930]), .rdlo_in(a10_wr[1931]),  .coef_in(coef[0]), .rdup_out(a11_wr[1930]), .rdlo_out(a11_wr[1931]));
			radix2 #(.width(width)) rd_st10_1932  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1932]), .rdlo_in(a10_wr[1933]),  .coef_in(coef[0]), .rdup_out(a11_wr[1932]), .rdlo_out(a11_wr[1933]));
			radix2 #(.width(width)) rd_st10_1934  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1934]), .rdlo_in(a10_wr[1935]),  .coef_in(coef[0]), .rdup_out(a11_wr[1934]), .rdlo_out(a11_wr[1935]));
			radix2 #(.width(width)) rd_st10_1936  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1936]), .rdlo_in(a10_wr[1937]),  .coef_in(coef[0]), .rdup_out(a11_wr[1936]), .rdlo_out(a11_wr[1937]));
			radix2 #(.width(width)) rd_st10_1938  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1938]), .rdlo_in(a10_wr[1939]),  .coef_in(coef[0]), .rdup_out(a11_wr[1938]), .rdlo_out(a11_wr[1939]));
			radix2 #(.width(width)) rd_st10_1940  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1940]), .rdlo_in(a10_wr[1941]),  .coef_in(coef[0]), .rdup_out(a11_wr[1940]), .rdlo_out(a11_wr[1941]));
			radix2 #(.width(width)) rd_st10_1942  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1942]), .rdlo_in(a10_wr[1943]),  .coef_in(coef[0]), .rdup_out(a11_wr[1942]), .rdlo_out(a11_wr[1943]));
			radix2 #(.width(width)) rd_st10_1944  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1944]), .rdlo_in(a10_wr[1945]),  .coef_in(coef[0]), .rdup_out(a11_wr[1944]), .rdlo_out(a11_wr[1945]));
			radix2 #(.width(width)) rd_st10_1946  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1946]), .rdlo_in(a10_wr[1947]),  .coef_in(coef[0]), .rdup_out(a11_wr[1946]), .rdlo_out(a11_wr[1947]));
			radix2 #(.width(width)) rd_st10_1948  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1948]), .rdlo_in(a10_wr[1949]),  .coef_in(coef[0]), .rdup_out(a11_wr[1948]), .rdlo_out(a11_wr[1949]));
			radix2 #(.width(width)) rd_st10_1950  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1950]), .rdlo_in(a10_wr[1951]),  .coef_in(coef[0]), .rdup_out(a11_wr[1950]), .rdlo_out(a11_wr[1951]));
			radix2 #(.width(width)) rd_st10_1952  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1952]), .rdlo_in(a10_wr[1953]),  .coef_in(coef[0]), .rdup_out(a11_wr[1952]), .rdlo_out(a11_wr[1953]));
			radix2 #(.width(width)) rd_st10_1954  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1954]), .rdlo_in(a10_wr[1955]),  .coef_in(coef[0]), .rdup_out(a11_wr[1954]), .rdlo_out(a11_wr[1955]));
			radix2 #(.width(width)) rd_st10_1956  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1956]), .rdlo_in(a10_wr[1957]),  .coef_in(coef[0]), .rdup_out(a11_wr[1956]), .rdlo_out(a11_wr[1957]));
			radix2 #(.width(width)) rd_st10_1958  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1958]), .rdlo_in(a10_wr[1959]),  .coef_in(coef[0]), .rdup_out(a11_wr[1958]), .rdlo_out(a11_wr[1959]));
			radix2 #(.width(width)) rd_st10_1960  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1960]), .rdlo_in(a10_wr[1961]),  .coef_in(coef[0]), .rdup_out(a11_wr[1960]), .rdlo_out(a11_wr[1961]));
			radix2 #(.width(width)) rd_st10_1962  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1962]), .rdlo_in(a10_wr[1963]),  .coef_in(coef[0]), .rdup_out(a11_wr[1962]), .rdlo_out(a11_wr[1963]));
			radix2 #(.width(width)) rd_st10_1964  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1964]), .rdlo_in(a10_wr[1965]),  .coef_in(coef[0]), .rdup_out(a11_wr[1964]), .rdlo_out(a11_wr[1965]));
			radix2 #(.width(width)) rd_st10_1966  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1966]), .rdlo_in(a10_wr[1967]),  .coef_in(coef[0]), .rdup_out(a11_wr[1966]), .rdlo_out(a11_wr[1967]));
			radix2 #(.width(width)) rd_st10_1968  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1968]), .rdlo_in(a10_wr[1969]),  .coef_in(coef[0]), .rdup_out(a11_wr[1968]), .rdlo_out(a11_wr[1969]));
			radix2 #(.width(width)) rd_st10_1970  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1970]), .rdlo_in(a10_wr[1971]),  .coef_in(coef[0]), .rdup_out(a11_wr[1970]), .rdlo_out(a11_wr[1971]));
			radix2 #(.width(width)) rd_st10_1972  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1972]), .rdlo_in(a10_wr[1973]),  .coef_in(coef[0]), .rdup_out(a11_wr[1972]), .rdlo_out(a11_wr[1973]));
			radix2 #(.width(width)) rd_st10_1974  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1974]), .rdlo_in(a10_wr[1975]),  .coef_in(coef[0]), .rdup_out(a11_wr[1974]), .rdlo_out(a11_wr[1975]));
			radix2 #(.width(width)) rd_st10_1976  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1976]), .rdlo_in(a10_wr[1977]),  .coef_in(coef[0]), .rdup_out(a11_wr[1976]), .rdlo_out(a11_wr[1977]));
			radix2 #(.width(width)) rd_st10_1978  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1978]), .rdlo_in(a10_wr[1979]),  .coef_in(coef[0]), .rdup_out(a11_wr[1978]), .rdlo_out(a11_wr[1979]));
			radix2 #(.width(width)) rd_st10_1980  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1980]), .rdlo_in(a10_wr[1981]),  .coef_in(coef[0]), .rdup_out(a11_wr[1980]), .rdlo_out(a11_wr[1981]));
			radix2 #(.width(width)) rd_st10_1982  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1982]), .rdlo_in(a10_wr[1983]),  .coef_in(coef[0]), .rdup_out(a11_wr[1982]), .rdlo_out(a11_wr[1983]));
			radix2 #(.width(width)) rd_st10_1984  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1984]), .rdlo_in(a10_wr[1985]),  .coef_in(coef[0]), .rdup_out(a11_wr[1984]), .rdlo_out(a11_wr[1985]));
			radix2 #(.width(width)) rd_st10_1986  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1986]), .rdlo_in(a10_wr[1987]),  .coef_in(coef[0]), .rdup_out(a11_wr[1986]), .rdlo_out(a11_wr[1987]));
			radix2 #(.width(width)) rd_st10_1988  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1988]), .rdlo_in(a10_wr[1989]),  .coef_in(coef[0]), .rdup_out(a11_wr[1988]), .rdlo_out(a11_wr[1989]));
			radix2 #(.width(width)) rd_st10_1990  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1990]), .rdlo_in(a10_wr[1991]),  .coef_in(coef[0]), .rdup_out(a11_wr[1990]), .rdlo_out(a11_wr[1991]));
			radix2 #(.width(width)) rd_st10_1992  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1992]), .rdlo_in(a10_wr[1993]),  .coef_in(coef[0]), .rdup_out(a11_wr[1992]), .rdlo_out(a11_wr[1993]));
			radix2 #(.width(width)) rd_st10_1994  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1994]), .rdlo_in(a10_wr[1995]),  .coef_in(coef[0]), .rdup_out(a11_wr[1994]), .rdlo_out(a11_wr[1995]));
			radix2 #(.width(width)) rd_st10_1996  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1996]), .rdlo_in(a10_wr[1997]),  .coef_in(coef[0]), .rdup_out(a11_wr[1996]), .rdlo_out(a11_wr[1997]));
			radix2 #(.width(width)) rd_st10_1998  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[1998]), .rdlo_in(a10_wr[1999]),  .coef_in(coef[0]), .rdup_out(a11_wr[1998]), .rdlo_out(a11_wr[1999]));
			radix2 #(.width(width)) rd_st10_2000  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[2000]), .rdlo_in(a10_wr[2001]),  .coef_in(coef[0]), .rdup_out(a11_wr[2000]), .rdlo_out(a11_wr[2001]));
			radix2 #(.width(width)) rd_st10_2002  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[2002]), .rdlo_in(a10_wr[2003]),  .coef_in(coef[0]), .rdup_out(a11_wr[2002]), .rdlo_out(a11_wr[2003]));
			radix2 #(.width(width)) rd_st10_2004  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[2004]), .rdlo_in(a10_wr[2005]),  .coef_in(coef[0]), .rdup_out(a11_wr[2004]), .rdlo_out(a11_wr[2005]));
			radix2 #(.width(width)) rd_st10_2006  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[2006]), .rdlo_in(a10_wr[2007]),  .coef_in(coef[0]), .rdup_out(a11_wr[2006]), .rdlo_out(a11_wr[2007]));
			radix2 #(.width(width)) rd_st10_2008  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[2008]), .rdlo_in(a10_wr[2009]),  .coef_in(coef[0]), .rdup_out(a11_wr[2008]), .rdlo_out(a11_wr[2009]));
			radix2 #(.width(width)) rd_st10_2010  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[2010]), .rdlo_in(a10_wr[2011]),  .coef_in(coef[0]), .rdup_out(a11_wr[2010]), .rdlo_out(a11_wr[2011]));
			radix2 #(.width(width)) rd_st10_2012  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[2012]), .rdlo_in(a10_wr[2013]),  .coef_in(coef[0]), .rdup_out(a11_wr[2012]), .rdlo_out(a11_wr[2013]));
			radix2 #(.width(width)) rd_st10_2014  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[2014]), .rdlo_in(a10_wr[2015]),  .coef_in(coef[0]), .rdup_out(a11_wr[2014]), .rdlo_out(a11_wr[2015]));
			radix2 #(.width(width)) rd_st10_2016  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[2016]), .rdlo_in(a10_wr[2017]),  .coef_in(coef[0]), .rdup_out(a11_wr[2016]), .rdlo_out(a11_wr[2017]));
			radix2 #(.width(width)) rd_st10_2018  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[2018]), .rdlo_in(a10_wr[2019]),  .coef_in(coef[0]), .rdup_out(a11_wr[2018]), .rdlo_out(a11_wr[2019]));
			radix2 #(.width(width)) rd_st10_2020  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[2020]), .rdlo_in(a10_wr[2021]),  .coef_in(coef[0]), .rdup_out(a11_wr[2020]), .rdlo_out(a11_wr[2021]));
			radix2 #(.width(width)) rd_st10_2022  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[2022]), .rdlo_in(a10_wr[2023]),  .coef_in(coef[0]), .rdup_out(a11_wr[2022]), .rdlo_out(a11_wr[2023]));
			radix2 #(.width(width)) rd_st10_2024  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[2024]), .rdlo_in(a10_wr[2025]),  .coef_in(coef[0]), .rdup_out(a11_wr[2024]), .rdlo_out(a11_wr[2025]));
			radix2 #(.width(width)) rd_st10_2026  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[2026]), .rdlo_in(a10_wr[2027]),  .coef_in(coef[0]), .rdup_out(a11_wr[2026]), .rdlo_out(a11_wr[2027]));
			radix2 #(.width(width)) rd_st10_2028  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[2028]), .rdlo_in(a10_wr[2029]),  .coef_in(coef[0]), .rdup_out(a11_wr[2028]), .rdlo_out(a11_wr[2029]));
			radix2 #(.width(width)) rd_st10_2030  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[2030]), .rdlo_in(a10_wr[2031]),  .coef_in(coef[0]), .rdup_out(a11_wr[2030]), .rdlo_out(a11_wr[2031]));
			radix2 #(.width(width)) rd_st10_2032  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[2032]), .rdlo_in(a10_wr[2033]),  .coef_in(coef[0]), .rdup_out(a11_wr[2032]), .rdlo_out(a11_wr[2033]));
			radix2 #(.width(width)) rd_st10_2034  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[2034]), .rdlo_in(a10_wr[2035]),  .coef_in(coef[0]), .rdup_out(a11_wr[2034]), .rdlo_out(a11_wr[2035]));
			radix2 #(.width(width)) rd_st10_2036  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[2036]), .rdlo_in(a10_wr[2037]),  .coef_in(coef[0]), .rdup_out(a11_wr[2036]), .rdlo_out(a11_wr[2037]));
			radix2 #(.width(width)) rd_st10_2038  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[2038]), .rdlo_in(a10_wr[2039]),  .coef_in(coef[0]), .rdup_out(a11_wr[2038]), .rdlo_out(a11_wr[2039]));
			radix2 #(.width(width)) rd_st10_2040  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[2040]), .rdlo_in(a10_wr[2041]),  .coef_in(coef[0]), .rdup_out(a11_wr[2040]), .rdlo_out(a11_wr[2041]));
			radix2 #(.width(width)) rd_st10_2042  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[2042]), .rdlo_in(a10_wr[2043]),  .coef_in(coef[0]), .rdup_out(a11_wr[2042]), .rdlo_out(a11_wr[2043]));
			radix2 #(.width(width)) rd_st10_2044  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[2044]), .rdlo_in(a10_wr[2045]),  .coef_in(coef[0]), .rdup_out(a11_wr[2044]), .rdlo_out(a11_wr[2045]));
			radix2 #(.width(width)) rd_st10_2046  (.clk(clk), .rst(rst),  .stall(comb_stall), .rdup_in(a10_wr[2046]), .rdlo_in(a10_wr[2047]),  .coef_in(coef[0]), .rdup_out(a11_wr[2046]), .rdlo_out(a11_wr[2047]));

		//--- output stage (bit reversal)
			assign x0_out       = a11_wr[0];                   
			assign x1_out       = a11_wr[1024];                
			assign x2_out       = a11_wr[512];                 
			assign x3_out       = a11_wr[1536];                
			assign x4_out       = a11_wr[256];                 
			assign x5_out       = a11_wr[1280];                
			assign x6_out       = a11_wr[768];                 
			assign x7_out       = a11_wr[1792];                
			assign x8_out       = a11_wr[128];                 
			assign x9_out       = a11_wr[1152];                
			assign x10_out      = a11_wr[640];                 
			assign x11_out      = a11_wr[1664];                
			assign x12_out      = a11_wr[384];                 
			assign x13_out      = a11_wr[1408];                
			assign x14_out      = a11_wr[896];                 
			assign x15_out      = a11_wr[1920];                
			assign x16_out      = a11_wr[64];                  
			assign x17_out      = a11_wr[1088];                
			assign x18_out      = a11_wr[576];                 
			assign x19_out      = a11_wr[1600];                
			assign x20_out      = a11_wr[320];                 
			assign x21_out      = a11_wr[1344];                
			assign x22_out      = a11_wr[832];                 
			assign x23_out      = a11_wr[1856];                
			assign x24_out      = a11_wr[192];                 
			assign x25_out      = a11_wr[1216];                
			assign x26_out      = a11_wr[704];                 
			assign x27_out      = a11_wr[1728];                
			assign x28_out      = a11_wr[448];                 
			assign x29_out      = a11_wr[1472];                
			assign x30_out      = a11_wr[960];                 
			assign x31_out      = a11_wr[1984];                
			assign x32_out      = a11_wr[32];                  
			assign x33_out      = a11_wr[1056];                
			assign x34_out      = a11_wr[544];                 
			assign x35_out      = a11_wr[1568];                
			assign x36_out      = a11_wr[288];                 
			assign x37_out      = a11_wr[1312];                
			assign x38_out      = a11_wr[800];                 
			assign x39_out      = a11_wr[1824];                
			assign x40_out      = a11_wr[160];                 
			assign x41_out      = a11_wr[1184];                
			assign x42_out      = a11_wr[672];                 
			assign x43_out      = a11_wr[1696];                
			assign x44_out      = a11_wr[416];                 
			assign x45_out      = a11_wr[1440];                
			assign x46_out      = a11_wr[928];                 
			assign x47_out      = a11_wr[1952];                
			assign x48_out      = a11_wr[96];                  
			assign x49_out      = a11_wr[1120];                
			assign x50_out      = a11_wr[608];                 
			assign x51_out      = a11_wr[1632];                
			assign x52_out      = a11_wr[352];                 
			assign x53_out      = a11_wr[1376];                
			assign x54_out      = a11_wr[864];                 
			assign x55_out      = a11_wr[1888];                
			assign x56_out      = a11_wr[224];                 
			assign x57_out      = a11_wr[1248];                
			assign x58_out      = a11_wr[736];                 
			assign x59_out      = a11_wr[1760];                
			assign x60_out      = a11_wr[480];                 
			assign x61_out      = a11_wr[1504];                
			assign x62_out      = a11_wr[992];                 
			assign x63_out      = a11_wr[2016];                
			assign x64_out      = a11_wr[16];                  
			assign x65_out      = a11_wr[1040];                
			assign x66_out      = a11_wr[528];                 
			assign x67_out      = a11_wr[1552];                
			assign x68_out      = a11_wr[272];                 
			assign x69_out      = a11_wr[1296];                
			assign x70_out      = a11_wr[784];                 
			assign x71_out      = a11_wr[1808];                
			assign x72_out      = a11_wr[144];                 
			assign x73_out      = a11_wr[1168];                
			assign x74_out      = a11_wr[656];                 
			assign x75_out      = a11_wr[1680];                
			assign x76_out      = a11_wr[400];                 
			assign x77_out      = a11_wr[1424];                
			assign x78_out      = a11_wr[912];                 
			assign x79_out      = a11_wr[1936];                
			assign x80_out      = a11_wr[80];                  
			assign x81_out      = a11_wr[1104];                
			assign x82_out      = a11_wr[592];                 
			assign x83_out      = a11_wr[1616];                
			assign x84_out      = a11_wr[336];                 
			assign x85_out      = a11_wr[1360];                
			assign x86_out      = a11_wr[848];                 
			assign x87_out      = a11_wr[1872];                
			assign x88_out      = a11_wr[208];                 
			assign x89_out      = a11_wr[1232];                
			assign x90_out      = a11_wr[720];                 
			assign x91_out      = a11_wr[1744];                
			assign x92_out      = a11_wr[464];                 
			assign x93_out      = a11_wr[1488];                
			assign x94_out      = a11_wr[976];                 
			assign x95_out      = a11_wr[2000];                
			assign x96_out      = a11_wr[48];                  
			assign x97_out      = a11_wr[1072];                
			assign x98_out      = a11_wr[560];                 
			assign x99_out      = a11_wr[1584];                
			assign x100_out     = a11_wr[304];                 
			assign x101_out     = a11_wr[1328];                
			assign x102_out     = a11_wr[816];                 
			assign x103_out     = a11_wr[1840];                
			assign x104_out     = a11_wr[176];                 
			assign x105_out     = a11_wr[1200];                
			assign x106_out     = a11_wr[688];                 
			assign x107_out     = a11_wr[1712];                
			assign x108_out     = a11_wr[432];                 
			assign x109_out     = a11_wr[1456];                
			assign x110_out     = a11_wr[944];                 
			assign x111_out     = a11_wr[1968];                
			assign x112_out     = a11_wr[112];                 
			assign x113_out     = a11_wr[1136];                
			assign x114_out     = a11_wr[624];                 
			assign x115_out     = a11_wr[1648];                
			assign x116_out     = a11_wr[368];                 
			assign x117_out     = a11_wr[1392];                
			assign x118_out     = a11_wr[880];                 
			assign x119_out     = a11_wr[1904];                
			assign x120_out     = a11_wr[240];                 
			assign x121_out     = a11_wr[1264];                
			assign x122_out     = a11_wr[752];                 
			assign x123_out     = a11_wr[1776];                
			assign x124_out     = a11_wr[496];                 
			assign x125_out     = a11_wr[1520];                
			assign x126_out     = a11_wr[1008];                
			assign x127_out     = a11_wr[2032];                
			assign x128_out     = a11_wr[8];                   
			assign x129_out     = a11_wr[1032];                
			assign x130_out     = a11_wr[520];                 
			assign x131_out     = a11_wr[1544];                
			assign x132_out     = a11_wr[264];                 
			assign x133_out     = a11_wr[1288];                
			assign x134_out     = a11_wr[776];                 
			assign x135_out     = a11_wr[1800];                
			assign x136_out     = a11_wr[136];                 
			assign x137_out     = a11_wr[1160];                
			assign x138_out     = a11_wr[648];                 
			assign x139_out     = a11_wr[1672];                
			assign x140_out     = a11_wr[392];                 
			assign x141_out     = a11_wr[1416];                
			assign x142_out     = a11_wr[904];                 
			assign x143_out     = a11_wr[1928];                
			assign x144_out     = a11_wr[72];                  
			assign x145_out     = a11_wr[1096];                
			assign x146_out     = a11_wr[584];                 
			assign x147_out     = a11_wr[1608];                
			assign x148_out     = a11_wr[328];                 
			assign x149_out     = a11_wr[1352];                
			assign x150_out     = a11_wr[840];                 
			assign x151_out     = a11_wr[1864];                
			assign x152_out     = a11_wr[200];                 
			assign x153_out     = a11_wr[1224];                
			assign x154_out     = a11_wr[712];                 
			assign x155_out     = a11_wr[1736];                
			assign x156_out     = a11_wr[456];                 
			assign x157_out     = a11_wr[1480];                
			assign x158_out     = a11_wr[968];                 
			assign x159_out     = a11_wr[1992];                
			assign x160_out     = a11_wr[40];                  
			assign x161_out     = a11_wr[1064];                
			assign x162_out     = a11_wr[552];                 
			assign x163_out     = a11_wr[1576];                
			assign x164_out     = a11_wr[296];                 
			assign x165_out     = a11_wr[1320];                
			assign x166_out     = a11_wr[808];                 
			assign x167_out     = a11_wr[1832];                
			assign x168_out     = a11_wr[168];                 
			assign x169_out     = a11_wr[1192];                
			assign x170_out     = a11_wr[680];                 
			assign x171_out     = a11_wr[1704];                
			assign x172_out     = a11_wr[424];                 
			assign x173_out     = a11_wr[1448];                
			assign x174_out     = a11_wr[936];                 
			assign x175_out     = a11_wr[1960];                
			assign x176_out     = a11_wr[104];                 
			assign x177_out     = a11_wr[1128];                
			assign x178_out     = a11_wr[616];                 
			assign x179_out     = a11_wr[1640];                
			assign x180_out     = a11_wr[360];                 
			assign x181_out     = a11_wr[1384];                
			assign x182_out     = a11_wr[872];                 
			assign x183_out     = a11_wr[1896];                
			assign x184_out     = a11_wr[232];                 
			assign x185_out     = a11_wr[1256];                
			assign x186_out     = a11_wr[744];                 
			assign x187_out     = a11_wr[1768];                
			assign x188_out     = a11_wr[488];                 
			assign x189_out     = a11_wr[1512];                
			assign x190_out     = a11_wr[1000];                
			assign x191_out     = a11_wr[2024];                
			assign x192_out     = a11_wr[24];                  
			assign x193_out     = a11_wr[1048];                
			assign x194_out     = a11_wr[536];                 
			assign x195_out     = a11_wr[1560];                
			assign x196_out     = a11_wr[280];                 
			assign x197_out     = a11_wr[1304];                
			assign x198_out     = a11_wr[792];                 
			assign x199_out     = a11_wr[1816];                
			assign x200_out     = a11_wr[152];                 
			assign x201_out     = a11_wr[1176];                
			assign x202_out     = a11_wr[664];                 
			assign x203_out     = a11_wr[1688];                
			assign x204_out     = a11_wr[408];                 
			assign x205_out     = a11_wr[1432];                
			assign x206_out     = a11_wr[920];                 
			assign x207_out     = a11_wr[1944];                
			assign x208_out     = a11_wr[88];                  
			assign x209_out     = a11_wr[1112];                
			assign x210_out     = a11_wr[600];                 
			assign x211_out     = a11_wr[1624];                
			assign x212_out     = a11_wr[344];                 
			assign x213_out     = a11_wr[1368];                
			assign x214_out     = a11_wr[856];                 
			assign x215_out     = a11_wr[1880];                
			assign x216_out     = a11_wr[216];                 
			assign x217_out     = a11_wr[1240];                
			assign x218_out     = a11_wr[728];                 
			assign x219_out     = a11_wr[1752];                
			assign x220_out     = a11_wr[472];                 
			assign x221_out     = a11_wr[1496];                
			assign x222_out     = a11_wr[984];                 
			assign x223_out     = a11_wr[2008];                
			assign x224_out     = a11_wr[56];                  
			assign x225_out     = a11_wr[1080];                
			assign x226_out     = a11_wr[568];                 
			assign x227_out     = a11_wr[1592];                
			assign x228_out     = a11_wr[312];                 
			assign x229_out     = a11_wr[1336];                
			assign x230_out     = a11_wr[824];                 
			assign x231_out     = a11_wr[1848];                
			assign x232_out     = a11_wr[184];                 
			assign x233_out     = a11_wr[1208];                
			assign x234_out     = a11_wr[696];                 
			assign x235_out     = a11_wr[1720];                
			assign x236_out     = a11_wr[440];                 
			assign x237_out     = a11_wr[1464];                
			assign x238_out     = a11_wr[952];                 
			assign x239_out     = a11_wr[1976];                
			assign x240_out     = a11_wr[120];                 
			assign x241_out     = a11_wr[1144];                
			assign x242_out     = a11_wr[632];                 
			assign x243_out     = a11_wr[1656];                
			assign x244_out     = a11_wr[376];                 
			assign x245_out     = a11_wr[1400];                
			assign x246_out     = a11_wr[888];                 
			assign x247_out     = a11_wr[1912];                
			assign x248_out     = a11_wr[248];                 
			assign x249_out     = a11_wr[1272];                
			assign x250_out     = a11_wr[760];                 
			assign x251_out     = a11_wr[1784];                
			assign x252_out     = a11_wr[504];                 
			assign x253_out     = a11_wr[1528];                
			assign x254_out     = a11_wr[1016];                
			assign x255_out     = a11_wr[2040];                
			assign x256_out     = a11_wr[4];                   
			assign x257_out     = a11_wr[1028];                
			assign x258_out     = a11_wr[516];                 
			assign x259_out     = a11_wr[1540];                
			assign x260_out     = a11_wr[260];                 
			assign x261_out     = a11_wr[1284];                
			assign x262_out     = a11_wr[772];                 
			assign x263_out     = a11_wr[1796];                
			assign x264_out     = a11_wr[132];                 
			assign x265_out     = a11_wr[1156];                
			assign x266_out     = a11_wr[644];                 
			assign x267_out     = a11_wr[1668];                
			assign x268_out     = a11_wr[388];                 
			assign x269_out     = a11_wr[1412];                
			assign x270_out     = a11_wr[900];                 
			assign x271_out     = a11_wr[1924];                
			assign x272_out     = a11_wr[68];                  
			assign x273_out     = a11_wr[1092];                
			assign x274_out     = a11_wr[580];                 
			assign x275_out     = a11_wr[1604];                
			assign x276_out     = a11_wr[324];                 
			assign x277_out     = a11_wr[1348];                
			assign x278_out     = a11_wr[836];                 
			assign x279_out     = a11_wr[1860];                
			assign x280_out     = a11_wr[196];                 
			assign x281_out     = a11_wr[1220];                
			assign x282_out     = a11_wr[708];                 
			assign x283_out     = a11_wr[1732];                
			assign x284_out     = a11_wr[452];                 
			assign x285_out     = a11_wr[1476];                
			assign x286_out     = a11_wr[964];                 
			assign x287_out     = a11_wr[1988];                
			assign x288_out     = a11_wr[36];                  
			assign x289_out     = a11_wr[1060];                
			assign x290_out     = a11_wr[548];                 
			assign x291_out     = a11_wr[1572];                
			assign x292_out     = a11_wr[292];                 
			assign x293_out     = a11_wr[1316];                
			assign x294_out     = a11_wr[804];                 
			assign x295_out     = a11_wr[1828];                
			assign x296_out     = a11_wr[164];                 
			assign x297_out     = a11_wr[1188];                
			assign x298_out     = a11_wr[676];                 
			assign x299_out     = a11_wr[1700];                
			assign x300_out     = a11_wr[420];                 
			assign x301_out     = a11_wr[1444];                
			assign x302_out     = a11_wr[932];                 
			assign x303_out     = a11_wr[1956];                
			assign x304_out     = a11_wr[100];                 
			assign x305_out     = a11_wr[1124];                
			assign x306_out     = a11_wr[612];                 
			assign x307_out     = a11_wr[1636];                
			assign x308_out     = a11_wr[356];                 
			assign x309_out     = a11_wr[1380];                
			assign x310_out     = a11_wr[868];                 
			assign x311_out     = a11_wr[1892];                
			assign x312_out     = a11_wr[228];                 
			assign x313_out     = a11_wr[1252];                
			assign x314_out     = a11_wr[740];                 
			assign x315_out     = a11_wr[1764];                
			assign x316_out     = a11_wr[484];                 
			assign x317_out     = a11_wr[1508];                
			assign x318_out     = a11_wr[996];                 
			assign x319_out     = a11_wr[2020];                
			assign x320_out     = a11_wr[20];                  
			assign x321_out     = a11_wr[1044];                
			assign x322_out     = a11_wr[532];                 
			assign x323_out     = a11_wr[1556];                
			assign x324_out     = a11_wr[276];                 
			assign x325_out     = a11_wr[1300];                
			assign x326_out     = a11_wr[788];                 
			assign x327_out     = a11_wr[1812];                
			assign x328_out     = a11_wr[148];                 
			assign x329_out     = a11_wr[1172];                
			assign x330_out     = a11_wr[660];                 
			assign x331_out     = a11_wr[1684];                
			assign x332_out     = a11_wr[404];                 
			assign x333_out     = a11_wr[1428];                
			assign x334_out     = a11_wr[916];                 
			assign x335_out     = a11_wr[1940];                
			assign x336_out     = a11_wr[84];                  
			assign x337_out     = a11_wr[1108];                
			assign x338_out     = a11_wr[596];                 
			assign x339_out     = a11_wr[1620];                
			assign x340_out     = a11_wr[340];                 
			assign x341_out     = a11_wr[1364];                
			assign x342_out     = a11_wr[852];                 
			assign x343_out     = a11_wr[1876];                
			assign x344_out     = a11_wr[212];                 
			assign x345_out     = a11_wr[1236];                
			assign x346_out     = a11_wr[724];                 
			assign x347_out     = a11_wr[1748];                
			assign x348_out     = a11_wr[468];                 
			assign x349_out     = a11_wr[1492];                
			assign x350_out     = a11_wr[980];                 
			assign x351_out     = a11_wr[2004];                
			assign x352_out     = a11_wr[52];                  
			assign x353_out     = a11_wr[1076];                
			assign x354_out     = a11_wr[564];                 
			assign x355_out     = a11_wr[1588];                
			assign x356_out     = a11_wr[308];                 
			assign x357_out     = a11_wr[1332];                
			assign x358_out     = a11_wr[820];                 
			assign x359_out     = a11_wr[1844];                
			assign x360_out     = a11_wr[180];                 
			assign x361_out     = a11_wr[1204];                
			assign x362_out     = a11_wr[692];                 
			assign x363_out     = a11_wr[1716];                
			assign x364_out     = a11_wr[436];                 
			assign x365_out     = a11_wr[1460];                
			assign x366_out     = a11_wr[948];                 
			assign x367_out     = a11_wr[1972];                
			assign x368_out     = a11_wr[116];                 
			assign x369_out     = a11_wr[1140];                
			assign x370_out     = a11_wr[628];                 
			assign x371_out     = a11_wr[1652];                
			assign x372_out     = a11_wr[372];                 
			assign x373_out     = a11_wr[1396];                
			assign x374_out     = a11_wr[884];                 
			assign x375_out     = a11_wr[1908];                
			assign x376_out     = a11_wr[244];                 
			assign x377_out     = a11_wr[1268];                
			assign x378_out     = a11_wr[756];                 
			assign x379_out     = a11_wr[1780];                
			assign x380_out     = a11_wr[500];                 
			assign x381_out     = a11_wr[1524];                
			assign x382_out     = a11_wr[1012];                
			assign x383_out     = a11_wr[2036];                
			assign x384_out     = a11_wr[12];                  
			assign x385_out     = a11_wr[1036];                
			assign x386_out     = a11_wr[524];                 
			assign x387_out     = a11_wr[1548];                
			assign x388_out     = a11_wr[268];                 
			assign x389_out     = a11_wr[1292];                
			assign x390_out     = a11_wr[780];                 
			assign x391_out     = a11_wr[1804];                
			assign x392_out     = a11_wr[140];                 
			assign x393_out     = a11_wr[1164];                
			assign x394_out     = a11_wr[652];                 
			assign x395_out     = a11_wr[1676];                
			assign x396_out     = a11_wr[396];                 
			assign x397_out     = a11_wr[1420];                
			assign x398_out     = a11_wr[908];                 
			assign x399_out     = a11_wr[1932];                
			assign x400_out     = a11_wr[76];                  
			assign x401_out     = a11_wr[1100];                
			assign x402_out     = a11_wr[588];                 
			assign x403_out     = a11_wr[1612];                
			assign x404_out     = a11_wr[332];                 
			assign x405_out     = a11_wr[1356];                
			assign x406_out     = a11_wr[844];                 
			assign x407_out     = a11_wr[1868];                
			assign x408_out     = a11_wr[204];                 
			assign x409_out     = a11_wr[1228];                
			assign x410_out     = a11_wr[716];                 
			assign x411_out     = a11_wr[1740];                
			assign x412_out     = a11_wr[460];                 
			assign x413_out     = a11_wr[1484];                
			assign x414_out     = a11_wr[972];                 
			assign x415_out     = a11_wr[1996];                
			assign x416_out     = a11_wr[44];                  
			assign x417_out     = a11_wr[1068];                
			assign x418_out     = a11_wr[556];                 
			assign x419_out     = a11_wr[1580];                
			assign x420_out     = a11_wr[300];                 
			assign x421_out     = a11_wr[1324];                
			assign x422_out     = a11_wr[812];                 
			assign x423_out     = a11_wr[1836];                
			assign x424_out     = a11_wr[172];                 
			assign x425_out     = a11_wr[1196];                
			assign x426_out     = a11_wr[684];                 
			assign x427_out     = a11_wr[1708];                
			assign x428_out     = a11_wr[428];                 
			assign x429_out     = a11_wr[1452];                
			assign x430_out     = a11_wr[940];                 
			assign x431_out     = a11_wr[1964];                
			assign x432_out     = a11_wr[108];                 
			assign x433_out     = a11_wr[1132];                
			assign x434_out     = a11_wr[620];                 
			assign x435_out     = a11_wr[1644];                
			assign x436_out     = a11_wr[364];                 
			assign x437_out     = a11_wr[1388];                
			assign x438_out     = a11_wr[876];                 
			assign x439_out     = a11_wr[1900];                
			assign x440_out     = a11_wr[236];                 
			assign x441_out     = a11_wr[1260];                
			assign x442_out     = a11_wr[748];                 
			assign x443_out     = a11_wr[1772];                
			assign x444_out     = a11_wr[492];                 
			assign x445_out     = a11_wr[1516];                
			assign x446_out     = a11_wr[1004];                
			assign x447_out     = a11_wr[2028];                
			assign x448_out     = a11_wr[28];                  
			assign x449_out     = a11_wr[1052];                
			assign x450_out     = a11_wr[540];                 
			assign x451_out     = a11_wr[1564];                
			assign x452_out     = a11_wr[284];                 
			assign x453_out     = a11_wr[1308];                
			assign x454_out     = a11_wr[796];                 
			assign x455_out     = a11_wr[1820];                
			assign x456_out     = a11_wr[156];                 
			assign x457_out     = a11_wr[1180];                
			assign x458_out     = a11_wr[668];                 
			assign x459_out     = a11_wr[1692];                
			assign x460_out     = a11_wr[412];                 
			assign x461_out     = a11_wr[1436];                
			assign x462_out     = a11_wr[924];                 
			assign x463_out     = a11_wr[1948];                
			assign x464_out     = a11_wr[92];                  
			assign x465_out     = a11_wr[1116];                
			assign x466_out     = a11_wr[604];                 
			assign x467_out     = a11_wr[1628];                
			assign x468_out     = a11_wr[348];                 
			assign x469_out     = a11_wr[1372];                
			assign x470_out     = a11_wr[860];                 
			assign x471_out     = a11_wr[1884];                
			assign x472_out     = a11_wr[220];                 
			assign x473_out     = a11_wr[1244];                
			assign x474_out     = a11_wr[732];                 
			assign x475_out     = a11_wr[1756];                
			assign x476_out     = a11_wr[476];                 
			assign x477_out     = a11_wr[1500];                
			assign x478_out     = a11_wr[988];                 
			assign x479_out     = a11_wr[2012];                
			assign x480_out     = a11_wr[60];                  
			assign x481_out     = a11_wr[1084];                
			assign x482_out     = a11_wr[572];                 
			assign x483_out     = a11_wr[1596];                
			assign x484_out     = a11_wr[316];                 
			assign x485_out     = a11_wr[1340];                
			assign x486_out     = a11_wr[828];                 
			assign x487_out     = a11_wr[1852];                
			assign x488_out     = a11_wr[188];                 
			assign x489_out     = a11_wr[1212];                
			assign x490_out     = a11_wr[700];                 
			assign x491_out     = a11_wr[1724];                
			assign x492_out     = a11_wr[444];                 
			assign x493_out     = a11_wr[1468];                
			assign x494_out     = a11_wr[956];                 
			assign x495_out     = a11_wr[1980];                
			assign x496_out     = a11_wr[124];                 
			assign x497_out     = a11_wr[1148];                
			assign x498_out     = a11_wr[636];                 
			assign x499_out     = a11_wr[1660];                
			assign x500_out     = a11_wr[380];                 
			assign x501_out     = a11_wr[1404];                
			assign x502_out     = a11_wr[892];                 
			assign x503_out     = a11_wr[1916];                
			assign x504_out     = a11_wr[252];                 
			assign x505_out     = a11_wr[1276];                
			assign x506_out     = a11_wr[764];                 
			assign x507_out     = a11_wr[1788];                
			assign x508_out     = a11_wr[508];                 
			assign x509_out     = a11_wr[1532];                
			assign x510_out     = a11_wr[1020];                
			assign x511_out     = a11_wr[2044];                
			assign x512_out     = a11_wr[2];                   
			assign x513_out     = a11_wr[1026];                
			assign x514_out     = a11_wr[514];                 
			assign x515_out     = a11_wr[1538];                
			assign x516_out     = a11_wr[258];                 
			assign x517_out     = a11_wr[1282];                
			assign x518_out     = a11_wr[770];                 
			assign x519_out     = a11_wr[1794];                
			assign x520_out     = a11_wr[130];                 
			assign x521_out     = a11_wr[1154];                
			assign x522_out     = a11_wr[642];                 
			assign x523_out     = a11_wr[1666];                
			assign x524_out     = a11_wr[386];                 
			assign x525_out     = a11_wr[1410];                
			assign x526_out     = a11_wr[898];                 
			assign x527_out     = a11_wr[1922];                
			assign x528_out     = a11_wr[66];                  
			assign x529_out     = a11_wr[1090];                
			assign x530_out     = a11_wr[578];                 
			assign x531_out     = a11_wr[1602];                
			assign x532_out     = a11_wr[322];                 
			assign x533_out     = a11_wr[1346];                
			assign x534_out     = a11_wr[834];                 
			assign x535_out     = a11_wr[1858];                
			assign x536_out     = a11_wr[194];                 
			assign x537_out     = a11_wr[1218];                
			assign x538_out     = a11_wr[706];                 
			assign x539_out     = a11_wr[1730];                
			assign x540_out     = a11_wr[450];                 
			assign x541_out     = a11_wr[1474];                
			assign x542_out     = a11_wr[962];                 
			assign x543_out     = a11_wr[1986];                
			assign x544_out     = a11_wr[34];                  
			assign x545_out     = a11_wr[1058];                
			assign x546_out     = a11_wr[546];                 
			assign x547_out     = a11_wr[1570];                
			assign x548_out     = a11_wr[290];                 
			assign x549_out     = a11_wr[1314];                
			assign x550_out     = a11_wr[802];                 
			assign x551_out     = a11_wr[1826];                
			assign x552_out     = a11_wr[162];                 
			assign x553_out     = a11_wr[1186];                
			assign x554_out     = a11_wr[674];                 
			assign x555_out     = a11_wr[1698];                
			assign x556_out     = a11_wr[418];                 
			assign x557_out     = a11_wr[1442];                
			assign x558_out     = a11_wr[930];                 
			assign x559_out     = a11_wr[1954];                
			assign x560_out     = a11_wr[98];                  
			assign x561_out     = a11_wr[1122];                
			assign x562_out     = a11_wr[610];                 
			assign x563_out     = a11_wr[1634];                
			assign x564_out     = a11_wr[354];                 
			assign x565_out     = a11_wr[1378];                
			assign x566_out     = a11_wr[866];                 
			assign x567_out     = a11_wr[1890];                
			assign x568_out     = a11_wr[226];                 
			assign x569_out     = a11_wr[1250];                
			assign x570_out     = a11_wr[738];                 
			assign x571_out     = a11_wr[1762];                
			assign x572_out     = a11_wr[482];                 
			assign x573_out     = a11_wr[1506];                
			assign x574_out     = a11_wr[994];                 
			assign x575_out     = a11_wr[2018];                
			assign x576_out     = a11_wr[18];                  
			assign x577_out     = a11_wr[1042];                
			assign x578_out     = a11_wr[530];                 
			assign x579_out     = a11_wr[1554];                
			assign x580_out     = a11_wr[274];                 
			assign x581_out     = a11_wr[1298];                
			assign x582_out     = a11_wr[786];                 
			assign x583_out     = a11_wr[1810];                
			assign x584_out     = a11_wr[146];                 
			assign x585_out     = a11_wr[1170];                
			assign x586_out     = a11_wr[658];                 
			assign x587_out     = a11_wr[1682];                
			assign x588_out     = a11_wr[402];                 
			assign x589_out     = a11_wr[1426];                
			assign x590_out     = a11_wr[914];                 
			assign x591_out     = a11_wr[1938];                
			assign x592_out     = a11_wr[82];                  
			assign x593_out     = a11_wr[1106];                
			assign x594_out     = a11_wr[594];                 
			assign x595_out     = a11_wr[1618];                
			assign x596_out     = a11_wr[338];                 
			assign x597_out     = a11_wr[1362];                
			assign x598_out     = a11_wr[850];                 
			assign x599_out     = a11_wr[1874];                
			assign x600_out     = a11_wr[210];                 
			assign x601_out     = a11_wr[1234];                
			assign x602_out     = a11_wr[722];                 
			assign x603_out     = a11_wr[1746];                
			assign x604_out     = a11_wr[466];                 
			assign x605_out     = a11_wr[1490];                
			assign x606_out     = a11_wr[978];                 
			assign x607_out     = a11_wr[2002];                
			assign x608_out     = a11_wr[50];                  
			assign x609_out     = a11_wr[1074];                
			assign x610_out     = a11_wr[562];                 
			assign x611_out     = a11_wr[1586];                
			assign x612_out     = a11_wr[306];                 
			assign x613_out     = a11_wr[1330];                
			assign x614_out     = a11_wr[818];                 
			assign x615_out     = a11_wr[1842];                
			assign x616_out     = a11_wr[178];                 
			assign x617_out     = a11_wr[1202];                
			assign x618_out     = a11_wr[690];                 
			assign x619_out     = a11_wr[1714];                
			assign x620_out     = a11_wr[434];                 
			assign x621_out     = a11_wr[1458];                
			assign x622_out     = a11_wr[946];                 
			assign x623_out     = a11_wr[1970];                
			assign x624_out     = a11_wr[114];                 
			assign x625_out     = a11_wr[1138];                
			assign x626_out     = a11_wr[626];                 
			assign x627_out     = a11_wr[1650];                
			assign x628_out     = a11_wr[370];                 
			assign x629_out     = a11_wr[1394];                
			assign x630_out     = a11_wr[882];                 
			assign x631_out     = a11_wr[1906];                
			assign x632_out     = a11_wr[242];                 
			assign x633_out     = a11_wr[1266];                
			assign x634_out     = a11_wr[754];                 
			assign x635_out     = a11_wr[1778];                
			assign x636_out     = a11_wr[498];                 
			assign x637_out     = a11_wr[1522];                
			assign x638_out     = a11_wr[1010];                
			assign x639_out     = a11_wr[2034];                
			assign x640_out     = a11_wr[10];                  
			assign x641_out     = a11_wr[1034];                
			assign x642_out     = a11_wr[522];                 
			assign x643_out     = a11_wr[1546];                
			assign x644_out     = a11_wr[266];                 
			assign x645_out     = a11_wr[1290];                
			assign x646_out     = a11_wr[778];                 
			assign x647_out     = a11_wr[1802];                
			assign x648_out     = a11_wr[138];                 
			assign x649_out     = a11_wr[1162];                
			assign x650_out     = a11_wr[650];                 
			assign x651_out     = a11_wr[1674];                
			assign x652_out     = a11_wr[394];                 
			assign x653_out     = a11_wr[1418];                
			assign x654_out     = a11_wr[906];                 
			assign x655_out     = a11_wr[1930];                
			assign x656_out     = a11_wr[74];                  
			assign x657_out     = a11_wr[1098];                
			assign x658_out     = a11_wr[586];                 
			assign x659_out     = a11_wr[1610];                
			assign x660_out     = a11_wr[330];                 
			assign x661_out     = a11_wr[1354];                
			assign x662_out     = a11_wr[842];                 
			assign x663_out     = a11_wr[1866];                
			assign x664_out     = a11_wr[202];                 
			assign x665_out     = a11_wr[1226];                
			assign x666_out     = a11_wr[714];                 
			assign x667_out     = a11_wr[1738];                
			assign x668_out     = a11_wr[458];                 
			assign x669_out     = a11_wr[1482];                
			assign x670_out     = a11_wr[970];                 
			assign x671_out     = a11_wr[1994];                
			assign x672_out     = a11_wr[42];                  
			assign x673_out     = a11_wr[1066];                
			assign x674_out     = a11_wr[554];                 
			assign x675_out     = a11_wr[1578];                
			assign x676_out     = a11_wr[298];                 
			assign x677_out     = a11_wr[1322];                
			assign x678_out     = a11_wr[810];                 
			assign x679_out     = a11_wr[1834];                
			assign x680_out     = a11_wr[170];                 
			assign x681_out     = a11_wr[1194];                
			assign x682_out     = a11_wr[682];                 
			assign x683_out     = a11_wr[1706];                
			assign x684_out     = a11_wr[426];                 
			assign x685_out     = a11_wr[1450];                
			assign x686_out     = a11_wr[938];                 
			assign x687_out     = a11_wr[1962];                
			assign x688_out     = a11_wr[106];                 
			assign x689_out     = a11_wr[1130];                
			assign x690_out     = a11_wr[618];                 
			assign x691_out     = a11_wr[1642];                
			assign x692_out     = a11_wr[362];                 
			assign x693_out     = a11_wr[1386];                
			assign x694_out     = a11_wr[874];                 
			assign x695_out     = a11_wr[1898];                
			assign x696_out     = a11_wr[234];                 
			assign x697_out     = a11_wr[1258];                
			assign x698_out     = a11_wr[746];                 
			assign x699_out     = a11_wr[1770];                
			assign x700_out     = a11_wr[490];                 
			assign x701_out     = a11_wr[1514];                
			assign x702_out     = a11_wr[1002];                
			assign x703_out     = a11_wr[2026];                
			assign x704_out     = a11_wr[26];                  
			assign x705_out     = a11_wr[1050];                
			assign x706_out     = a11_wr[538];                 
			assign x707_out     = a11_wr[1562];                
			assign x708_out     = a11_wr[282];                 
			assign x709_out     = a11_wr[1306];                
			assign x710_out     = a11_wr[794];                 
			assign x711_out     = a11_wr[1818];                
			assign x712_out     = a11_wr[154];                 
			assign x713_out     = a11_wr[1178];                
			assign x714_out     = a11_wr[666];                 
			assign x715_out     = a11_wr[1690];                
			assign x716_out     = a11_wr[410];                 
			assign x717_out     = a11_wr[1434];                
			assign x718_out     = a11_wr[922];                 
			assign x719_out     = a11_wr[1946];                
			assign x720_out     = a11_wr[90];                  
			assign x721_out     = a11_wr[1114];                
			assign x722_out     = a11_wr[602];                 
			assign x723_out     = a11_wr[1626];                
			assign x724_out     = a11_wr[346];                 
			assign x725_out     = a11_wr[1370];                
			assign x726_out     = a11_wr[858];                 
			assign x727_out     = a11_wr[1882];                
			assign x728_out     = a11_wr[218];                 
			assign x729_out     = a11_wr[1242];                
			assign x730_out     = a11_wr[730];                 
			assign x731_out     = a11_wr[1754];                
			assign x732_out     = a11_wr[474];                 
			assign x733_out     = a11_wr[1498];                
			assign x734_out     = a11_wr[986];                 
			assign x735_out     = a11_wr[2010];                
			assign x736_out     = a11_wr[58];                  
			assign x737_out     = a11_wr[1082];                
			assign x738_out     = a11_wr[570];                 
			assign x739_out     = a11_wr[1594];                
			assign x740_out     = a11_wr[314];                 
			assign x741_out     = a11_wr[1338];                
			assign x742_out     = a11_wr[826];                 
			assign x743_out     = a11_wr[1850];                
			assign x744_out     = a11_wr[186];                 
			assign x745_out     = a11_wr[1210];                
			assign x746_out     = a11_wr[698];                 
			assign x747_out     = a11_wr[1722];                
			assign x748_out     = a11_wr[442];                 
			assign x749_out     = a11_wr[1466];                
			assign x750_out     = a11_wr[954];                 
			assign x751_out     = a11_wr[1978];                
			assign x752_out     = a11_wr[122];                 
			assign x753_out     = a11_wr[1146];                
			assign x754_out     = a11_wr[634];                 
			assign x755_out     = a11_wr[1658];                
			assign x756_out     = a11_wr[378];                 
			assign x757_out     = a11_wr[1402];                
			assign x758_out     = a11_wr[890];                 
			assign x759_out     = a11_wr[1914];                
			assign x760_out     = a11_wr[250];                 
			assign x761_out     = a11_wr[1274];                
			assign x762_out     = a11_wr[762];                 
			assign x763_out     = a11_wr[1786];                
			assign x764_out     = a11_wr[506];                 
			assign x765_out     = a11_wr[1530];                
			assign x766_out     = a11_wr[1018];                
			assign x767_out     = a11_wr[2042];                
			assign x768_out     = a11_wr[6];                   
			assign x769_out     = a11_wr[1030];                
			assign x770_out     = a11_wr[518];                 
			assign x771_out     = a11_wr[1542];                
			assign x772_out     = a11_wr[262];                 
			assign x773_out     = a11_wr[1286];                
			assign x774_out     = a11_wr[774];                 
			assign x775_out     = a11_wr[1798];                
			assign x776_out     = a11_wr[134];                 
			assign x777_out     = a11_wr[1158];                
			assign x778_out     = a11_wr[646];                 
			assign x779_out     = a11_wr[1670];                
			assign x780_out     = a11_wr[390];                 
			assign x781_out     = a11_wr[1414];                
			assign x782_out     = a11_wr[902];                 
			assign x783_out     = a11_wr[1926];                
			assign x784_out     = a11_wr[70];                  
			assign x785_out     = a11_wr[1094];                
			assign x786_out     = a11_wr[582];                 
			assign x787_out     = a11_wr[1606];                
			assign x788_out     = a11_wr[326];                 
			assign x789_out     = a11_wr[1350];                
			assign x790_out     = a11_wr[838];                 
			assign x791_out     = a11_wr[1862];                
			assign x792_out     = a11_wr[198];                 
			assign x793_out     = a11_wr[1222];                
			assign x794_out     = a11_wr[710];                 
			assign x795_out     = a11_wr[1734];                
			assign x796_out     = a11_wr[454];                 
			assign x797_out     = a11_wr[1478];                
			assign x798_out     = a11_wr[966];                 
			assign x799_out     = a11_wr[1990];                
			assign x800_out     = a11_wr[38];                  
			assign x801_out     = a11_wr[1062];                
			assign x802_out     = a11_wr[550];                 
			assign x803_out     = a11_wr[1574];                
			assign x804_out     = a11_wr[294];                 
			assign x805_out     = a11_wr[1318];                
			assign x806_out     = a11_wr[806];                 
			assign x807_out     = a11_wr[1830];                
			assign x808_out     = a11_wr[166];                 
			assign x809_out     = a11_wr[1190];                
			assign x810_out     = a11_wr[678];                 
			assign x811_out     = a11_wr[1702];                
			assign x812_out     = a11_wr[422];                 
			assign x813_out     = a11_wr[1446];                
			assign x814_out     = a11_wr[934];                 
			assign x815_out     = a11_wr[1958];                
			assign x816_out     = a11_wr[102];                 
			assign x817_out     = a11_wr[1126];                
			assign x818_out     = a11_wr[614];                 
			assign x819_out     = a11_wr[1638];                
			assign x820_out     = a11_wr[358];                 
			assign x821_out     = a11_wr[1382];                
			assign x822_out     = a11_wr[870];                 
			assign x823_out     = a11_wr[1894];                
			assign x824_out     = a11_wr[230];                 
			assign x825_out     = a11_wr[1254];                
			assign x826_out     = a11_wr[742];                 
			assign x827_out     = a11_wr[1766];                
			assign x828_out     = a11_wr[486];                 
			assign x829_out     = a11_wr[1510];                
			assign x830_out     = a11_wr[998];                 
			assign x831_out     = a11_wr[2022];                
			assign x832_out     = a11_wr[22];                  
			assign x833_out     = a11_wr[1046];                
			assign x834_out     = a11_wr[534];                 
			assign x835_out     = a11_wr[1558];                
			assign x836_out     = a11_wr[278];                 
			assign x837_out     = a11_wr[1302];                
			assign x838_out     = a11_wr[790];                 
			assign x839_out     = a11_wr[1814];                
			assign x840_out     = a11_wr[150];                 
			assign x841_out     = a11_wr[1174];                
			assign x842_out     = a11_wr[662];                 
			assign x843_out     = a11_wr[1686];                
			assign x844_out     = a11_wr[406];                 
			assign x845_out     = a11_wr[1430];                
			assign x846_out     = a11_wr[918];                 
			assign x847_out     = a11_wr[1942];                
			assign x848_out     = a11_wr[86];                  
			assign x849_out     = a11_wr[1110];                
			assign x850_out     = a11_wr[598];                 
			assign x851_out     = a11_wr[1622];                
			assign x852_out     = a11_wr[342];                 
			assign x853_out     = a11_wr[1366];                
			assign x854_out     = a11_wr[854];                 
			assign x855_out     = a11_wr[1878];                
			assign x856_out     = a11_wr[214];                 
			assign x857_out     = a11_wr[1238];                
			assign x858_out     = a11_wr[726];                 
			assign x859_out     = a11_wr[1750];                
			assign x860_out     = a11_wr[470];                 
			assign x861_out     = a11_wr[1494];                
			assign x862_out     = a11_wr[982];                 
			assign x863_out     = a11_wr[2006];                
			assign x864_out     = a11_wr[54];                  
			assign x865_out     = a11_wr[1078];                
			assign x866_out     = a11_wr[566];                 
			assign x867_out     = a11_wr[1590];                
			assign x868_out     = a11_wr[310];                 
			assign x869_out     = a11_wr[1334];                
			assign x870_out     = a11_wr[822];                 
			assign x871_out     = a11_wr[1846];                
			assign x872_out     = a11_wr[182];                 
			assign x873_out     = a11_wr[1206];                
			assign x874_out     = a11_wr[694];                 
			assign x875_out     = a11_wr[1718];                
			assign x876_out     = a11_wr[438];                 
			assign x877_out     = a11_wr[1462];                
			assign x878_out     = a11_wr[950];                 
			assign x879_out     = a11_wr[1974];                
			assign x880_out     = a11_wr[118];                 
			assign x881_out     = a11_wr[1142];                
			assign x882_out     = a11_wr[630];                 
			assign x883_out     = a11_wr[1654];                
			assign x884_out     = a11_wr[374];                 
			assign x885_out     = a11_wr[1398];                
			assign x886_out     = a11_wr[886];                 
			assign x887_out     = a11_wr[1910];                
			assign x888_out     = a11_wr[246];                 
			assign x889_out     = a11_wr[1270];                
			assign x890_out     = a11_wr[758];                 
			assign x891_out     = a11_wr[1782];                
			assign x892_out     = a11_wr[502];                 
			assign x893_out     = a11_wr[1526];                
			assign x894_out     = a11_wr[1014];                
			assign x895_out     = a11_wr[2038];                
			assign x896_out     = a11_wr[14];                  
			assign x897_out     = a11_wr[1038];                
			assign x898_out     = a11_wr[526];                 
			assign x899_out     = a11_wr[1550];                
			assign x900_out     = a11_wr[270];                 
			assign x901_out     = a11_wr[1294];                
			assign x902_out     = a11_wr[782];                 
			assign x903_out     = a11_wr[1806];                
			assign x904_out     = a11_wr[142];                 
			assign x905_out     = a11_wr[1166];                
			assign x906_out     = a11_wr[654];                 
			assign x907_out     = a11_wr[1678];                
			assign x908_out     = a11_wr[398];                 
			assign x909_out     = a11_wr[1422];                
			assign x910_out     = a11_wr[910];                 
			assign x911_out     = a11_wr[1934];                
			assign x912_out     = a11_wr[78];                  
			assign x913_out     = a11_wr[1102];                
			assign x914_out     = a11_wr[590];                 
			assign x915_out     = a11_wr[1614];                
			assign x916_out     = a11_wr[334];                 
			assign x917_out     = a11_wr[1358];                
			assign x918_out     = a11_wr[846];                 
			assign x919_out     = a11_wr[1870];                
			assign x920_out     = a11_wr[206];                 
			assign x921_out     = a11_wr[1230];                
			assign x922_out     = a11_wr[718];                 
			assign x923_out     = a11_wr[1742];                
			assign x924_out     = a11_wr[462];                 
			assign x925_out     = a11_wr[1486];                
			assign x926_out     = a11_wr[974];                 
			assign x927_out     = a11_wr[1998];                
			assign x928_out     = a11_wr[46];                  
			assign x929_out     = a11_wr[1070];                
			assign x930_out     = a11_wr[558];                 
			assign x931_out     = a11_wr[1582];                
			assign x932_out     = a11_wr[302];                 
			assign x933_out     = a11_wr[1326];                
			assign x934_out     = a11_wr[814];                 
			assign x935_out     = a11_wr[1838];                
			assign x936_out     = a11_wr[174];                 
			assign x937_out     = a11_wr[1198];                
			assign x938_out     = a11_wr[686];                 
			assign x939_out     = a11_wr[1710];                
			assign x940_out     = a11_wr[430];                 
			assign x941_out     = a11_wr[1454];                
			assign x942_out     = a11_wr[942];                 
			assign x943_out     = a11_wr[1966];                
			assign x944_out     = a11_wr[110];                 
			assign x945_out     = a11_wr[1134];                
			assign x946_out     = a11_wr[622];                 
			assign x947_out     = a11_wr[1646];                
			assign x948_out     = a11_wr[366];                 
			assign x949_out     = a11_wr[1390];                
			assign x950_out     = a11_wr[878];                 
			assign x951_out     = a11_wr[1902];                
			assign x952_out     = a11_wr[238];                 
			assign x953_out     = a11_wr[1262];                
			assign x954_out     = a11_wr[750];                 
			assign x955_out     = a11_wr[1774];                
			assign x956_out     = a11_wr[494];                 
			assign x957_out     = a11_wr[1518];                
			assign x958_out     = a11_wr[1006];                
			assign x959_out     = a11_wr[2030];                
			assign x960_out     = a11_wr[30];                  
			assign x961_out     = a11_wr[1054];                
			assign x962_out     = a11_wr[542];                 
			assign x963_out     = a11_wr[1566];                
			assign x964_out     = a11_wr[286];                 
			assign x965_out     = a11_wr[1310];                
			assign x966_out     = a11_wr[798];                 
			assign x967_out     = a11_wr[1822];                
			assign x968_out     = a11_wr[158];                 
			assign x969_out     = a11_wr[1182];                
			assign x970_out     = a11_wr[670];                 
			assign x971_out     = a11_wr[1694];                
			assign x972_out     = a11_wr[414];                 
			assign x973_out     = a11_wr[1438];                
			assign x974_out     = a11_wr[926];                 
			assign x975_out     = a11_wr[1950];                
			assign x976_out     = a11_wr[94];                  
			assign x977_out     = a11_wr[1118];                
			assign x978_out     = a11_wr[606];                 
			assign x979_out     = a11_wr[1630];                
			assign x980_out     = a11_wr[350];                 
			assign x981_out     = a11_wr[1374];                
			assign x982_out     = a11_wr[862];                 
			assign x983_out     = a11_wr[1886];                
			assign x984_out     = a11_wr[222];                 
			assign x985_out     = a11_wr[1246];                
			assign x986_out     = a11_wr[734];                 
			assign x987_out     = a11_wr[1758];                
			assign x988_out     = a11_wr[478];                 
			assign x989_out     = a11_wr[1502];                
			assign x990_out     = a11_wr[990];                 
			assign x991_out     = a11_wr[2014];                
			assign x992_out     = a11_wr[62];                  
			assign x993_out     = a11_wr[1086];                
			assign x994_out     = a11_wr[574];                 
			assign x995_out     = a11_wr[1598];                
			assign x996_out     = a11_wr[318];                 
			assign x997_out     = a11_wr[1342];                
			assign x998_out     = a11_wr[830];                 
			assign x999_out     = a11_wr[1854];                
			assign x1000_out    = a11_wr[190];                 
			assign x1001_out    = a11_wr[1214];                
			assign x1002_out    = a11_wr[702];                 
			assign x1003_out    = a11_wr[1726];                
			assign x1004_out    = a11_wr[446];                 
			assign x1005_out    = a11_wr[1470];                
			assign x1006_out    = a11_wr[958];                 
			assign x1007_out    = a11_wr[1982];                
			assign x1008_out    = a11_wr[126];                 
			assign x1009_out    = a11_wr[1150];                
			assign x1010_out    = a11_wr[638];                 
			assign x1011_out    = a11_wr[1662];                
			assign x1012_out    = a11_wr[382];                 
			assign x1013_out    = a11_wr[1406];                
			assign x1014_out    = a11_wr[894];                 
			assign x1015_out    = a11_wr[1918];                
			assign x1016_out    = a11_wr[254];                 
			assign x1017_out    = a11_wr[1278];                
			assign x1018_out    = a11_wr[766];                 
			assign x1019_out    = a11_wr[1790];                
			assign x1020_out    = a11_wr[510];                 
			assign x1021_out    = a11_wr[1534];                
			assign x1022_out    = a11_wr[1022];                
			assign x1023_out    = a11_wr[2046];                
			assign x1024_out    = a11_wr[1];                   
			assign x1025_out    = a11_wr[1025];                
			assign x1026_out    = a11_wr[513];                 
			assign x1027_out    = a11_wr[1537];                
			assign x1028_out    = a11_wr[257];                 
			assign x1029_out    = a11_wr[1281];                
			assign x1030_out    = a11_wr[769];                 
			assign x1031_out    = a11_wr[1793];                
			assign x1032_out    = a11_wr[129];                 
			assign x1033_out    = a11_wr[1153];                
			assign x1034_out    = a11_wr[641];                 
			assign x1035_out    = a11_wr[1665];                
			assign x1036_out    = a11_wr[385];                 
			assign x1037_out    = a11_wr[1409];                
			assign x1038_out    = a11_wr[897];                 
			assign x1039_out    = a11_wr[1921];                
			assign x1040_out    = a11_wr[65];                  
			assign x1041_out    = a11_wr[1089];                
			assign x1042_out    = a11_wr[577];                 
			assign x1043_out    = a11_wr[1601];                
			assign x1044_out    = a11_wr[321];                 
			assign x1045_out    = a11_wr[1345];                
			assign x1046_out    = a11_wr[833];                 
			assign x1047_out    = a11_wr[1857];                
			assign x1048_out    = a11_wr[193];                 
			assign x1049_out    = a11_wr[1217];                
			assign x1050_out    = a11_wr[705];                 
			assign x1051_out    = a11_wr[1729];                
			assign x1052_out    = a11_wr[449];                 
			assign x1053_out    = a11_wr[1473];                
			assign x1054_out    = a11_wr[961];                 
			assign x1055_out    = a11_wr[1985];                
			assign x1056_out    = a11_wr[33];                  
			assign x1057_out    = a11_wr[1057];                
			assign x1058_out    = a11_wr[545];                 
			assign x1059_out    = a11_wr[1569];                
			assign x1060_out    = a11_wr[289];                 
			assign x1061_out    = a11_wr[1313];                
			assign x1062_out    = a11_wr[801];                 
			assign x1063_out    = a11_wr[1825];                
			assign x1064_out    = a11_wr[161];                 
			assign x1065_out    = a11_wr[1185];                
			assign x1066_out    = a11_wr[673];                 
			assign x1067_out    = a11_wr[1697];                
			assign x1068_out    = a11_wr[417];                 
			assign x1069_out    = a11_wr[1441];                
			assign x1070_out    = a11_wr[929];                 
			assign x1071_out    = a11_wr[1953];                
			assign x1072_out    = a11_wr[97];                  
			assign x1073_out    = a11_wr[1121];                
			assign x1074_out    = a11_wr[609];                 
			assign x1075_out    = a11_wr[1633];                
			assign x1076_out    = a11_wr[353];                 
			assign x1077_out    = a11_wr[1377];                
			assign x1078_out    = a11_wr[865];                 
			assign x1079_out    = a11_wr[1889];                
			assign x1080_out    = a11_wr[225];                 
			assign x1081_out    = a11_wr[1249];                
			assign x1082_out    = a11_wr[737];                 
			assign x1083_out    = a11_wr[1761];                
			assign x1084_out    = a11_wr[481];                 
			assign x1085_out    = a11_wr[1505];                
			assign x1086_out    = a11_wr[993];                 
			assign x1087_out    = a11_wr[2017];                
			assign x1088_out    = a11_wr[17];                  
			assign x1089_out    = a11_wr[1041];                
			assign x1090_out    = a11_wr[529];                 
			assign x1091_out    = a11_wr[1553];                
			assign x1092_out    = a11_wr[273];                 
			assign x1093_out    = a11_wr[1297];                
			assign x1094_out    = a11_wr[785];                 
			assign x1095_out    = a11_wr[1809];                
			assign x1096_out    = a11_wr[145];                 
			assign x1097_out    = a11_wr[1169];                
			assign x1098_out    = a11_wr[657];                 
			assign x1099_out    = a11_wr[1681];                
			assign x1100_out    = a11_wr[401];                 
			assign x1101_out    = a11_wr[1425];                
			assign x1102_out    = a11_wr[913];                 
			assign x1103_out    = a11_wr[1937];                
			assign x1104_out    = a11_wr[81];                  
			assign x1105_out    = a11_wr[1105];                
			assign x1106_out    = a11_wr[593];                 
			assign x1107_out    = a11_wr[1617];                
			assign x1108_out    = a11_wr[337];                 
			assign x1109_out    = a11_wr[1361];                
			assign x1110_out    = a11_wr[849];                 
			assign x1111_out    = a11_wr[1873];                
			assign x1112_out    = a11_wr[209];                 
			assign x1113_out    = a11_wr[1233];                
			assign x1114_out    = a11_wr[721];                 
			assign x1115_out    = a11_wr[1745];                
			assign x1116_out    = a11_wr[465];                 
			assign x1117_out    = a11_wr[1489];                
			assign x1118_out    = a11_wr[977];                 
			assign x1119_out    = a11_wr[2001];                
			assign x1120_out    = a11_wr[49];                  
			assign x1121_out    = a11_wr[1073];                
			assign x1122_out    = a11_wr[561];                 
			assign x1123_out    = a11_wr[1585];                
			assign x1124_out    = a11_wr[305];                 
			assign x1125_out    = a11_wr[1329];                
			assign x1126_out    = a11_wr[817];                 
			assign x1127_out    = a11_wr[1841];                
			assign x1128_out    = a11_wr[177];                 
			assign x1129_out    = a11_wr[1201];                
			assign x1130_out    = a11_wr[689];                 
			assign x1131_out    = a11_wr[1713];                
			assign x1132_out    = a11_wr[433];                 
			assign x1133_out    = a11_wr[1457];                
			assign x1134_out    = a11_wr[945];                 
			assign x1135_out    = a11_wr[1969];                
			assign x1136_out    = a11_wr[113];                 
			assign x1137_out    = a11_wr[1137];                
			assign x1138_out    = a11_wr[625];                 
			assign x1139_out    = a11_wr[1649];                
			assign x1140_out    = a11_wr[369];                 
			assign x1141_out    = a11_wr[1393];                
			assign x1142_out    = a11_wr[881];                 
			assign x1143_out    = a11_wr[1905];                
			assign x1144_out    = a11_wr[241];                 
			assign x1145_out    = a11_wr[1265];                
			assign x1146_out    = a11_wr[753];                 
			assign x1147_out    = a11_wr[1777];                
			assign x1148_out    = a11_wr[497];                 
			assign x1149_out    = a11_wr[1521];                
			assign x1150_out    = a11_wr[1009];                
			assign x1151_out    = a11_wr[2033];                
			assign x1152_out    = a11_wr[9];                   
			assign x1153_out    = a11_wr[1033];                
			assign x1154_out    = a11_wr[521];                 
			assign x1155_out    = a11_wr[1545];                
			assign x1156_out    = a11_wr[265];                 
			assign x1157_out    = a11_wr[1289];                
			assign x1158_out    = a11_wr[777];                 
			assign x1159_out    = a11_wr[1801];                
			assign x1160_out    = a11_wr[137];                 
			assign x1161_out    = a11_wr[1161];                
			assign x1162_out    = a11_wr[649];                 
			assign x1163_out    = a11_wr[1673];                
			assign x1164_out    = a11_wr[393];                 
			assign x1165_out    = a11_wr[1417];                
			assign x1166_out    = a11_wr[905];                 
			assign x1167_out    = a11_wr[1929];                
			assign x1168_out    = a11_wr[73];                  
			assign x1169_out    = a11_wr[1097];                
			assign x1170_out    = a11_wr[585];                 
			assign x1171_out    = a11_wr[1609];                
			assign x1172_out    = a11_wr[329];                 
			assign x1173_out    = a11_wr[1353];                
			assign x1174_out    = a11_wr[841];                 
			assign x1175_out    = a11_wr[1865];                
			assign x1176_out    = a11_wr[201];                 
			assign x1177_out    = a11_wr[1225];                
			assign x1178_out    = a11_wr[713];                 
			assign x1179_out    = a11_wr[1737];                
			assign x1180_out    = a11_wr[457];                 
			assign x1181_out    = a11_wr[1481];                
			assign x1182_out    = a11_wr[969];                 
			assign x1183_out    = a11_wr[1993];                
			assign x1184_out    = a11_wr[41];                  
			assign x1185_out    = a11_wr[1065];                
			assign x1186_out    = a11_wr[553];                 
			assign x1187_out    = a11_wr[1577];                
			assign x1188_out    = a11_wr[297];                 
			assign x1189_out    = a11_wr[1321];                
			assign x1190_out    = a11_wr[809];                 
			assign x1191_out    = a11_wr[1833];                
			assign x1192_out    = a11_wr[169];                 
			assign x1193_out    = a11_wr[1193];                
			assign x1194_out    = a11_wr[681];                 
			assign x1195_out    = a11_wr[1705];                
			assign x1196_out    = a11_wr[425];                 
			assign x1197_out    = a11_wr[1449];                
			assign x1198_out    = a11_wr[937];                 
			assign x1199_out    = a11_wr[1961];                
			assign x1200_out    = a11_wr[105];                 
			assign x1201_out    = a11_wr[1129];                
			assign x1202_out    = a11_wr[617];                 
			assign x1203_out    = a11_wr[1641];                
			assign x1204_out    = a11_wr[361];                 
			assign x1205_out    = a11_wr[1385];                
			assign x1206_out    = a11_wr[873];                 
			assign x1207_out    = a11_wr[1897];                
			assign x1208_out    = a11_wr[233];                 
			assign x1209_out    = a11_wr[1257];                
			assign x1210_out    = a11_wr[745];                 
			assign x1211_out    = a11_wr[1769];                
			assign x1212_out    = a11_wr[489];                 
			assign x1213_out    = a11_wr[1513];                
			assign x1214_out    = a11_wr[1001];                
			assign x1215_out    = a11_wr[2025];                
			assign x1216_out    = a11_wr[25];                  
			assign x1217_out    = a11_wr[1049];                
			assign x1218_out    = a11_wr[537];                 
			assign x1219_out    = a11_wr[1561];                
			assign x1220_out    = a11_wr[281];                 
			assign x1221_out    = a11_wr[1305];                
			assign x1222_out    = a11_wr[793];                 
			assign x1223_out    = a11_wr[1817];                
			assign x1224_out    = a11_wr[153];                 
			assign x1225_out    = a11_wr[1177];                
			assign x1226_out    = a11_wr[665];                 
			assign x1227_out    = a11_wr[1689];                
			assign x1228_out    = a11_wr[409];                 
			assign x1229_out    = a11_wr[1433];                
			assign x1230_out    = a11_wr[921];                 
			assign x1231_out    = a11_wr[1945];                
			assign x1232_out    = a11_wr[89];                  
			assign x1233_out    = a11_wr[1113];                
			assign x1234_out    = a11_wr[601];                 
			assign x1235_out    = a11_wr[1625];                
			assign x1236_out    = a11_wr[345];                 
			assign x1237_out    = a11_wr[1369];                
			assign x1238_out    = a11_wr[857];                 
			assign x1239_out    = a11_wr[1881];                
			assign x1240_out    = a11_wr[217];                 
			assign x1241_out    = a11_wr[1241];                
			assign x1242_out    = a11_wr[729];                 
			assign x1243_out    = a11_wr[1753];                
			assign x1244_out    = a11_wr[473];                 
			assign x1245_out    = a11_wr[1497];                
			assign x1246_out    = a11_wr[985];                 
			assign x1247_out    = a11_wr[2009];                
			assign x1248_out    = a11_wr[57];                  
			assign x1249_out    = a11_wr[1081];                
			assign x1250_out    = a11_wr[569];                 
			assign x1251_out    = a11_wr[1593];                
			assign x1252_out    = a11_wr[313];                 
			assign x1253_out    = a11_wr[1337];                
			assign x1254_out    = a11_wr[825];                 
			assign x1255_out    = a11_wr[1849];                
			assign x1256_out    = a11_wr[185];                 
			assign x1257_out    = a11_wr[1209];                
			assign x1258_out    = a11_wr[697];                 
			assign x1259_out    = a11_wr[1721];                
			assign x1260_out    = a11_wr[441];                 
			assign x1261_out    = a11_wr[1465];                
			assign x1262_out    = a11_wr[953];                 
			assign x1263_out    = a11_wr[1977];                
			assign x1264_out    = a11_wr[121];                 
			assign x1265_out    = a11_wr[1145];                
			assign x1266_out    = a11_wr[633];                 
			assign x1267_out    = a11_wr[1657];                
			assign x1268_out    = a11_wr[377];                 
			assign x1269_out    = a11_wr[1401];                
			assign x1270_out    = a11_wr[889];                 
			assign x1271_out    = a11_wr[1913];                
			assign x1272_out    = a11_wr[249];                 
			assign x1273_out    = a11_wr[1273];                
			assign x1274_out    = a11_wr[761];                 
			assign x1275_out    = a11_wr[1785];                
			assign x1276_out    = a11_wr[505];                 
			assign x1277_out    = a11_wr[1529];                
			assign x1278_out    = a11_wr[1017];                
			assign x1279_out    = a11_wr[2041];                
			assign x1280_out    = a11_wr[5];                   
			assign x1281_out    = a11_wr[1029];                
			assign x1282_out    = a11_wr[517];                 
			assign x1283_out    = a11_wr[1541];                
			assign x1284_out    = a11_wr[261];                 
			assign x1285_out    = a11_wr[1285];                
			assign x1286_out    = a11_wr[773];                 
			assign x1287_out    = a11_wr[1797];                
			assign x1288_out    = a11_wr[133];                 
			assign x1289_out    = a11_wr[1157];                
			assign x1290_out    = a11_wr[645];                 
			assign x1291_out    = a11_wr[1669];                
			assign x1292_out    = a11_wr[389];                 
			assign x1293_out    = a11_wr[1413];                
			assign x1294_out    = a11_wr[901];                 
			assign x1295_out    = a11_wr[1925];                
			assign x1296_out    = a11_wr[69];                  
			assign x1297_out    = a11_wr[1093];                
			assign x1298_out    = a11_wr[581];                 
			assign x1299_out    = a11_wr[1605];                
			assign x1300_out    = a11_wr[325];                 
			assign x1301_out    = a11_wr[1349];                
			assign x1302_out    = a11_wr[837];                 
			assign x1303_out    = a11_wr[1861];                
			assign x1304_out    = a11_wr[197];                 
			assign x1305_out    = a11_wr[1221];                
			assign x1306_out    = a11_wr[709];                 
			assign x1307_out    = a11_wr[1733];                
			assign x1308_out    = a11_wr[453];                 
			assign x1309_out    = a11_wr[1477];                
			assign x1310_out    = a11_wr[965];                 
			assign x1311_out    = a11_wr[1989];                
			assign x1312_out    = a11_wr[37];                  
			assign x1313_out    = a11_wr[1061];                
			assign x1314_out    = a11_wr[549];                 
			assign x1315_out    = a11_wr[1573];                
			assign x1316_out    = a11_wr[293];                 
			assign x1317_out    = a11_wr[1317];                
			assign x1318_out    = a11_wr[805];                 
			assign x1319_out    = a11_wr[1829];                
			assign x1320_out    = a11_wr[165];                 
			assign x1321_out    = a11_wr[1189];                
			assign x1322_out    = a11_wr[677];                 
			assign x1323_out    = a11_wr[1701];                
			assign x1324_out    = a11_wr[421];                 
			assign x1325_out    = a11_wr[1445];                
			assign x1326_out    = a11_wr[933];                 
			assign x1327_out    = a11_wr[1957];                
			assign x1328_out    = a11_wr[101];                 
			assign x1329_out    = a11_wr[1125];                
			assign x1330_out    = a11_wr[613];                 
			assign x1331_out    = a11_wr[1637];                
			assign x1332_out    = a11_wr[357];                 
			assign x1333_out    = a11_wr[1381];                
			assign x1334_out    = a11_wr[869];                 
			assign x1335_out    = a11_wr[1893];                
			assign x1336_out    = a11_wr[229];                 
			assign x1337_out    = a11_wr[1253];                
			assign x1338_out    = a11_wr[741];                 
			assign x1339_out    = a11_wr[1765];                
			assign x1340_out    = a11_wr[485];                 
			assign x1341_out    = a11_wr[1509];                
			assign x1342_out    = a11_wr[997];                 
			assign x1343_out    = a11_wr[2021];                
			assign x1344_out    = a11_wr[21];                  
			assign x1345_out    = a11_wr[1045];                
			assign x1346_out    = a11_wr[533];                 
			assign x1347_out    = a11_wr[1557];                
			assign x1348_out    = a11_wr[277];                 
			assign x1349_out    = a11_wr[1301];                
			assign x1350_out    = a11_wr[789];                 
			assign x1351_out    = a11_wr[1813];                
			assign x1352_out    = a11_wr[149];                 
			assign x1353_out    = a11_wr[1173];                
			assign x1354_out    = a11_wr[661];                 
			assign x1355_out    = a11_wr[1685];                
			assign x1356_out    = a11_wr[405];                 
			assign x1357_out    = a11_wr[1429];                
			assign x1358_out    = a11_wr[917];                 
			assign x1359_out    = a11_wr[1941];                
			assign x1360_out    = a11_wr[85];                  
			assign x1361_out    = a11_wr[1109];                
			assign x1362_out    = a11_wr[597];                 
			assign x1363_out    = a11_wr[1621];                
			assign x1364_out    = a11_wr[341];                 
			assign x1365_out    = a11_wr[1365];                
			assign x1366_out    = a11_wr[853];                 
			assign x1367_out    = a11_wr[1877];                
			assign x1368_out    = a11_wr[213];                 
			assign x1369_out    = a11_wr[1237];                
			assign x1370_out    = a11_wr[725];                 
			assign x1371_out    = a11_wr[1749];                
			assign x1372_out    = a11_wr[469];                 
			assign x1373_out    = a11_wr[1493];                
			assign x1374_out    = a11_wr[981];                 
			assign x1375_out    = a11_wr[2005];                
			assign x1376_out    = a11_wr[53];                  
			assign x1377_out    = a11_wr[1077];                
			assign x1378_out    = a11_wr[565];                 
			assign x1379_out    = a11_wr[1589];                
			assign x1380_out    = a11_wr[309];                 
			assign x1381_out    = a11_wr[1333];                
			assign x1382_out    = a11_wr[821];                 
			assign x1383_out    = a11_wr[1845];                
			assign x1384_out    = a11_wr[181];                 
			assign x1385_out    = a11_wr[1205];                
			assign x1386_out    = a11_wr[693];                 
			assign x1387_out    = a11_wr[1717];                
			assign x1388_out    = a11_wr[437];                 
			assign x1389_out    = a11_wr[1461];                
			assign x1390_out    = a11_wr[949];                 
			assign x1391_out    = a11_wr[1973];                
			assign x1392_out    = a11_wr[117];                 
			assign x1393_out    = a11_wr[1141];                
			assign x1394_out    = a11_wr[629];                 
			assign x1395_out    = a11_wr[1653];                
			assign x1396_out    = a11_wr[373];                 
			assign x1397_out    = a11_wr[1397];                
			assign x1398_out    = a11_wr[885];                 
			assign x1399_out    = a11_wr[1909];                
			assign x1400_out    = a11_wr[245];                 
			assign x1401_out    = a11_wr[1269];                
			assign x1402_out    = a11_wr[757];                 
			assign x1403_out    = a11_wr[1781];                
			assign x1404_out    = a11_wr[501];                 
			assign x1405_out    = a11_wr[1525];                
			assign x1406_out    = a11_wr[1013];                
			assign x1407_out    = a11_wr[2037];                
			assign x1408_out    = a11_wr[13];                  
			assign x1409_out    = a11_wr[1037];                
			assign x1410_out    = a11_wr[525];                 
			assign x1411_out    = a11_wr[1549];                
			assign x1412_out    = a11_wr[269];                 
			assign x1413_out    = a11_wr[1293];                
			assign x1414_out    = a11_wr[781];                 
			assign x1415_out    = a11_wr[1805];                
			assign x1416_out    = a11_wr[141];                 
			assign x1417_out    = a11_wr[1165];                
			assign x1418_out    = a11_wr[653];                 
			assign x1419_out    = a11_wr[1677];                
			assign x1420_out    = a11_wr[397];                 
			assign x1421_out    = a11_wr[1421];                
			assign x1422_out    = a11_wr[909];                 
			assign x1423_out    = a11_wr[1933];                
			assign x1424_out    = a11_wr[77];                  
			assign x1425_out    = a11_wr[1101];                
			assign x1426_out    = a11_wr[589];                 
			assign x1427_out    = a11_wr[1613];                
			assign x1428_out    = a11_wr[333];                 
			assign x1429_out    = a11_wr[1357];                
			assign x1430_out    = a11_wr[845];                 
			assign x1431_out    = a11_wr[1869];                
			assign x1432_out    = a11_wr[205];                 
			assign x1433_out    = a11_wr[1229];                
			assign x1434_out    = a11_wr[717];                 
			assign x1435_out    = a11_wr[1741];                
			assign x1436_out    = a11_wr[461];                 
			assign x1437_out    = a11_wr[1485];                
			assign x1438_out    = a11_wr[973];                 
			assign x1439_out    = a11_wr[1997];                
			assign x1440_out    = a11_wr[45];                  
			assign x1441_out    = a11_wr[1069];                
			assign x1442_out    = a11_wr[557];                 
			assign x1443_out    = a11_wr[1581];                
			assign x1444_out    = a11_wr[301];                 
			assign x1445_out    = a11_wr[1325];                
			assign x1446_out    = a11_wr[813];                 
			assign x1447_out    = a11_wr[1837];                
			assign x1448_out    = a11_wr[173];                 
			assign x1449_out    = a11_wr[1197];                
			assign x1450_out    = a11_wr[685];                 
			assign x1451_out    = a11_wr[1709];                
			assign x1452_out    = a11_wr[429];                 
			assign x1453_out    = a11_wr[1453];                
			assign x1454_out    = a11_wr[941];                 
			assign x1455_out    = a11_wr[1965];                
			assign x1456_out    = a11_wr[109];                 
			assign x1457_out    = a11_wr[1133];                
			assign x1458_out    = a11_wr[621];                 
			assign x1459_out    = a11_wr[1645];                
			assign x1460_out    = a11_wr[365];                 
			assign x1461_out    = a11_wr[1389];                
			assign x1462_out    = a11_wr[877];                 
			assign x1463_out    = a11_wr[1901];                
			assign x1464_out    = a11_wr[237];                 
			assign x1465_out    = a11_wr[1261];                
			assign x1466_out    = a11_wr[749];                 
			assign x1467_out    = a11_wr[1773];                
			assign x1468_out    = a11_wr[493];                 
			assign x1469_out    = a11_wr[1517];                
			assign x1470_out    = a11_wr[1005];                
			assign x1471_out    = a11_wr[2029];                
			assign x1472_out    = a11_wr[29];                  
			assign x1473_out    = a11_wr[1053];                
			assign x1474_out    = a11_wr[541];                 
			assign x1475_out    = a11_wr[1565];                
			assign x1476_out    = a11_wr[285];                 
			assign x1477_out    = a11_wr[1309];                
			assign x1478_out    = a11_wr[797];                 
			assign x1479_out    = a11_wr[1821];                
			assign x1480_out    = a11_wr[157];                 
			assign x1481_out    = a11_wr[1181];                
			assign x1482_out    = a11_wr[669];                 
			assign x1483_out    = a11_wr[1693];                
			assign x1484_out    = a11_wr[413];                 
			assign x1485_out    = a11_wr[1437];                
			assign x1486_out    = a11_wr[925];                 
			assign x1487_out    = a11_wr[1949];                
			assign x1488_out    = a11_wr[93];                  
			assign x1489_out    = a11_wr[1117];                
			assign x1490_out    = a11_wr[605];                 
			assign x1491_out    = a11_wr[1629];                
			assign x1492_out    = a11_wr[349];                 
			assign x1493_out    = a11_wr[1373];                
			assign x1494_out    = a11_wr[861];                 
			assign x1495_out    = a11_wr[1885];                
			assign x1496_out    = a11_wr[221];                 
			assign x1497_out    = a11_wr[1245];                
			assign x1498_out    = a11_wr[733];                 
			assign x1499_out    = a11_wr[1757];                
			assign x1500_out    = a11_wr[477];                 
			assign x1501_out    = a11_wr[1501];                
			assign x1502_out    = a11_wr[989];                 
			assign x1503_out    = a11_wr[2013];                
			assign x1504_out    = a11_wr[61];                  
			assign x1505_out    = a11_wr[1085];                
			assign x1506_out    = a11_wr[573];                 
			assign x1507_out    = a11_wr[1597];                
			assign x1508_out    = a11_wr[317];                 
			assign x1509_out    = a11_wr[1341];                
			assign x1510_out    = a11_wr[829];                 
			assign x1511_out    = a11_wr[1853];                
			assign x1512_out    = a11_wr[189];                 
			assign x1513_out    = a11_wr[1213];                
			assign x1514_out    = a11_wr[701];                 
			assign x1515_out    = a11_wr[1725];                
			assign x1516_out    = a11_wr[445];                 
			assign x1517_out    = a11_wr[1469];                
			assign x1518_out    = a11_wr[957];                 
			assign x1519_out    = a11_wr[1981];                
			assign x1520_out    = a11_wr[125];                 
			assign x1521_out    = a11_wr[1149];                
			assign x1522_out    = a11_wr[637];                 
			assign x1523_out    = a11_wr[1661];                
			assign x1524_out    = a11_wr[381];                 
			assign x1525_out    = a11_wr[1405];                
			assign x1526_out    = a11_wr[893];                 
			assign x1527_out    = a11_wr[1917];                
			assign x1528_out    = a11_wr[253];                 
			assign x1529_out    = a11_wr[1277];                
			assign x1530_out    = a11_wr[765];                 
			assign x1531_out    = a11_wr[1789];                
			assign x1532_out    = a11_wr[509];                 
			assign x1533_out    = a11_wr[1533];                
			assign x1534_out    = a11_wr[1021];                
			assign x1535_out    = a11_wr[2045];                
			assign x1536_out    = a11_wr[3];                   
			assign x1537_out    = a11_wr[1027];                
			assign x1538_out    = a11_wr[515];                 
			assign x1539_out    = a11_wr[1539];                
			assign x1540_out    = a11_wr[259];                 
			assign x1541_out    = a11_wr[1283];                
			assign x1542_out    = a11_wr[771];                 
			assign x1543_out    = a11_wr[1795];                
			assign x1544_out    = a11_wr[131];                 
			assign x1545_out    = a11_wr[1155];                
			assign x1546_out    = a11_wr[643];                 
			assign x1547_out    = a11_wr[1667];                
			assign x1548_out    = a11_wr[387];                 
			assign x1549_out    = a11_wr[1411];                
			assign x1550_out    = a11_wr[899];                 
			assign x1551_out    = a11_wr[1923];                
			assign x1552_out    = a11_wr[67];                  
			assign x1553_out    = a11_wr[1091];                
			assign x1554_out    = a11_wr[579];                 
			assign x1555_out    = a11_wr[1603];                
			assign x1556_out    = a11_wr[323];                 
			assign x1557_out    = a11_wr[1347];                
			assign x1558_out    = a11_wr[835];                 
			assign x1559_out    = a11_wr[1859];                
			assign x1560_out    = a11_wr[195];                 
			assign x1561_out    = a11_wr[1219];                
			assign x1562_out    = a11_wr[707];                 
			assign x1563_out    = a11_wr[1731];                
			assign x1564_out    = a11_wr[451];                 
			assign x1565_out    = a11_wr[1475];                
			assign x1566_out    = a11_wr[963];                 
			assign x1567_out    = a11_wr[1987];                
			assign x1568_out    = a11_wr[35];                  
			assign x1569_out    = a11_wr[1059];                
			assign x1570_out    = a11_wr[547];                 
			assign x1571_out    = a11_wr[1571];                
			assign x1572_out    = a11_wr[291];                 
			assign x1573_out    = a11_wr[1315];                
			assign x1574_out    = a11_wr[803];                 
			assign x1575_out    = a11_wr[1827];                
			assign x1576_out    = a11_wr[163];                 
			assign x1577_out    = a11_wr[1187];                
			assign x1578_out    = a11_wr[675];                 
			assign x1579_out    = a11_wr[1699];                
			assign x1580_out    = a11_wr[419];                 
			assign x1581_out    = a11_wr[1443];                
			assign x1582_out    = a11_wr[931];                 
			assign x1583_out    = a11_wr[1955];                
			assign x1584_out    = a11_wr[99];                  
			assign x1585_out    = a11_wr[1123];                
			assign x1586_out    = a11_wr[611];                 
			assign x1587_out    = a11_wr[1635];                
			assign x1588_out    = a11_wr[355];                 
			assign x1589_out    = a11_wr[1379];                
			assign x1590_out    = a11_wr[867];                 
			assign x1591_out    = a11_wr[1891];                
			assign x1592_out    = a11_wr[227];                 
			assign x1593_out    = a11_wr[1251];                
			assign x1594_out    = a11_wr[739];                 
			assign x1595_out    = a11_wr[1763];                
			assign x1596_out    = a11_wr[483];                 
			assign x1597_out    = a11_wr[1507];                
			assign x1598_out    = a11_wr[995];                 
			assign x1599_out    = a11_wr[2019];                
			assign x1600_out    = a11_wr[19];                  
			assign x1601_out    = a11_wr[1043];                
			assign x1602_out    = a11_wr[531];                 
			assign x1603_out    = a11_wr[1555];                
			assign x1604_out    = a11_wr[275];                 
			assign x1605_out    = a11_wr[1299];                
			assign x1606_out    = a11_wr[787];                 
			assign x1607_out    = a11_wr[1811];                
			assign x1608_out    = a11_wr[147];                 
			assign x1609_out    = a11_wr[1171];                
			assign x1610_out    = a11_wr[659];                 
			assign x1611_out    = a11_wr[1683];                
			assign x1612_out    = a11_wr[403];                 
			assign x1613_out    = a11_wr[1427];                
			assign x1614_out    = a11_wr[915];                 
			assign x1615_out    = a11_wr[1939];                
			assign x1616_out    = a11_wr[83];                  
			assign x1617_out    = a11_wr[1107];                
			assign x1618_out    = a11_wr[595];                 
			assign x1619_out    = a11_wr[1619];                
			assign x1620_out    = a11_wr[339];                 
			assign x1621_out    = a11_wr[1363];                
			assign x1622_out    = a11_wr[851];                 
			assign x1623_out    = a11_wr[1875];                
			assign x1624_out    = a11_wr[211];                 
			assign x1625_out    = a11_wr[1235];                
			assign x1626_out    = a11_wr[723];                 
			assign x1627_out    = a11_wr[1747];                
			assign x1628_out    = a11_wr[467];                 
			assign x1629_out    = a11_wr[1491];                
			assign x1630_out    = a11_wr[979];                 
			assign x1631_out    = a11_wr[2003];                
			assign x1632_out    = a11_wr[51];                  
			assign x1633_out    = a11_wr[1075];                
			assign x1634_out    = a11_wr[563];                 
			assign x1635_out    = a11_wr[1587];                
			assign x1636_out    = a11_wr[307];                 
			assign x1637_out    = a11_wr[1331];                
			assign x1638_out    = a11_wr[819];                 
			assign x1639_out    = a11_wr[1843];                
			assign x1640_out    = a11_wr[179];                 
			assign x1641_out    = a11_wr[1203];                
			assign x1642_out    = a11_wr[691];                 
			assign x1643_out    = a11_wr[1715];                
			assign x1644_out    = a11_wr[435];                 
			assign x1645_out    = a11_wr[1459];                
			assign x1646_out    = a11_wr[947];                 
			assign x1647_out    = a11_wr[1971];                
			assign x1648_out    = a11_wr[115];                 
			assign x1649_out    = a11_wr[1139];                
			assign x1650_out    = a11_wr[627];                 
			assign x1651_out    = a11_wr[1651];                
			assign x1652_out    = a11_wr[371];                 
			assign x1653_out    = a11_wr[1395];                
			assign x1654_out    = a11_wr[883];                 
			assign x1655_out    = a11_wr[1907];                
			assign x1656_out    = a11_wr[243];                 
			assign x1657_out    = a11_wr[1267];                
			assign x1658_out    = a11_wr[755];                 
			assign x1659_out    = a11_wr[1779];                
			assign x1660_out    = a11_wr[499];                 
			assign x1661_out    = a11_wr[1523];                
			assign x1662_out    = a11_wr[1011];                
			assign x1663_out    = a11_wr[2035];                
			assign x1664_out    = a11_wr[11];                  
			assign x1665_out    = a11_wr[1035];                
			assign x1666_out    = a11_wr[523];                 
			assign x1667_out    = a11_wr[1547];                
			assign x1668_out    = a11_wr[267];                 
			assign x1669_out    = a11_wr[1291];                
			assign x1670_out    = a11_wr[779];                 
			assign x1671_out    = a11_wr[1803];                
			assign x1672_out    = a11_wr[139];                 
			assign x1673_out    = a11_wr[1163];                
			assign x1674_out    = a11_wr[651];                 
			assign x1675_out    = a11_wr[1675];                
			assign x1676_out    = a11_wr[395];                 
			assign x1677_out    = a11_wr[1419];                
			assign x1678_out    = a11_wr[907];                 
			assign x1679_out    = a11_wr[1931];                
			assign x1680_out    = a11_wr[75];                  
			assign x1681_out    = a11_wr[1099];                
			assign x1682_out    = a11_wr[587];                 
			assign x1683_out    = a11_wr[1611];                
			assign x1684_out    = a11_wr[331];                 
			assign x1685_out    = a11_wr[1355];                
			assign x1686_out    = a11_wr[843];                 
			assign x1687_out    = a11_wr[1867];                
			assign x1688_out    = a11_wr[203];                 
			assign x1689_out    = a11_wr[1227];                
			assign x1690_out    = a11_wr[715];                 
			assign x1691_out    = a11_wr[1739];                
			assign x1692_out    = a11_wr[459];                 
			assign x1693_out    = a11_wr[1483];                
			assign x1694_out    = a11_wr[971];                 
			assign x1695_out    = a11_wr[1995];                
			assign x1696_out    = a11_wr[43];                  
			assign x1697_out    = a11_wr[1067];                
			assign x1698_out    = a11_wr[555];                 
			assign x1699_out    = a11_wr[1579];                
			assign x1700_out    = a11_wr[299];                 
			assign x1701_out    = a11_wr[1323];                
			assign x1702_out    = a11_wr[811];                 
			assign x1703_out    = a11_wr[1835];                
			assign x1704_out    = a11_wr[171];                 
			assign x1705_out    = a11_wr[1195];                
			assign x1706_out    = a11_wr[683];                 
			assign x1707_out    = a11_wr[1707];                
			assign x1708_out    = a11_wr[427];                 
			assign x1709_out    = a11_wr[1451];                
			assign x1710_out    = a11_wr[939];                 
			assign x1711_out    = a11_wr[1963];                
			assign x1712_out    = a11_wr[107];                 
			assign x1713_out    = a11_wr[1131];                
			assign x1714_out    = a11_wr[619];                 
			assign x1715_out    = a11_wr[1643];                
			assign x1716_out    = a11_wr[363];                 
			assign x1717_out    = a11_wr[1387];                
			assign x1718_out    = a11_wr[875];                 
			assign x1719_out    = a11_wr[1899];                
			assign x1720_out    = a11_wr[235];                 
			assign x1721_out    = a11_wr[1259];                
			assign x1722_out    = a11_wr[747];                 
			assign x1723_out    = a11_wr[1771];                
			assign x1724_out    = a11_wr[491];                 
			assign x1725_out    = a11_wr[1515];                
			assign x1726_out    = a11_wr[1003];                
			assign x1727_out    = a11_wr[2027];                
			assign x1728_out    = a11_wr[27];                  
			assign x1729_out    = a11_wr[1051];                
			assign x1730_out    = a11_wr[539];                 
			assign x1731_out    = a11_wr[1563];                
			assign x1732_out    = a11_wr[283];                 
			assign x1733_out    = a11_wr[1307];                
			assign x1734_out    = a11_wr[795];                 
			assign x1735_out    = a11_wr[1819];                
			assign x1736_out    = a11_wr[155];                 
			assign x1737_out    = a11_wr[1179];                
			assign x1738_out    = a11_wr[667];                 
			assign x1739_out    = a11_wr[1691];                
			assign x1740_out    = a11_wr[411];                 
			assign x1741_out    = a11_wr[1435];                
			assign x1742_out    = a11_wr[923];                 
			assign x1743_out    = a11_wr[1947];                
			assign x1744_out    = a11_wr[91];                  
			assign x1745_out    = a11_wr[1115];                
			assign x1746_out    = a11_wr[603];                 
			assign x1747_out    = a11_wr[1627];                
			assign x1748_out    = a11_wr[347];                 
			assign x1749_out    = a11_wr[1371];                
			assign x1750_out    = a11_wr[859];                 
			assign x1751_out    = a11_wr[1883];                
			assign x1752_out    = a11_wr[219];                 
			assign x1753_out    = a11_wr[1243];                
			assign x1754_out    = a11_wr[731];                 
			assign x1755_out    = a11_wr[1755];                
			assign x1756_out    = a11_wr[475];                 
			assign x1757_out    = a11_wr[1499];                
			assign x1758_out    = a11_wr[987];                 
			assign x1759_out    = a11_wr[2011];                
			assign x1760_out    = a11_wr[59];                  
			assign x1761_out    = a11_wr[1083];                
			assign x1762_out    = a11_wr[571];                 
			assign x1763_out    = a11_wr[1595];                
			assign x1764_out    = a11_wr[315];                 
			assign x1765_out    = a11_wr[1339];                
			assign x1766_out    = a11_wr[827];                 
			assign x1767_out    = a11_wr[1851];                
			assign x1768_out    = a11_wr[187];                 
			assign x1769_out    = a11_wr[1211];                
			assign x1770_out    = a11_wr[699];                 
			assign x1771_out    = a11_wr[1723];                
			assign x1772_out    = a11_wr[443];                 
			assign x1773_out    = a11_wr[1467];                
			assign x1774_out    = a11_wr[955];                 
			assign x1775_out    = a11_wr[1979];                
			assign x1776_out    = a11_wr[123];                 
			assign x1777_out    = a11_wr[1147];                
			assign x1778_out    = a11_wr[635];                 
			assign x1779_out    = a11_wr[1659];                
			assign x1780_out    = a11_wr[379];                 
			assign x1781_out    = a11_wr[1403];                
			assign x1782_out    = a11_wr[891];                 
			assign x1783_out    = a11_wr[1915];                
			assign x1784_out    = a11_wr[251];                 
			assign x1785_out    = a11_wr[1275];                
			assign x1786_out    = a11_wr[763];                 
			assign x1787_out    = a11_wr[1787];                
			assign x1788_out    = a11_wr[507];                 
			assign x1789_out    = a11_wr[1531];                
			assign x1790_out    = a11_wr[1019];                
			assign x1791_out    = a11_wr[2043];                
			assign x1792_out    = a11_wr[7];                   
			assign x1793_out    = a11_wr[1031];                
			assign x1794_out    = a11_wr[519];                 
			assign x1795_out    = a11_wr[1543];                
			assign x1796_out    = a11_wr[263];                 
			assign x1797_out    = a11_wr[1287];                
			assign x1798_out    = a11_wr[775];                 
			assign x1799_out    = a11_wr[1799];                
			assign x1800_out    = a11_wr[135];                 
			assign x1801_out    = a11_wr[1159];                
			assign x1802_out    = a11_wr[647];                 
			assign x1803_out    = a11_wr[1671];                
			assign x1804_out    = a11_wr[391];                 
			assign x1805_out    = a11_wr[1415];                
			assign x1806_out    = a11_wr[903];                 
			assign x1807_out    = a11_wr[1927];                
			assign x1808_out    = a11_wr[71];                  
			assign x1809_out    = a11_wr[1095];                
			assign x1810_out    = a11_wr[583];                 
			assign x1811_out    = a11_wr[1607];                
			assign x1812_out    = a11_wr[327];                 
			assign x1813_out    = a11_wr[1351];                
			assign x1814_out    = a11_wr[839];                 
			assign x1815_out    = a11_wr[1863];                
			assign x1816_out    = a11_wr[199];                 
			assign x1817_out    = a11_wr[1223];                
			assign x1818_out    = a11_wr[711];                 
			assign x1819_out    = a11_wr[1735];                
			assign x1820_out    = a11_wr[455];                 
			assign x1821_out    = a11_wr[1479];                
			assign x1822_out    = a11_wr[967];                 
			assign x1823_out    = a11_wr[1991];                
			assign x1824_out    = a11_wr[39];                  
			assign x1825_out    = a11_wr[1063];                
			assign x1826_out    = a11_wr[551];                 
			assign x1827_out    = a11_wr[1575];                
			assign x1828_out    = a11_wr[295];                 
			assign x1829_out    = a11_wr[1319];                
			assign x1830_out    = a11_wr[807];                 
			assign x1831_out    = a11_wr[1831];                
			assign x1832_out    = a11_wr[167];                 
			assign x1833_out    = a11_wr[1191];                
			assign x1834_out    = a11_wr[679];                 
			assign x1835_out    = a11_wr[1703];                
			assign x1836_out    = a11_wr[423];                 
			assign x1837_out    = a11_wr[1447];                
			assign x1838_out    = a11_wr[935];                 
			assign x1839_out    = a11_wr[1959];                
			assign x1840_out    = a11_wr[103];                 
			assign x1841_out    = a11_wr[1127];                
			assign x1842_out    = a11_wr[615];                 
			assign x1843_out    = a11_wr[1639];                
			assign x1844_out    = a11_wr[359];                 
			assign x1845_out    = a11_wr[1383];                
			assign x1846_out    = a11_wr[871];                 
			assign x1847_out    = a11_wr[1895];                
			assign x1848_out    = a11_wr[231];                 
			assign x1849_out    = a11_wr[1255];                
			assign x1850_out    = a11_wr[743];                 
			assign x1851_out    = a11_wr[1767];                
			assign x1852_out    = a11_wr[487];                 
			assign x1853_out    = a11_wr[1511];                
			assign x1854_out    = a11_wr[999];                 
			assign x1855_out    = a11_wr[2023];                
			assign x1856_out    = a11_wr[23];                  
			assign x1857_out    = a11_wr[1047];                
			assign x1858_out    = a11_wr[535];                 
			assign x1859_out    = a11_wr[1559];                
			assign x1860_out    = a11_wr[279];                 
			assign x1861_out    = a11_wr[1303];                
			assign x1862_out    = a11_wr[791];                 
			assign x1863_out    = a11_wr[1815];                
			assign x1864_out    = a11_wr[151];                 
			assign x1865_out    = a11_wr[1175];                
			assign x1866_out    = a11_wr[663];                 
			assign x1867_out    = a11_wr[1687];                
			assign x1868_out    = a11_wr[407];                 
			assign x1869_out    = a11_wr[1431];                
			assign x1870_out    = a11_wr[919];                 
			assign x1871_out    = a11_wr[1943];                
			assign x1872_out    = a11_wr[87];                  
			assign x1873_out    = a11_wr[1111];                
			assign x1874_out    = a11_wr[599];                 
			assign x1875_out    = a11_wr[1623];                
			assign x1876_out    = a11_wr[343];                 
			assign x1877_out    = a11_wr[1367];                
			assign x1878_out    = a11_wr[855];                 
			assign x1879_out    = a11_wr[1879];                
			assign x1880_out    = a11_wr[215];                 
			assign x1881_out    = a11_wr[1239];                
			assign x1882_out    = a11_wr[727];                 
			assign x1883_out    = a11_wr[1751];                
			assign x1884_out    = a11_wr[471];                 
			assign x1885_out    = a11_wr[1495];                
			assign x1886_out    = a11_wr[983];                 
			assign x1887_out    = a11_wr[2007];                
			assign x1888_out    = a11_wr[55];                  
			assign x1889_out    = a11_wr[1079];                
			assign x1890_out    = a11_wr[567];                 
			assign x1891_out    = a11_wr[1591];                
			assign x1892_out    = a11_wr[311];                 
			assign x1893_out    = a11_wr[1335];                
			assign x1894_out    = a11_wr[823];                 
			assign x1895_out    = a11_wr[1847];                
			assign x1896_out    = a11_wr[183];                 
			assign x1897_out    = a11_wr[1207];                
			assign x1898_out    = a11_wr[695];                 
			assign x1899_out    = a11_wr[1719];                
			assign x1900_out    = a11_wr[439];                 
			assign x1901_out    = a11_wr[1463];                
			assign x1902_out    = a11_wr[951];                 
			assign x1903_out    = a11_wr[1975];                
			assign x1904_out    = a11_wr[119];                 
			assign x1905_out    = a11_wr[1143];                
			assign x1906_out    = a11_wr[631];                 
			assign x1907_out    = a11_wr[1655];                
			assign x1908_out    = a11_wr[375];                 
			assign x1909_out    = a11_wr[1399];                
			assign x1910_out    = a11_wr[887];                 
			assign x1911_out    = a11_wr[1911];                
			assign x1912_out    = a11_wr[247];                 
			assign x1913_out    = a11_wr[1271];                
			assign x1914_out    = a11_wr[759];                 
			assign x1915_out    = a11_wr[1783];                
			assign x1916_out    = a11_wr[503];                 
			assign x1917_out    = a11_wr[1527];                
			assign x1918_out    = a11_wr[1015];                
			assign x1919_out    = a11_wr[2039];                
			assign x1920_out    = a11_wr[15];                  
			assign x1921_out    = a11_wr[1039];                
			assign x1922_out    = a11_wr[527];                 
			assign x1923_out    = a11_wr[1551];                
			assign x1924_out    = a11_wr[271];                 
			assign x1925_out    = a11_wr[1295];                
			assign x1926_out    = a11_wr[783];                 
			assign x1927_out    = a11_wr[1807];                
			assign x1928_out    = a11_wr[143];                 
			assign x1929_out    = a11_wr[1167];                
			assign x1930_out    = a11_wr[655];                 
			assign x1931_out    = a11_wr[1679];                
			assign x1932_out    = a11_wr[399];                 
			assign x1933_out    = a11_wr[1423];                
			assign x1934_out    = a11_wr[911];                 
			assign x1935_out    = a11_wr[1935];                
			assign x1936_out    = a11_wr[79];                  
			assign x1937_out    = a11_wr[1103];                
			assign x1938_out    = a11_wr[591];                 
			assign x1939_out    = a11_wr[1615];                
			assign x1940_out    = a11_wr[335];                 
			assign x1941_out    = a11_wr[1359];                
			assign x1942_out    = a11_wr[847];                 
			assign x1943_out    = a11_wr[1871];                
			assign x1944_out    = a11_wr[207];                 
			assign x1945_out    = a11_wr[1231];                
			assign x1946_out    = a11_wr[719];                 
			assign x1947_out    = a11_wr[1743];                
			assign x1948_out    = a11_wr[463];                 
			assign x1949_out    = a11_wr[1487];                
			assign x1950_out    = a11_wr[975];                 
			assign x1951_out    = a11_wr[1999];                
			assign x1952_out    = a11_wr[47];                  
			assign x1953_out    = a11_wr[1071];                
			assign x1954_out    = a11_wr[559];                 
			assign x1955_out    = a11_wr[1583];                
			assign x1956_out    = a11_wr[303];                 
			assign x1957_out    = a11_wr[1327];                
			assign x1958_out    = a11_wr[815];                 
			assign x1959_out    = a11_wr[1839];                
			assign x1960_out    = a11_wr[175];                 
			assign x1961_out    = a11_wr[1199];                
			assign x1962_out    = a11_wr[687];                 
			assign x1963_out    = a11_wr[1711];                
			assign x1964_out    = a11_wr[431];                 
			assign x1965_out    = a11_wr[1455];                
			assign x1966_out    = a11_wr[943];                 
			assign x1967_out    = a11_wr[1967];                
			assign x1968_out    = a11_wr[111];                 
			assign x1969_out    = a11_wr[1135];                
			assign x1970_out    = a11_wr[623];                 
			assign x1971_out    = a11_wr[1647];                
			assign x1972_out    = a11_wr[367];                 
			assign x1973_out    = a11_wr[1391];                
			assign x1974_out    = a11_wr[879];                 
			assign x1975_out    = a11_wr[1903];                
			assign x1976_out    = a11_wr[239];                 
			assign x1977_out    = a11_wr[1263];                
			assign x1978_out    = a11_wr[751];                 
			assign x1979_out    = a11_wr[1775];                
			assign x1980_out    = a11_wr[495];                 
			assign x1981_out    = a11_wr[1519];                
			assign x1982_out    = a11_wr[1007];                
			assign x1983_out    = a11_wr[2031];                
			assign x1984_out    = a11_wr[31];                  
			assign x1985_out    = a11_wr[1055];                
			assign x1986_out    = a11_wr[543];                 
			assign x1987_out    = a11_wr[1567];                
			assign x1988_out    = a11_wr[287];                 
			assign x1989_out    = a11_wr[1311];                
			assign x1990_out    = a11_wr[799];                 
			assign x1991_out    = a11_wr[1823];                
			assign x1992_out    = a11_wr[159];                 
			assign x1993_out    = a11_wr[1183];                
			assign x1994_out    = a11_wr[671];                 
			assign x1995_out    = a11_wr[1695];                
			assign x1996_out    = a11_wr[415];                 
			assign x1997_out    = a11_wr[1439];                
			assign x1998_out    = a11_wr[927];                 
			assign x1999_out    = a11_wr[1951];                
			assign x2000_out    = a11_wr[95];                  
			assign x2001_out    = a11_wr[1119];                
			assign x2002_out    = a11_wr[607];                 
			assign x2003_out    = a11_wr[1631];                
			assign x2004_out    = a11_wr[351];                 
			assign x2005_out    = a11_wr[1375];                
			assign x2006_out    = a11_wr[863];                 
			assign x2007_out    = a11_wr[1887];                
			assign x2008_out    = a11_wr[223];                 
			assign x2009_out    = a11_wr[1247];                
			assign x2010_out    = a11_wr[735];                 
			assign x2011_out    = a11_wr[1759];                
			assign x2012_out    = a11_wr[479];                 
			assign x2013_out    = a11_wr[1503];                
			assign x2014_out    = a11_wr[991];                 
			assign x2015_out    = a11_wr[2015];                
			assign x2016_out    = a11_wr[63];                  
			assign x2017_out    = a11_wr[1087];                
			assign x2018_out    = a11_wr[575];                 
			assign x2019_out    = a11_wr[1599];                
			assign x2020_out    = a11_wr[319];                 
			assign x2021_out    = a11_wr[1343];                
			assign x2022_out    = a11_wr[831];                 
			assign x2023_out    = a11_wr[1855];                
			assign x2024_out    = a11_wr[191];                 
			assign x2025_out    = a11_wr[1215];                
			assign x2026_out    = a11_wr[703];                 
			assign x2027_out    = a11_wr[1727];                
			assign x2028_out    = a11_wr[447];                 
			assign x2029_out    = a11_wr[1471];                
			assign x2030_out    = a11_wr[959];                 
			assign x2031_out    = a11_wr[1983];                
			assign x2032_out    = a11_wr[127];                 
			assign x2033_out    = a11_wr[1151];                
			assign x2034_out    = a11_wr[639];                 
			assign x2035_out    = a11_wr[1663];                
			assign x2036_out    = a11_wr[383];                 
			assign x2037_out    = a11_wr[1407];                
			assign x2038_out    = a11_wr[895];                 
			assign x2039_out    = a11_wr[1919];                
			assign x2040_out    = a11_wr[255];                 
			assign x2041_out    = a11_wr[1279];                
			assign x2042_out    = a11_wr[767];                 
			assign x2043_out    = a11_wr[1791];                
			assign x2044_out    = a11_wr[511];                 
			assign x2045_out    = a11_wr[1535];                
			assign x2046_out    = a11_wr[1023];                
			assign x2047_out    = a11_wr[2047];                


endmodule
