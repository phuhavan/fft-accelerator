`include "localmem_defines.h"

//======================================================

module mul_tw
(
	input	[`DM_BANK_COLS-1:0] in0,
	input	[`DM_BANK_COLS-1:0] in1,
	output	[`DM_BANK_COLS-1:0] out0
);

endmodule